`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
KknvL6SYSb5dRFuWP4AJqBhO3b64YXO1jXJrKEg0Z3ikGAO3obMtU40YwJiJW7ipQ08/Y8WRYNWh
nV2LdqH0dA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QLUbVPatcj7IWeOM7GaVpOxxKXKrfEAPdOAPmfRnpcapAKHnvWUhcysRYZ/rY/73FKWInR8HJilV
JFgxROZVCNWQ1zJhGgmKt04WHahOu9miHsfm8H7yNJ6k3TsDqjbc8beG5UCVgF6x/gDB8LRb2Vlo
OYeUOl3UjHyll8Sbd9I=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4fDulW+j2qCXqz735RjXksliYlPtal97cQEPC5accAQtxDw7TbdSqrHOiG5KctOIuaRzvRMOO5x
8R7f4K2bkMvIUjiiFP5Xw/fjJySLFuOiZoiNxxNdz5n6QQgBWYDepruKbEU7yj9zlmf0zEFmWZo2
ShS1WpLwP3B9Mcm5hJ+0GZ0wSeVmrvJEKp8kqO3uW6EVpKbiSMmBugVkGUzz9ZrIbzEZlELi+wJ/
HVgQM4hNwGKaRhAKNMJGLkgs6Mi/pI+CqjdrjRYK0X20OxPYi7+y3i6gUy//rkWJVRVSqqxJt07h
XfBm/2egXCeHNQMVyg/cuW80bFPZUcKb/tb28A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eEHF/HRqboErONr15dWGPiKIhHmEp89NzpKM1HVNOPxPMAhm5Q7SHcs30Gyp606YzPvXAWOwIhp6
yShxWJQDMNzjx8XLNdk6Hk4q1OFOlxJvftzg6IwFePhX6CX5M/h6gWDjhSncOnYuNt1s46FrBJGA
DJZ7AbtD39aEQbpRrtRqPKdh74/RGoSXOsksuOHq//+3LZGY5WN1wdVNJTew5IKMLtb98TYlHOO4
w28CobD4NywkdWMYWBeN1weCfLySyzftQavfk/dRUoBAG4mBbSm67pDUnjTuzD/BMIiEezbjKgGt
v5JKng8K28aaFylCDbrjWbQ4f0E0MG89P9bqcQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LBodvKMdQLsL3NITg6iyfn6uEr0nsFsSECbcpJ0VM9GPtNyhu1PCIqop74QUK0jX7gNod2kXTA0j
UPAVU1VbFsW+W9odvoIvVhgiIvptX2ncKxVnQVrYamDTZTPdFxs85ZcmhfukKF1ctZJMx5QHtsT8
/fgDo9EnaiAwUK6EH1vPn8nlJtMakUlaKARMU1hnWHBUkjruM2J062f3fYCx1Fc0yI51VXZXtNw2
A35SpeR68WKPmXnaWtRfYcT55OhdStBuASxbBHMItu7IQi56vUWP8LJm5L8r7e0VPvAGmJGTHM8m
DRb2QSYwaQDB32Ac/WNT/HueDTeVlvRT+cXLnQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RTdH2QVRkLMNeDjWHM39MNQI9JpZeMEnnaFqgJIEgBuj3R1/oXRV+h+0yVRQ+SMug8jz9no0jCSS
W3wRM89ooYAXiOYt8RwiQibqZKat+R7T7m3thhmgMEI8uoi9fGuXrcwO/YAOvNwNOuRc5iytwydq
EbyW4aM2m+CrXKFlD7s=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hNd+z0nXH9GYvgjnhDJoJvhFhK8AT6oUoCmTuJoXrdeSPSICu0d2AmfE/9zKTVob1byyZNQ+dZJb
Ma+7SxXV1+3xFvececBxzrOjVMq4geH8T4yeo12KR/tsEogGtiBVtNuwOoiOTxmMqj4v1JDOa2o8
G9PU/lTBUSoEzibdcIpQyhvP7Mdz6AOWlVWthHuCNvffk52oBkFkYg/wxqRli9uZ+ljnrd6rXIeN
pcjEkI9ALbBEAZnGGMY3do4kdn+d4UrzbiC/0FwIrw+uZYeWK2+A1bCZ3JcBMczd2lYYJYQOACWj
1dr/Sij9Dnl2NTdY6Acp6dQAwn2oASr3Hs8Onw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2480)
`pragma protect data_block
F4D6nIAHG9w7CzDjTOGl433b/ii9ahOx8+IfkLmcfM8G6T7LM4/Frrx3cn9UsUko2x/qD8Q/qCyu
TrwRUdjKWMC4Fc5bAjjUZgbTWgyAHHAy2hpz4B4ocPTIwHvLZuJapDRkAxNr73Z3OCc++uPgjOBZ
3zuq0xrZCwMgFBuyBAqR/HUQYa1mO04ylZjdZ2SeeVKy6es8A/SeJzrlRq9JqfOHIIQCN+3g4Tav
U7uCMrg0Urbno/NQ2/vPldi+sbj2P+dqztE0RJ6Hd3opBpPfdafqoR6virfk3FL0K0pD7vFUUlDC
i9ukhwJaekkdaxmnVWXuPD6v5jVTYdnqPoiLuAv4KYVg61F45h6B3JPj/9ixgb3T313LGOueFfxg
LfmwHwnSqsczI9IoBQ45ZCaaY+U4Tb0jZHDjandZ6XzRYV9kIKIBj3RIzomdgv4PIA7bXvIAOdsH
V+xbeUDty/38RX4D7W/j65yxN9sK5KVA7yLrjuy60qeM68FcakKx6HTf2ztRpJB1ke72nXdvmhCh
ItrlyyHkFh8EcBE9r0/Zl0NATDNjFZ5V5k4A47kuNGUs5h8x8ENVHNyQGywLieEVu80Q/lbDMMAn
cYpK4b41a+H9rcFnCEEETzaH6k02qt4L9xtej5bbv7TZmkiBKsCB/cQ6RmVQOT4scIo9j3mD+41U
FgM/9l/XKo2vJD+W2uOTpXkdSYNak2zu5kSYfPvcB66speAoizwaah33sCPkz9XGgzsdI+wZYnux
saKJmJBdTXYhz0F2B1oC4eCg/zuc4kDXTCcipT42+ZJqXif4/1NSHaBorZBe0slMxY9s816/vtDJ
kbFb9ExYXaGJK2LQ5atYrFmFAFl+uHK61vaRoJoOwGXKd69PDkNxbbq6tqysW2XQBBzyHNTcQP66
m/CTxYH6BLZEFcsmSd+h/wCta7CuQaqOL+srwC+D5/pzHQCPtNrl7uUtU2ilsteycK/NZZa7f5N8
bmTcFTXt8IcVk1mWE5uMcwtCbVg14c+AInOhUPgpiu55ycLi2HWLvDuK5K/YQKyK7p06jtXm8nc1
B3ltgFe2FvWbxeFmMWwF/X+C2Ro5S/yEanaXRG/k0PPzKTBW6+tYy5qR6RSNBdp6JdAxB4Kcht7U
6pkjPOjdgfjJXRqGuUixkChL9g+2MQupYLH/lX33P8/IQM7AgiqQmJbhLxg6mLo3WCnt0f19gzW1
BtgiezRIS+tp6q6DCCVJrjQNJFgRIdpg0um0lhhRpyfoLBHsxUt4i5dqfpG4t/7nVZp25yHvGAz8
ImN5SIxD4hTf5hc/RjBzJs3ppytIHJ21q66sQqVoShEsmBbyjr72pIlmza3DzlAnne5yQ9H3NfDB
d6XkZ6tLUDa3cX7Ydrldeb3bNkxEr0kNOypGdTebb9a5si211GlztvgAQOhxm2fj4Swgjxd2F+tk
TuZNAVtX1tFaCtBYUICgpUyIUV2eXdrM0j4+OEGUQNzgKqS2wOBMAnOupUGQY91ocfZMvCIjplp9
LzHzsCwpWCYucEnWrHJk5eSUZ5Zop/9FIgjuIQ+VvDItYdsJPgvvwN7vYOfBfSjU3qgyWERbl1jb
eT7aAsni5a62PeBY7X9ZgNLvF+EaudNlj6DWKUi7mvoIIK+vrVpUBlw2UEL8XILqo/15Gf6EKMhO
+FU7zVxiw7vQc2GrLmIrnJ9w5x0CM/Awpt4M51+CDeUGN5WTW6CnNAMjBvGb9E3EfTDKeay5l5NP
jeBcpcVbDMnPxOZpm01x3FvW8Rk+NXPt8fvFrFKvFg8wC85lsyYirHKQPXItxKO9pIodsfv47uKY
LYKfye4Tb4bbukmGjPGx0VpLOU81Ms6X70LYFZk1Yh4a8UkATYiT2fIVDkwX8cUiK8ifZ/VRsBHi
VE7zBZhd5Kp49aogU2no5ISQKdd3yblHk6uriBgU3DxCPyl9RSYrOg56iQyXijPuS4M63lRiL4kd
pkCXjulr32X5WK11NSd3NNQkNuO1bWdAAwC0b4ZXmFYAE2BMuK/uDEvvJvupmruOZS8+T4SDewGB
ouhRIx4lQJ+3ozhlAxMWOnpgiaKI5JIu6ITSTfHPnchpR0QqClMZ7xlh8qWFTZsiUXHBV8iENPP0
AdcWALHFUX7cnd2cvvJd/1pjHl7ORyBgNoropb0U9N3La80U4PkNxYfkBDXwCvqj/aMMkT5DYfQx
zkSf6bMLEgMn8JJ832iqJUi6nRcJSFp8SKj3tNNRIkTx+G+H5UmYMuP37X0NggkXoj2lj51mbxyR
8VCoCt1F+Pu74/iXCXCvrHsj+omwMTVElebwmQsycYeovn/7fGJjKVpjcZuG91NjLhvOFlN2vosd
nhfq7unr3ttxu9b2M8abVHIVdajp5RWT4FGiEhhtS+dbwGUQs9tRFXl4QoJ3WqlJUqyb93TdHIQM
t2Qut+SNQglqly5Gh6iVEkcmVNpf8588juoEYGWCKQEXBppKgihtFWU0p7Fcw5opHFlv0dZVTFTu
fs037/Obt9uQ6XHjEHiSNRMdiKy1RaYPLPjP82y7wlKnOmIzpdSlHPVqvfSDSxclo5+JFfW07bMv
QheQ/+dDWy+Pkgi4HyhnMywzYUFa1YPe7KoosdcbVJl6AKLytYHEq8S701MP+dIUv4asnfZ1uZgY
mjsJYGGUqOmNb3kx0Qvlf0bGdfgTo7gLZBm3rvpxrEAtldBuZSHA6Qozsoq6NrOOKMBIbMECyhzo
sf/T3MRSVmWbiCMsnTklGMZV39e1O6mL2wvkv9Ek++O/Lp+tN5fjk29DAAdOxKACKlwFywEx89cE
XfEqScgQvCeMvixVMOItTVdHEVh4gFbb36xajc0GInVPzvcL4KsMrd6u94CgjMNWCclXexDfA8Bk
XPfV+z+dDW1CNOTe5IVQKTqMd3I+q3XQkwjegw53SQQQSZiOV2GnnTsht+GN4wEcSrR+MoAwdDG4
gzi2eJEy5T15uWggR0R2RmIncZeGB0HPRh9LfmDUwaPicIRX9TZOJXjVA7aRvrWvWhs+wIEhuruj
BvPk1nnG4iQZLKrkk2AA4r+Mxi5xp/vInnUAjDuHODQr0HB9+TOInOHkIM6vogd6xWc0iiUuTaUf
kjX2EmFSYCzfSVQ793zvfa1Zdm3GOKm3LS4PkTKjQPjCYqcWUOhJZc0SZ30DCjgdmppsJqV1CzSG
UGw5Jy2cyvQ/n1sculIDezD0srykh8lVvQIpWUVs93dwLUW1+uFll8YIk1q7tVoXBhmNuFzG8DQP
gVDnquP/uoN6pM7/GyrA6QbidwI2Wp2krKQiYbw=
`pragma protect end_protected
