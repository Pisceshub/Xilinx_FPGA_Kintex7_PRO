`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69264)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9JR+2FTwzOkJ1yLmnse46t3GbkqvKGdMPXCsVU97ufEdNV6W4u47IL58
Jnz8MyoPlqMjtlqhzRXXLit4FW7q1CEeRroKbHBJmfNijs1tjBaOT7URGEqz/N/ORUCJc7b6YDID
flYJi5KZgm+BbtWEB22qHAKg3jeiS3/tmCorTq1805PglLyk/xUU69tOBuB0vkPOt41Q6NgevKCm
Q8rcnqlfQ24FC+0kus0sHxmFPiVPkxd64IUpPdhMsAPzX21ILChmMZDqvWW5PtTqz7EJSX7cQCxI
/oO2hT9FNVIw3ilpb2ctfg9y5wYDfCm+8IwtY8REssF4bcjUbDBND3s1yg3PMmCVJ6+c83nR8zHd
zG3035fdmQ7u2GOZB2WDcOEFPC2mT/epggNvW8vI8m33oENF7Tz8ihEOLvbxpPkif5DaKWkQmyPU
4CV9cnHX7uwVXU0LUA01dotoM1fL9+gvyV0GRwAIDeRJn0EvvGixmMtlqIe1Wn8tOskKK6tPO758
zaLIsV1mEAZ0jnwsi0WMQo2bAKlJ+JDhURLsk1Oy6uJZ90bpSgFP6JSddk6gJRnaxfsU9a3X0rBp
pUx5szbACvpU5L4im5MaKipLwD2C+o8Slt7SWKiNaztZCVyLjgXAY9+jDaDkHdmsNfVqOHmyeAAI
fwjd1RmER3T6UGdv03yAJrh/w0UGjKWO3vi+ZSDu6GDldeDGf8DKDGRsSnAduHpY9vSawEThAbsa
EJ//RhIJZKi1/BOWX00uHqFmyAqDna5PwsacGX0z3CMFPIN7Mlk165plQvg4FvbNA9Vbi4wGRuTl
heeProYy9laMNRPLKYwp7tIprmSOJtrsch8xktcy6W558AKpP1Y2wJ3BgOqScZqiwFa1NS70M9Wl
tfo+GA3Ck6g5gopAFTa/g3q9WVHMPOvVWdvQByegfABs7AJPLIuAVFoDBIC66OdSX3KzRJyn0uaa
v0ecYgZ06DDCtnEfj0Ev19cuqdQ9kbzSxNPxmEsw2eC5hjYScsRAO+psBDsCSf+72yz5b2F9WYWy
WayY7Vq7d6gPm1MScSBfFDkGDMnOKNYWWyyMDPRwuYfNA9z4K+RzRThNTcABxFytHjlPrSsxhc1P
AcefD9T0xbJdGGaTEv0HPhwbLNTpqx0e9k+K/q2U77ldVPhOzrtAMSNwfh+ieWeZ8/Bri0Vf8iQ2
4RAR/Ilp0xVcLh9J7/V8t3MFoYNqbPOQAvYXeLSYxTb1HBKgxyT+EMUrSHeZOYX/Tq3iFVQdySQ+
TlHKgzjmNDoISe3ex80Q0J3FQrAMJ6QXmuQ+80SwJtW1mk5OJwUtalH9C+VudOYPC0gcY2y6bCWT
9ztt8sKYSc5ZK+vRiMu2/ib254KvyliVMr2LjpEfz/L1oarH2+vWzyx90CZ2zonuOT0nSuqBb9D6
tFW4ArD6JcjI10h4WSiu4Ulb9v/UAaQv6uTNQCLGMj6d9/3piaht0JclC/sYZToy7WmvOTM9KIKK
KO1JMoIsUpZ29MzQiL3gdV9lRDw6ENDfrQHtef4QyblG/ZtvhRdFYzDA73YewBQjNJGU+a9OPRcI
VKY4CGWnQNIe8TIhkBOXt60IJiBI4+mwDlJiVTvp7f3JJoijskbkWfgXpGY42YGuW+21K2eY9roY
RBo0WT7nR9FMzeQ8v7uOtXLh7lAu9j97YBy6/2Q/gU4hpOVCw5f5lcJ3clNC/yYwj7AR0w/69jKx
CvDqnfXeTuk40JN34HcIrzIacSzqqgBaDomfgz0A5HcT9xKFl/37ixBc4WMFpeVjJ2C18FyrwujJ
AlX3gln9nOzhp7knoKzkvfsVfZvbcbM6vqzLnVlu/SbtmkYKVcp6fb35SQxmL9+TGfvKahTWxLT4
M0BQkP5dZlrimaCv59iXQfU1FWzSX3QPKXoL6vtEamYK7zzVC7NWebdgjonHko7irJQpjUC4xIZ4
f/ypOd/vNEYshm8xpdhL7bcPN06v1UitouODVU7V5k8BoNOb1fQRNHH8D4VD2v7KNG94ZitcjXLP
gTVLyxZlQDtYv/C6fL0F35xLyQ1SBIVn0lYzLZwbvCY/qvAU1yrri0TsiOwjBGkbJGpECE+ADYRs
Jbl2tv4Qo66RpGVNXA/7FyzcVLV3ISmsz1EUwq9Po1RwCQ5xXlQ5iR+4zZvhC5HpoFxe/bwz3KOK
UvXV9At3NPdi9QGJYErSnuyMxMZbfKXMtz2wjz4DPcUu6BzPJEkxUy9yzN3qlnIWXZt01UNsnsni
GYdyU32OlbDD/DvPxVaq6gepMw/a2ePIdgLcSMCtpYbdDb1u3g0u0Ywp/uaOZBHpEJ62mrHcAwv9
BBIX0zwVuIZiUsraERoVmuPkp7lixGtMPtxnQB+z4kbVrcdxmKMhyBYFU3p7WfP8dIc8p5gpDHwi
ux1G+r4TdnJ1u37QUyb3FAXDHdS9Gzg/71NBEiGVacbZiTLZ8Z5mX56jPRZVii4bs21u1zMlM3Yi
4dTRqtzDQODXBzTfE4dMTsR2AXHlnihg4UkgQ1LYOLtoMEc4OYWAdB5ynQYxQtCCehAcWGOrKSFG
0BRae7eGTxA6OvborWS9bJ68bGGq/udYJwbGf4RzD9TqrtCtlGN6o+XkAZBgND20R2OftmVg1h/I
06zUqM/aIsC2x6BBSjfQR/4I0JJve/BPRoWGQvE032bzltpDQW+fKpwc0k8E7p2IfoROWI92/qF3
3vhGsCaupAMyFjMXUmGWdVlxbd4M2mGGHRn2Mjzw77W71goy+rFvspNAbVPH44R+5m/xjvIHjFgL
ueUtok45R+4OlTdi/0r29RPxn1vPyO2Ciuns7uBTTxg5jcWFPwCz8ir15ObAQYiuhnI8VUUuO19l
m71hhBHHqe1+D0vG9f4Uw0JEdcNsYpAUMWFmb8C2Q83q5UjWB+sS6v4j7eh/Co0iKDdobt4BmYFZ
yOtdhpjKdvJ3eGD0NI2jMBSs3W5ooIl2x53V/VZmfvSL+KlahmjZ4W8erurzyY0BZoe5trl4OpzQ
5Hm3TvYBO+PF3vYxhnJ9hntHT+NLpFk8NAy8dw7LKE0hoPyCn10n+ApOTZtqb8BP33YGckLNKXUe
SAxRQBzh9UbtcM5+S+Y4g0eHo5vZQpZ0PKFoMOTxISwUnQPvIM5ufo7dQbsoVXKVdtl5ft7m3L77
sk70s0JM79K0f8jX4XgCKIeacHYGwLCI8n79F9rcv56LPf48SQoRx0C1GMfSszwpg/3MPhe1F7pD
Ce2uDt8d8b43B4QDJz//VCW0PtG+HlJkvo5np2zHryN+n7iTtp8OeE9XXxJsao9LOyHQyw3uO8jJ
pYoBk+S6XVVaaZmUJsthtn0XXweneR5dZ7JQ0x50BSeIbbL9YMlE1tmT2X73LHpvldoL8os728zM
leU5y1pRL2z+tOWjIlvC+n8UEiinOUquOI7krgCijV+3WSRy5bv0ewck5Ap2WG98J0HTg2VDwPQd
2My73ZmqltYgn0HHu+HC95hfPG7qGj2u5y0gENAg/2f8qcnkbKSGlypdwe/EQA+33zphnlg5Ul+H
DSgwb/Y5v7I0qPdTLnYF7CThy6XXLzyCN68dRzm4cWtv1ACFFN9SDhbucWrAEW3w9o+Rqkv1uirD
j9YLS8i23KEl1MZ0rHFPXULhS0+nqVpRq0UPXocy4ku8qLItY19JhcwItKxc7oQcgItDNZMk10SS
+vkeAu/QUbe+7Zc8bcJlpzXikUZWzVOoZFU5bO+6KYYg6fK/gFD82kGDWjwcW9tl0k3PIZlKgqoD
bVzWXNkazNQLLPVlGskq//S5LwjO69UTKkUGPXjCvYhtAuXVTQm3z6eLyncBhdhR2WKJrW1AdbAm
FNAJwlG90FJ2K2UXjVk+u9m0IhTU1Hpc9vtQ4sQEKNEsZRzMvd9bkcMYbvNHWKu6vRz2vvQTZtaG
jCqbrnNxk/oc00unkNS8PqzH1vLDbnarDmiDF8net0eGvy7KKe6qpOZC/T+p9zngFL/BAq9iIgAY
ClQZ08jlbSdtH1cs6xxjcWu76gRZNdCnfltj+mICcscItELpn32w/rMwCHRUAX22pUqC2cazpxJu
VDFg9bT6yLfuYjS20DaeNlOsjslIcqRGticYG7nUwuHOX6mv8k1LW6pSSQZ0vjyTVXuuMJ4t5m/6
aHBgnlYFq2S+CGgVdx4zCp+lTpxuOtmmrpQ/XqThG5bHf09jKhNFp6UBeaZP+qQHDLk4TC9N/U1P
tgmzIK7hXbsorqSN8ckLTyn6KX2tlUADMyOSZ80nH0Cg4xeoZdvKUI7d68ZaLsyoJ92ZwHlsq8Ys
7sytie6iEHgVwqvQZ1PKT3ADFDECl+mBndo6gWAYMxF2DViYZaZ9MoeDBFDLMjRIFC4D6e4OwNCK
cJg/cXDuD16pGdKgEb+rEHvH/lGITCIcnggKpn7vaTC4m1I+lPDwcFuJf4kK+H5gjgCScjc3nW9T
F+RO3VyxyTisjFGTTYVx+b/tK94EEOUyS2YgClBImMk1OthAMOP0XIRvJIaa7bCqsRR2Kh/jdprn
kYN5lqVQzSWx8QAxd2XGNwqWx7UnsX4f7FosDEFHLzMiMp0XijxGsvPd7XpokJbr8ipTZPGNS4wl
YoXCQyQ9lY6Apqe81zW0EwX1jXNCNZX5ofieHzUwWOSqvewKHOW+HvdyN32Ig2CpOO1qXi10O9cT
SvXjdo51CML++MmAAdgA+rtVSddfhU1sclHRXl0+AbLoWuqCfLc74HyXIN3mAChrJbRkVzfSH9tW
vW2ByElglvto0iGU/lyoZqRcEUCkR2U6TPD6y2Q3eecK3m+0ieLW4y03EqAbYYURAaWEaMRw7lAy
DnMdWR05fHAa2toDu5HMTPRM2RS/t1uJeJUnxYDKcNwIcw9nqPlZ9ONDARQGMqwyXi4E5UHpfKCy
oQIU1WL9z5UmLLEC5vTxYjfo1cf+rgQUjLHj6Fi5e5Po9oQEqjx/XXMD+tgUi29OuBYXTIM+HYfx
JtX/zgMr0foNdDdTn3wW5csYWzqWsZ70kBCrnBIPqPzpgHPZpswlat3Gk+yPLc7P/RrNjfX/sxY+
ofOmjmWAYzLHYNWz89UzUHme57evloRtGyulhz9SayOfHLxJhm2IwmuKXs84ybgz3g8qxlr0+c/o
1nvVxBMsIgzzEPUPUzrbPcraUNrDZ9ICmhI63ZfXrBL4OeXrGMppLkEK9WKBUvJvd8bjq52d2rBM
2WOvVqxclmNs0Whv8aQwFffsWKpfQ38XHpeMUlOlxPO0z8feMxRO7xsZCPn9xkG+Vo/jPwMwC92w
uXYNDfReaV7Cy2r0ESsTfzSLH9igmlMFmtI8tdhC/eNBDk0agnocceJVBQcDI5fnO5d4k5IIVYmv
++habUDseo0BTNmwahTUsrQfHMECSptDivdyuJgBqURioJ5YJ3widMijxTMQktxY773MxVT8MCQI
XAgiyDMr23gqfwmDmuEY26lHiE2/PQwfFsJVIk+ni0M5O6IhXqkwMqHH8iH8KprKPIDRPTzxkzGN
TWphppPhY7S7i3jmUq3yOu+iu+5M2sQ3cAd3HEi8aErN01VC6YzWP5Zij/lJhfOH5QZ2YoW7TzE9
4kNeAQ4m5JCaJcHO9KZI3xe17+A/RQGWSuJSFFTbIzfbnSEGt+yPMJLdUAHCNVczamiU6JCMQjbm
it1/QR2w7sojVsWZzxGUbCH2NBxZtzyVVyBKvvPtRs7LUo/FnBDtJoe3sdnyIukouMIv1gyzL9+H
wSbfPB2OMTUp478KO3z8djvL8Pyu3SQTDqnBgW4K1Haebbmjn56aXBV/dEfdoLzwIfWbScyUDQ2r
C5MB6D1BnPotlxehgVy8Nt7IqbGC8h3/VX70DrD2+yDeuG9ZF4KNVGy2prLHQbGepTG+UXSSg3n5
8fSZubMyS4PhnuJ6UlltWQCYtiJ7wGTP7N8ou6vEQnq6lexz/UIAh5c9CieLC0Ppj4oIbo3PZRxW
1bQ5QBf/ubJfG0eZy7cKZOfB4LoCcegXtKkdHA4JuOej6AyPB5+EjkbvZYC4ye6WCDbgui2svn9J
UksBvoNt2ExOc8kaYqzyoLcBp5J2GJn4p0d0X+LShHPbKSq6GH9mWEObHzHhXsDVs4UvoukHCRVa
FO9v1GVGUCPP4L49FrdVKqLk6dTOdr1D/9/1obYpsRDkOQwwWWmIeDUKLPRFcP2sbHGShfeeBPLb
ZLCFU8YfuMs+ga5qRc0Me5sg9wX6lWwQv6g5qGxs0dpZszkEopu13I0KPeLhdzWxpRbsg85bhORM
p8mJhJ2uPYw5xb8YGDbVEOr/BJDjp5+yAIS793/JbtGYg0D8mYyVpRKjYGB3kCXZW5RglftPTVCF
JN+BforXMlD9uEO7JZWYpufNSCXIKlDkgSDJ+OF06qLDKGhW8e1z1eV4LAGlfGJ5ERemMhkQ7fvy
5u5JrcySloD25w4aGfDL2hEwU8qOWYgUDmIwnjRd3ey7udsZkixep9jXzn70Xrz0hXPIv/6+ChWS
pZVf1tFKYr4LsuQijsXjEC4XnzqOaKCAqWbdOEV84naFx2nlUM1ZYwCaoj8ti+MG8RA4jQMR5AgD
PGxUkRyKm++J8AOfe9dQligTHpIZHOvkAUXEQ0eqyA7IPy5Y1CdTKSGWBh+/2S+7vsQmksTEiuQm
pm6G/AqxU/ceU75wy/LZszLLbYsBTSH+VHJ42HAXnHjVqGP5Vme5GtOB1ack5TcT5Zah8kMwlxDt
yAW/ZRy/wkJm0egFdnW7F88t15ZhgN6p27GxKSezsAywPZmJ0bgyhaWRwRi/4Qpq0S9wnvF30s8S
Fs43QteL1tPLEdW3ng11NQMeVJ78f34S8MfJDBtAboelDOeyp32XcLpwJJehu9OwsKiR81QuEg+1
pft0LshZjO7YdJSq5xZjB6cnStCQ7VCwjhUbCVjIGmirI3hGtRtKHTLVl/Zmq1Z3Rb/HCSXt/YPy
TPLj7ZEZn7Lx/7qL/kfVqCqlWAPSvm/I305vK1dK9A49Z0AQf6w9sHgmcxo40DJtrOEc4DjRwLfi
EK4NIFNrD/i2JS5nQMbIYqwvqbFsfC3Q+O1/q9FrfzkQMEK6rbgQx5UUWWJbvNJhZaDaOVp7pap6
PBLQ8EZRmigfuclBOfrILKEy182Er2wDpqhjyMECR8ddHwPqB83RsSC2zTbGhaMjGGuPZvFask8h
mChJCz5vxUsPJ95iFAAdDR+OX2zXVsbHZ8VF1m+IXMdhmjvUKX6kNp9nCiD2/78vAPKoha0bICDl
MF3j0MF8GHpLsy3Neebq73E+ArO89fDux+JCNtu9tMLg2GbgcU+66rDiyiq1hIZcWIzr0JyySR2o
U/tHpMwxzIi+uilWDScLxfMRFInxcnURiNX/O3opEeYX7SCIkJxs7F482hwqL93fs4X5WPv+X+2L
dInkw4tIwIQ17yYBEkrQNAOVgRwWmO9ouw2Ac565qrTaAlNtOpKYRhZx96pA7CWmcYlhF9eiZfQp
B/zDlcqLwYvxF/7Y2L4LE6X0v/NkybkvWiJtkzfeRdVSsJc2v/vE2J8j7bO9E6zzBZ11oXRXDclP
XYVDMjoKGF+ygiKjOwBrLBw1lZdqh6RSroEwFX2DwulwJzPKpsv+jBU0/4HTvWETB+rlv6KsCVLj
iN8LXoFjTe9SLF6N3Z84Atxhb+N7TvNmfcYEE51qRGOtYE7evGaLHxipSAKLVuNiwRFQm4ynbi6+
U8M4DXHOvh5H6pAViLtFJsJQl11sBi+huXyTdPhPNQXFld3/rgNoF066hbn9xI5jWTB+GrEuJnPc
6UppoOv5cHNgLPM+IFb3P3tWPq5EPk/P59eWYwT8Ts5wpR5pi/OElkd186bynzcqKS0USMTfZHjc
nli5XKfgpc6i0B8vLcxsbPlsl+yghZgHHhK/IGq+3GbnVBI9flFTHWoLt0ZcmVNrYd04dfmoD8pW
GykRoLSWC6BHW+qcRTJChz9YShAeYp8/clr234lIjRI5HAJ54LQ/U0ZqM0ltakfwKRUy6IEvuHaV
L0nztZIWSNop4ZjfW3/Kg2+E/SRpNDl20Z+iNY7umQnFtin0R7jJ2H7e45psLw9h7hFFseeluwIT
tnnROtnk+pUpjzGkGcnXJCTzGa0FsL7V9bHQtKwTwU7CdmySl7HZJ4KMuPgIjSrwoGdBJR5pS1P5
bs5pJQsOii5XPPega+WsHnJjKtyRi4BkOg13CkXaTTSJPPFfQC69Ibnp7kwjMTAIM4TFdlTQG4nF
elwbtmJ3wgyIDFloNq/eAyLpICIeRq6S4PNHOQIgbl2O7HrAKOLchIrWA65oIxqRWVs0sXYznI1l
MWj3q61nu9s4/L8Le1UOFsfLmf4l+2jKaYrKn10M52WX/+Ge+8SCcWZCe+yYXt2VsklJ8FUb5a0a
lOO6nT4u1IK6ryoWa3CKQZW1vyuY/BnKWR5qL3dkRd3jIg2yexIaCSLalxaS4obeL9Y8rc6gsdO1
cd2mFjngMBVmB0GQE+jGm5afNqS+UaVU2S7yUzjyDYPeqqGnY919Ukg6YBOxIbcWb66gwQtAXFFa
8dtax6mEEe/m06TfZ9Aa6v7hjiwNnucD77pFNze543dXB4eN/KUx7ktvhPYKuqA2PxBfxxcYkFr+
NJW91e7ugr3Uo3udh52Rtq/UK/gnhuhcZEi3wo2Sln4gZGZlugLtI39kGf2hi2krOvK6rErUhBy4
HqN9AYunI9zKR4k+5ifaeaX+G4/BOcrNmpAxH8rAvA5wpJ/JHJR8d5ygRC0MCgeU3D0g1Bfd0pdP
uuLylAXFUaluxD1wtofdicAf6LU4xHcP9KQ4swdXFHxp0IewMGjtK9H0uhILjG6Fma2GDgQNv9po
kdLFskgHg3L8mK2TMVB4jTOauBg0fQT8gmldhzNoy4uzau7ELtMadmzYuNLHZKfCb2PPz0zUmA4U
LmPWP9ozT7Op8uou6X2cRKxGuu4Fgamu8vaHlKYeYXucKhwdl5I8gGreGxj6LIUc5nPN4hF68p7s
y1inKcPUJEGraNI7B59ZVuEHBtHv+d+cqs0QfArGkf/rXvrPtXwzMW/vLDJsOxpnAvhbaWNntv/z
NTXl/UfWe4nmwuOdDfFtuFmuWwQshtvqKXRuXosWk6dxRNc7UHtvyvb93vRgosfekRDIOazHoNQu
s5XUPsF7BIC83/Ij/APRFMqJ1NM1B7X5/IqT9HoXPX+IXVyar8be092il/835aEnpCITvArNlEp5
6QWwwAJjJHYMGeG5UqKbB/nKf0eQILNaOP7B2yQENc+YjPqPacsQ+tMI1mbDA7vomXwwrAVJUT3H
o/xKRCQgK+q7TIEq0yyy5yQkRAFQikotKTGwv+54Dr06ywKFHgIRQkbFK2mQ+F9eCCzyqSEzo4nW
77Q/rYhFonJiDaoV4jye4Nj5lmmAJBVcK7Z47YNt79Hinj0UHY61cyPLzN51AeJicoMOUGFonJ2z
DAEw0Q2jJx3j1m47JiHEjWqjRjgTDMZtZwfd2pXMFInxskL1BM8X8ouoQfBqLoqhGut/pGUGYYOn
rIiKBAnmVUQdqmoUijOG/T4/1W8rfQQfFRPjV/mtu3jDC0ZQt9ktS2cS71O2LxOYpblDNoAqm2x/
GUkp3Fd81KtCeehULG3p59esE/pe9/yeJods2oDqF/I7v+zmaOZcjjeYhMz1w1DrDbq9wWnArjdp
iADLFUEpN0AF/tYv4L4lpQiF3ZYeZcSv+DxXsqmJVe/ss8/FmppZZYAGPmVCJ7Po47a55yrH2A2L
9OzZ/uHqsfwcLPocMAotvmSg8qVEGCNNb6eijUQQeQCqf4QQCtQrkm4g+mw30fO5lNPtwp+GcEsJ
JtWUiendPFvSqe3HZhjDvVdtJ1CZ+eCd3/p3VtVwIzF+IoLLcSr/z5JWMzLej+wh5WDdn258FPX2
0Rz3mBGCsA+KZoKzVPtzBaspw0JEPJCTqmfVfDQepbWAdmYIGymLWrTQGENrNSeX+UY7TvPzMFOM
ert/ojB4f6lIWZUbit8jrwkqMtGoNT4k08spJCnB5gq3oZZo9ml0oYYMOYqeMycwHd67bDECq94Y
y64IpLuRZmJV5A6EhMZjchO6dCT1xIrKmsGmRQ2oyXJOBLGM4AlSniOmxPqQJQhOs5jaLD1QjF8K
mCbc3OlPCMGYCTDT0G9+v4avGpJL5KhEoMbLehM1zRQFvEdXL9KblBlcjD001Qoa8dHDb1YGJnm4
q3qzlVF89e1Pa/ujfhwxSNt4SfA4NF/ROSF/5+A9dwns/+N1LMmAUICvzhVGPzMszKy9BRyNTmU8
FHGbZJEc9lnv1O4eLTnQIs5F/I5hJAdtetUAjJHBRjJpXxhpOGmcyZ2/bcj6I/vo1xzMOY9Lrwe0
KM+Amt6QajXSOmDPAl6TTh+4KZU16TXOVNVqMPNeMNZ1rYZqQS7Pf4qTML9pt+kh7e+nYN5qGmJq
ezbHSMdh6JliKgTcB0Qva4r7P1PFAeJOcMuwlEIVnZgXBwFDlx3OmrFxws9VRVfi29hEtJlU+5B8
BOYKH9uGa3I7QKZrxeZ8I8IIFBeApM7y45dyCk928dc4lcr5yEFdpc3oogeFkH7qagAUWCv3eNB9
4le6P1/13WoHBYSW+jqb6GYDNDqiLRsxoLFnVk6G/OD88z4Dq1Gp1pEG6Rw8QcLCfIFRBvi0EHM/
LLmG8xVKwJ7wuyWD9UWXzW8KjBjoKswHwRE5ivJQtRvVDdWeo4ZmM4ZKdkN7MmWxf0to2Jhcf68J
9FohTBw47gFt9eaBQWzWm6SPB50FnQx0fGRHVsf/KsU8BXpzfK5K2eAX+8ATpqgtvgWBLKmIvgW4
AtyVha2t8U36yTyJNi2t6SgDXcJg7vYvj0jXzvCIIe6A9WoKglh+my9CcAJSJf5d1AdalFXFX5Cz
Sztw2mZcYNTpxMaJxGrEKxgGLvifpsLtT4FI25G/udiBqjSYXJitcSndL6IpJQzTO69k3cb99SoM
UMKwK+4A7EiVVkJnn4Fa0uzzotGN0ojCTNh61zlRV6wuqq64v/9loFz2sVZm+1Oql8Mf51C8TgFW
UZ9gbGKUiW/vH8GpMzDkrFqd+1rmnBnEV0iPQzetwyCPbnkL4/zRsQZU5XrP1GFEZi631VAJYgfx
sF9kwTWrAkjGmZej9DUp4rnVkjaZdnSArSiSumRAzFsC3U7UgatYod1fVdAcMBUl7Y2/9eAKGpht
vs+9ZxcLaAcSac2U5DihDfgS9qZSc/xeTU2PUGGDd7VEgnlpM+qN4Yb6Cotf/MvaUjbDs93ymPj7
EnE8kAEJF3QnSTFDc/GiKV+o95tMMu9Oa4sPSKZ/2UlmCj2NNEq16EyW4PncOmVIHk/Wb8kJD1b4
5hJpciLhG9VOHXNoBT8AtlEmG0QevEs7NgCQvDuSeW+0B1/z+4Y2hBMNH5g4+hhAwuxm7C9Pq1cU
OYDyZT4KU+TDcouGlcgqa8VQd6ATrPcFGr0xLd+V/BURa23qToIqHNzWQpERogSzb9RNIM63pruq
+CiIuS2Jbu4fl/BHvxwWv6UDPGtaSCRJ+x5dHRGJXKX/SmENJvjYC8iCHEgKJmHeu5Dv84NNcN/j
Hh8png9bIUf3RakenHURvaZ/qCllHpWXYyBwnD3SFO6xvgyjpCgg4RCxnDLWIV88zToIvuvnaMaq
EUKthQGWlTq7Q3MSgyo0g9URFe9/kH77MomECDvtmbT4rVisIUcWIAnchRHqmEsIn7ZfaC/aLetB
StFrjj2auiTAXtIxVhXNkk2B6645lP6w6AO0Y6lADwRRzH7OuiqS441G6axG8jhS3kQbzFlWTPq9
FLqaTIEwkrXa/DW3xzuTrv2CAcdb96I8YJ2gm5SW0bMnCfD7oIEHQ/oIKLcsLdZqOqn/0hr8RKLC
o9Onpn58rrBVg7UOm1D2ZCXVcLne5DBbBs5QVpvsDGB92v9GRkCVy5aAgOUA130GrHYqKXg+sm+V
EqWWhrs3lOsLmGnAmkc8bGmhWpt1vXrxWFX0pewz5fBTT3YwHTa9bFiznmhXXLc5RKawqeOXARC0
ZvTYAOVA7WkhTmiRHpiWBJnbXCXKq/BlOxHtk7Pr35nX46gt+JJdhYJFkFohJ/m/WJYrAbfc7ol/
2I9V/EtoILvHz6Fm3PrRzn4SwztknC/ergd88mAM5iRzRkvMqCAZFKQKgwePI+xizzbw44Ckn5Y5
5OtA8Iw/sDtnS2gmRNym8NjvG6LIQPY0AtdJ+d7R93FAffQ2VRo557lfeScIm5/lNSpJP+1XjZUP
XI/seRPhLJiRehpsmlcPIuF3w6yROfqCcYSCYY013vM++GGfLx+Axf9w/w/o8VNFFMNs3n6/cb+s
7sXrW0RWjko+zYc5+FwPzTdKxrbzXsvkMJCY2Y2Yj3uXZimyvXJaqTBWRXsIQbwn2aV96+3skyrM
pguKTTYJkA6DWlFWqNrXK+TPdwGdaj21kTKSt46mPJZJ4Vx7Wf7nsR9wFZCCI5DUcmRcZm6nHTQ4
WqkZ5ioz9FXWXvlxc0gyAoWOBOqjrXv+qUPDmHYLTT90b85NIT+aWzfBUCqykVh2oTMkM3Ap1LXW
PSJ9Wj+VNktJsSqdA/kpnAUnQu9+oYx3EKYYDpQrQpydcdNUEAQaMGIVuVaTL/+P7iSg35kxjsjv
ggQfGT6DsYEmPADp/pDjBgZYj724LUxkQlXpM7ZbgmZbBU3oyca2oC8TUkDhefvGADnlddiybJLX
6nMJ2GmeQ/HSYUwVfishclRC2XvJt4VTsmCbnFE2RimTIbEcb54XRbQxO4yknfFwUQqgz2znDF5Z
0Y6eHfoVdScO+2XgJWtlzp1oLx0MXyR9UERqhOJJegRYpb+sck1bgYEeGuVIcxfu7ODTuLbCMMFy
92nf2mIv+S5RDgZHlTGEcz+hKMuC1oEePyFwKK4eEXZSs9LiuU7caID7EPuzWTLSHNzMT6gQqqqH
dKDHWkfV03ZvYDtKP8VorfL452DapI0cHCM9IMSc0iYvKi6rqsSXSAY7Pd+7Ap06I/j+OrlsuNTe
qkJyRtkDI3q4NMdSIpU2rrrtaC7wXwj9vGmCMROYdDDYqebjNbc8GFUObn4o9Eek+E+/XkFXAM8j
o/1T/B1PukHQl+ELZ2G277zPjE8wcFTyN2uoic8jjXTOpclQMm0n00eg2o3SX22yxy7pIRP8sjtS
ASLqPwk99iWuHH3mGfNrg7sZ8ir5kf8O+cp4ixwSOTZ/BEMNBi6GMX2wnS1aR/XfgbTDMh32GtTm
I7PMDbk3X8k8bDUG0VUSmhLAPPvCoPIXOCgNRChioMvjAxECIosTYsAVdnSyyAKEkgG5NeV1tik9
V6IjA6T19Fpg+dqFBI2QZDJx7bAQck7edMvUW9DG+8McDgVX9wPLZdhBeY79TpXavewlmwF/e3VC
CUED7gdXy/pWKVHRTQtNK0JyYHD44eqf6z7V6Mhq0Zq+hTmfURraKfP91az+F4fndw2/6fbPa0RL
xIt9KpYgaxKl9DRT4fIhZtVrpg0XgXSQqbn6Bi/OejAVGjex+bcSquyhri4ZdLmtsZnfqEcLhmya
joPCPUsTpfnI/c22gMoT3KtQGZM0nv2gPw2i9/Elou1qedObrFC5LseK519IIlrRiSIY1L9fe1oo
OJqr0HSEfkHUCpHKhdV94EQdITfCt0VElqMg/myWur+4xL+yrxSHQyWCkE+Vto3RYhJBa985NR/t
3ookojynZzop2pTJu9f9XlEVEvXvbovIFR9ZdbML6lArjRvpGB6EXiNBTTvkB2nCaUkLTFJ6gMZF
BHuEEieSKialwybsN6d9Am84cpNvxNfs8SQlCa2qG6xy4DubNmta3pUJRrse5UYxuWtG6+o3okgM
tIGc1LeMkLUKlDgXcikzPPJSgV2Pqzn0beeDCmffCL+mp3fXI5sYklcRNJzCROSRkpszbRxhrlhH
PT/ArRzKtOmE5qnnuNaVU3SW10KO2SWhUUCgPDkwvCSOzEW7YImI9pJfWJ9jCOEAyaoDytCTQVhZ
nuDYr6DcpfsR410vEXgxyGGNsqjUBdq8wJs/Pruxhv6GRjMhUikEVhu8TkP+IEjzLODqntbdF8vP
0qjUYm6ZqNACneYbDG4k3g/k9nhSuNMGeHL5N82hhyRHTDyTu4g8nKeqTyKvfQ++d2BZYY2FC0uJ
nwTydrVmh29ig+0RhLTCVLcrxoWWMzJrlN6bie2v+3WUFzngr7/4cx/V1CqQwABqyndP5pg4HcsQ
GpBFcrXL+J/scZCxAcKHcR96FRJBBazYHmskPFk0EnxSvnUwJTILFhM5ruPbgQcwVjMSmjDJmxWW
HOtizerha+jQ4CRL3EoLIDhDKpTcOkuV8PP9xkLLgiqn7PGY9Z+SXGOWfnG+6oGsjIzznklh3VBB
n+/Su3d7W/ExqL8dcwTgPoo6eJWnLuvFaSYQ4Hg8C/BxosB8Z173/Y48H9KBNSPdHQbDl/cHQIoz
2kNMUkk7sNPm9h4UjKCqtlYeESl/XDNP0gLSZWBpJ6gbT86rQk7XrVOfeJ96xEAHrtwWITF6/lIi
i+q2M20pX80OyomnRsn0T1nQ0r3NC55pEq2H/IY32+UOo9Ab5Q4yExsIPzNOgMRla3qnULOxnwPo
22wkUvdlgzgBYAE78RdAYAKmGDH7bcAwMUDzv2YzxqTFsfLWMdXhWMo0M56GYJFEZKhOqsGB0ESs
StAVruLo4F7rlyTRWFJXv9e+vw9YlZ266yWeMRNnlIhZKtBDfMzV4xxLfS1A+8R1jAZDP/OZZWbQ
RgC5ViBkoY4XW83EpztPnGJ7PYc7dFkdP4j7dd05/Nt7i0RuIrJuT9KWsXPKwcWDyf6KZfVVUAIh
dKxh0wJjYRWpYLS9vK9GhKSqvt9PJvlTtNqg3gnH29eGEw6QhGoubteq9vvGv4AIaPr9v0hJbbCH
EFwxSXOtip3CUvGF9qwl6SC+pTtBzQ4F94qStjxHUsT5LcPRAcSFoCl7No23o1E+3a49JgFB/R7Q
s5F9RdgB85pdqX+NEYv2ulSLqxZd/Nj56YaVO2mrRfIqzkVs0IjjB0bo9kg9WlbEVNg069xXfn+a
FcKhfZ+fkSy6kp79kojgjXXim9uKjL1XZiVOj+dDlhRYGAX2Z9M2clctvt4Zka5U7XLV5SD+ArL8
iLD3M6rtHfoaBNYdgPo739xtax+x962YCu6Pkb+7I4gCoi6+aZMV6WBL2/JyraPot1/e8bGk4EfZ
NnBnOiWAbWDb0uF2zqdsAVdjrfjeExRBkpbX9WfUXkfUwLoWIrSYjZIm3ZDXwlnaOyMtG5w1j5xf
Wx0J220YAFdk8BmIh+LB76rZAFT7H1O3ySRCUYXPQZ2vRAQ+YGVhWFYHS4soohE7me/QuJQG/Ihn
NeI5iBiJXEr+k90Zb3pZMnQ6seo8euA04XeyFAg0ma41yoKUJC5HzwdueBir7z7DA121vCmwfHxB
QTLLhIl7xOzdUsqo8bKwDPitLRoMElXBOl7YqScx8tUSO664cQak1Ex/pIaQGipmV2qyTFy5jCX2
RCBmOXFC42HJHrZMglIHMqeflAUI+ki3fSMSvtVLz1nh12UkVvtNB59HEwbgjLRsF/avB3UJkzC3
sbXPF18wRWqZiA1Q9YstSjsbwDq6sgC0Vsl41wbXu8u4X0sR0xTOjJaMiEIUHRBPjcc+ji11GBL+
gfL6OUcQwCD4XN54Wj0j5qP6ZHZlXRnk2sBxgYItVFUKE7pebS9+YPpTY3PNlNnHEYsULjpTQ/Xu
EDoGiXkvsYZ7hSKNpIufCBRQ4gL4BWoQVuyHM7AC+z5seGp6JzS3tbH0ckyMg6OkO/h1lIin2KH4
DUVtXpYxh0Tlo7PF08ct5TXLVyF44s5pFlzoGlsBHC9gHZol/+oIkcsFJ/XIxiOyydeFU1fQuE8k
/4+avLp8XIGH4G5eT8Yx7TozAblS+vatvhOVbjxzWTagp4KnVVKjp6ecM3/BkKs1M9dhcciBPyEd
IOfFdbeX4ntfKybiRS/D0rOnvPcv/nYD26Pjmj7XZp4i0BzydwtXYpbPZpPNVSmoW/qesXA8lBIf
2DxIUXKbhlJcQ85G0SUfq/O6gEZD1HcMWwsFgPPp5iV139dkV/7cIuhAIXDO0kYUzufe7CcgkXTJ
LJykxDUkUIL788IlK8D0pfNLrZyZnABuLRrb8UkNiY4BAlTbnBSGYpGeWrXnvbpVHuIuClxLJDMV
Hvzl1ZUXttvGWGML7g4usZSma74tzlNRrp4nLCCConvXY0GTHuQ49QAQvviiO7b0Ba5av1hGGNCp
k/qMqEzwR23Mu8AD7PweabkgT+aIoeOdh8QdaeGRDOtz3yAQEEUBB88cTPans+k762TOw80xOidP
RzOf7iF3GS7pHMpx5bc6OlA0ZICqUeZV4sR/vpBbYHi0oNTG9QPWFCkJFWxin1H7q9VIXkUZpYiB
n/Vn428BHBcVF+q9LuoMQ0TOSghxuLa0TgQrzK0qgkr7T5kDp1m7892lklwQjBThf04Kq6C7t+6p
zBeal2OUh5Buze99iPlDDDrcnfPTKVjzqOAcmDUokOUw4g3cmhau0NBs7AdXYAYSXzxuKyUkGmXX
8AouQh/lpj5MDpHxg/QNbe/v/a8xQszVwSdKulLhfc/5yBYodR5XFq70DKqQDMEdYsrMWnmFh0cK
U0mNvs5Yh9qJEaZTWCnrEUBXR9P9a6H8aLf8/rnhGiXG9IsiUqRdliWZ/5GAOHnt01JhPYduH7hJ
VKxqwKLZdhTpl7MxOjxnpr3QCkvM9wed7E5rzu2HQtNwrq/5BbznWQ8eRBdhRB+28VuhRquRrUev
M8b7urJRvKzxVWzGTU+t+8OQoh7SFPKG1Z+D4yxrz/ltsxUpWZF4EiTMTAiS2W8oWF7PLOn5mdUW
KZzxLo27P+ceeQ0IYG6FKOctimCkohFPaPk8CqQcE7/IpCPy66loIBOtRD83pEH+zeKVyepguY6C
JWyaACzxB8IfloeEDrR9kBTYVFDKlYmlXCS1XDOiVZz5jWlTaSsR4cNIbuQwlH3bclT5tZ6XhINr
L+HqLNjJBRgnRW25B6d8vierNJFD3FuQyb+a8oLManE1bPZBmsn+PgfU+oR+nTCOPUG/cNspNa9y
OLMaFS/kpCeGyODd59mnmqJJXYt2QJMr9XOLA6KRzQbGhnMPkLspIVD+qadXlZaUq7KD/yjPi77i
F7A2rbwfPwEN7oHcrR5eMPi4m35BoWxRPhLTvY5FxILDcHTloE/JghmOupheYrP2uXRW2uaR9G+6
vPAPrvj3dfuLL8ajKP0YiYoPr+x5FsLh9EnGQ63siCiXxO+4RscpBkMQ2T6yTVLxYHTIG6orTNeu
pznGVg/zz0e7VIOtGSYBH5HYttRu93P+CF7UydZ/keEaxeHYw+yCA/aiGrRb9vzn0UR6kEMKUTOb
56PlYIrLm6Pe5pfdSFZnVYN8lz5CLhvn/Z5ryiqorwfVdl7Ub/fYtjVezjqugrLBTPOMrkxfmHMB
AdaANpDz9SwYyvrQF/W9C5AgItG6QWBst5BmwkWZem5T19qiLf+RfERw0I8LY2eG1JsaRsyYxD3Z
1x9eZDev8gBA0mkrj+Z33HmE0Ck/ca0ExC3TStZd9YFx1/u/3DSvSJ1q21xudXbGtuBox+zxjTf6
pSDnZocGVMkcIjZq2vBSPlW9+/t7CvoHFKMrjDj5v5c6b0QA+whO5KLgs9imYGxExbID5J+HgUu5
dBFoFfPOH5EvfbKLi9JofcdceV63Bf2vTLROHyc/F6labkrTdTZKb5D3aobQzS+8gRbW872aIgYU
9ra40gMBxwaRWQYUtPiE13pB2Ugq7J8sEe+M5pELxuUIRap1OhEF05MmjqGm3hkmkio6pnnGUkBs
hHOdy+8ldDcp2bswhWML01GNJymftg9avOxpsXdqRmpnBG5mYti+NFvhNnLh451BHsC09eSrPNxd
9F9/sOyGMxuuut/FpeMNIaUswpur/TqscNMNOlk8hXiwrfNyywSHmQkxk3Ga8ojlaufN/dAnIGAp
FRmHR1cC0nrIBAg3tG9jue7JDJ63FepCMQUDH1Je1KQI2X+NyX6XJ/nJwrtpmR7GKoq8UpeE2pZJ
ashPJQdWTRZNFliOZS8P0sZRrTa7Xju5zdKNgV+rMBPj2+mmk/AEVzmicOPC/p+Mf/3GqJTJqYnP
jIfQ2XawYLwBXmTpBz0rlC48i4ETyI3jB/Q7iL5a9/XMRWvz3mdV1Kxj7zrPUvItAgmgCLxX9mh2
vxh/PvKhuDb3x841X12KNzbckJ1dg56CJ4WYcBM4xwMEclOdhi7DoksWaKu7PCXf4agtyoVeFyw+
VxW5uFWS9LTcjLo6zwjJEm9RPkCRFsnRM8hHdQXjeoXCwBiSuZLxO8vgDKzn97MilpaSP+gXYWKK
m1BvwOfGUjM3fFo4SsalEzvlLOgGRzwHSvmM4jEy8sqGWKu9Fity7SMv6zIKvMzhQqe+Sjme1/a2
lgWer5ocJZqaWu9hoYVnHo6Pf166gW1KrORoGsaHE6NLnqWC4UTXnpFa+2fioLYB71BRdrtwiNed
0VYhKqVm3VPRvzogWTDR6YZyjxikdTVXC/Jj33XZ38joDcmutFw/af/St88D9v6LqlcifBlxhvPz
sT6VHePf5oxAkmXbo//fedJE4/u1BtN0RVONOb0UUOBW9x+4AEbQ64tyD52mahOnes42j6/EEcsC
7YFHMvl66hFIxlCAka/QVJLU7175H01umqM7y1jcX8r+EH9dxe6HXYyBhlSVifGk9Ztt2cx4ZB4q
lSnVDQ81o+Z25HbWFbP48UyD6YM9fr2rVQKgBThADdnLm3LkyjaBZbdWNluqsLKYuvwqvmFQLmhX
qD5zdam5Td7sscdLAajhIb3GcelAis0TJ3YHGV+4KlR6dpSIIpVCDkirU+mrL8EK69MXQYpEYLEi
OWF0LZc5sqikK6EI84dQvMDDqufuhT+9FXi7eoTHV0sScQWMpDkAb1piSf3zzlsBkbNT9wo8B3Mk
4QZaqZrxS5dA5LDJExdqnWgOAURIkF/bgPt5PXo4Tq5JA4tHajoanmfj2sKkLQEwtz0qohLbJBCy
yCxdZuWUnvJ4kFfVM7P4kT/m6osPpPgbekn2jbMmhw91uEm/QDDATW9F+MkJKB4DTVQReIDd8YNy
ElkRnErFZXZpQd6R6Hpif/OTheYr27Wv3ARr8/lMUFNM8tcUlGZ5sIKD4ZFoEllCO4Hx/4kWGeLR
YKkrmmq/cKxWQUJuRP33E+Ff0E1wphNn6Als7C22a27FdNB8uzZmULqB4+sB67Wh3eYzhC+ZrX7U
IyHFYNMk/XzztPZpizBr7iQUg6cUyiDkFvATU8CM1y0J5ZWsFZiufLviRR9LNHRh6W+SaX/Czn/8
g8F/c03Ztx2VEakAjQfQoKY1Np729wDwjy9v0zbJzkE6J8QTjXl++h1bsRWwoac2K+14NoK8/FVU
tXT06VT0lKWoPL8/xL6U1H/O3GXTeFPyQcPPsXTjA7ImnW4IMokfhzveeEfwPj9yCazR7GWuBDHF
caJQ+SfqVKLTZtwP4ta7LmNgyYL9Q3mNVXcCwNGMe6DdUffUvmMEUcqvIGBgmH/qfnSddN+lXtTi
/iyL51fjysOnMnJdBztLJwcl5ovLyBOKGjntoMoEPC4G4ERRUYiLKY6vY1iU+TpO1Wi57Wj0YYt1
ZhWB6a8xfwM9NJQLFLLigN1FwoXga8Qi2qPmRLNHhCjq1NY0E91BRry7UgpekqFtDIS5LQIM+gTF
FsRDb2OaHj490Ca3U9vook/d26haqwtj4LtFNR7Kf+7XMHKpYpLm2MRVd/uNJSYhi7qSv9A6h8zX
RYPeUbymM7EPgtz/upQrgc0eKyIDVeoUn7H73rvmB85wwhe+6yr20G6AqICFfOxBzDXA2Bm5r9UB
ElPzIrtgIyDBoH+CvByGjm6DFbIq4qAxbZam1Try5jbNwcOIIx0IH9L+9XjLaUP5UrtXFmoJmtc6
+r8/e+00N1b48RBxmYm9pvq1mcYX7STQs+0PlXnbtypt2HhfXsgNDKlX8H/pIxRQAnfac6FkiN99
8vYomvOHy5vXIVaYtI4wbO6PHKzTcEvMHU7p1wMdU02hVNLKXUmbzlVfpb+j4ad0xxwx6eQOYIIX
DcDKqoZHS9tDGXua32WYyRSsr4zws2d0AYtf36+lM6YI8JByGEngV6GyDOua86uRjGU494aSppkN
yAflwghEHLjXXDGZRxofm8QVoPURSHLreh8sbpuQxBHBf2D0ZOGw4jynFrkgUwM+h0b3f42dSDV/
d2SnOKLyh9/d16Q7XZmubF5MJeU7fhNaCjIMZT9YAVNt6v5JsyHwaLXjem8AY9nak2oCCXNXOtvu
0z7TwbxQXakDiX8FHbP5Q0pxmZTIq/ii41nwxWRMvyUhCtGAhN6x7tjTuTOUIOvLHgRORHXqH8q2
IvMV0CtUOg1iyrHgYTKgSEmnS6EcpO6pLNWZnUEcvJSZqbABZ+B2RMvqcQ535StWJCf5ja+sVRyy
M5FkgZvY4F1Wd+YMTcqSjza9i27xGvmpEHVjVajEr0A0gvYqIT2PwMjXG8hvAyDeOsQHNd0ojW4D
F2I/+w4cW9U+DiDNNUHrxeEqUagBdo11v+2jovZQpg3EHW00F4WvM4xcIS/hbItpyYYSLZk+qaL6
OMYjDDAQ4m59r9xNRzuaNXfNwEt1ztTLP0P1Audael5bE7ADPs30OZb9q+J9BxmDdLglAqdXhGd9
VBOYiKJzXKbpDPY4QrwpKOoLOOWFTpW+Us8gc/pqBUdpsvBCR8cO+GdlcC/j2uWyiMy+c4j0ltdZ
/ACh1BFw4+mQWX5lIhPme1Aq4m0WBPOjQq0RaXNlMB6JKyi73ZaYgMw0/yO0oKXJJgOF53serisN
fwxThImMohhrKG6O1Sm7o4ZZH3UC7KRP4PqmLlx+DZmuMWCgX5hVD0PnwOZb/ThnyXiELsoHV84Z
LEH6zV+fhxotSFAhYpyKXvymBnFCxUqw/JZOsrzvUrO7Wq04i/XlTzvGx7EG79Sgj0IUPUPFEbEh
UuNev2xUTAigfOzxbIahylmdHJObn+Ej3GDZ6c9Td+OriQrY1ZG2HfYsywKPKkqZWQ2JAU0gd0RM
hVd9pcvZoWBANtWXng0nH4WeC7L+4Bb/69ivYRIzaPQuATb404ygl6f2yKTbMwNtASoVdu2GOjj7
yuN7A/Swc0DlicRSka+63P53nY8V5UTKIDk8eyxa+TzWVGvu+ghzC6tEf17WsGFJzIjAfuVJRkuO
AlHlTcUwnGfdoehliQ2zE0owPwDIIxxP6r7zBvkd9B9ZWPI/bXw5DgEjcpU5kBJZ7X6y0HMkeLhL
Q4UoBMbYPZVWlmIQfQPAE0nqrc8m82Qet88kMH+uJYyTGQKwt629a6SWuv/BYqbxw/H7y1zhtGer
7RNe4GXaIfkhYgxJoHGeItsBmdq2LMpeNxy0q2XmI1iCC5Wrim/oyvESR+Wchw0y73FpWNTxOIIl
jj0F0HTBpauY/EAbAMXgePr/yQ2CvjwOqJsoZkwgF9gXN0GTG1d1vANpnvZWn+5XdWhuXJTkOBbR
6rynAcBdAiokNCT1k07ahNM5TK+kFcmPfp6QAMJzMfpVcoIF1fmT1oLvJgYFlbu+T7G0KVxjM2Zd
DJoxzCs1TK7KVZpqZEJUphwTeoV57+wIuCEB5gtDoLiKVpvsqQfM2Xp3eEvNcyxYp2iX/4uFixko
3z30H/CNdQMH+tNr8842QRJmIRL6KoogAcUacqzU87pYjAVU4yiznxdyBvmltUBmP0qPw7FlnACN
Xbddk+RMlD0boQHEquxdRej/NzmnblkLMue6JqLfAq9VG9WFYald2vu97zQmvJT+B+FkXHHQ+yi3
XNa9UtQkwPcmH2QTyYUAkx40ox7lwqoKjgFqStJiKZ0GN0cx2jXt2lnXQBxg8GVkQjcFWAOg3eis
wTh7WFavsSrTlQPv4zhXlBj3grKp/v/huu1jxbtVfcWdJ4IkyJCDNl9puC9Z/tV0Ji6fGL83TSCh
Z9PgmtghrtejTj7yt9sev3JJP5bDlJuh1ZA8nsadM9Q3GjbAR64HBsJHL3tJRTuRaHubVA4dZPps
DTBSrv7kioUTiR8+7Op/AnceT65Ur9tsPG2RwAjpOlmwZ+OKYUyFfmF3n+b7uw7YUJBqUMxTIECQ
Oi6vAvSuIMmhBLD5zPzwkS0CHmRSwa/j4YFt9kqcOFNrxG/YWNt+90XSTHBJNrdtTbiJnbot+p9m
2iJBJN7xFgDsI73iXmp44C080pqp5Gah2NaXr8bK07ovdOKD+lJS10SFJFKjDdyarNIo0xTNOuN/
BCf8Dn8R3C+ToJ1T41zEr9+RWbCc8VecVzVIDfc4W9PAgthFf7IWTZ1TqJekDUtWymQXYpjgpbOo
8xFuWSdmT/svl6YRLN83apVpe9dCry6OSRUb1y4jmdkZ5PoKjDd+oh38HmP65FRUNmmYKZkKVTMk
9xQcJGDqQXqncd7duC4qL4MEhka0XhWhdgXU1KdL/ANznzmNMhQgxi7Ltq8JJ1UdRmpUIX9R/1o7
aNl+Uvz/KGyTOkKsaJLwNg+wP9JI6royyuAw9BNzpLEZJmsbs+CXjbQ8v25/rDIYwjoZZjELziIN
cdZB6v9kP/TqtcFncbNNdLJBOudyPuBPsqk0QUGDHceVxFVhVUYZlZ4lHmJxs+DiSj0aiYswFEMU
H0CwE9oJ4ViShSpNWPdLJYVh5Zu2+4HRqVmYuannsNF4F0XynAZA1n3Ccte0s5VTnOqMdID2/OGC
frqqOcES/ahxx/kyWarI/jfZsnZjcFd4kAlqs9xioCQNSF8rR7A7rh7PQE3+1AEGUc71mRcMHnPE
dhzLLCBbohZjWFc5B+rNCDgJOV1CIDbA/fm9NMIsiLkjc4aIgGa/txF0FI2wwS77kZgjwAMCg6Da
SYCAkt9g2ANtVID4mVNO4+nbOM/tmA1MWiP3jtx1/9DatD/hX6XfFcGpNA16blq8A9Xxg/i+CcZV
CawV/JdMgB6lf6krtlbYWndFJr2K/C8Vj23ypDHvoGCJLABx2Ym55DLM9m9XwK6fGT37fjIKS6Km
56jmKl3Bk7P8dtbHIYPptLAedfsZEkuXoHHhQCjE5o0eepwfID2T2zCJMW/Gc/tuEESkJC6jEii2
Cp1F/VQ1NRcNO99/gnbRI4hbcGKNZ/0mUDhr0rckSoWbBr5aVVmJ6q+2qXyR6pf4ZV+5+Zm2LQUv
skvsS1OtKqRl95TUa1HZ0Topm4ZCQufS69VLWE+DE39/sm+CBLl06nuEx4MFYyw40KH+G17SzSAQ
SUzxjLv8Hn4+OJwljtTEQi2SXsZaLyFLdYoIFSlCV+WFRIZwOPqz5JzwKhDcJAZxUu0niUE3YnYv
C3BetRzowGXhWEbgnD0skwRwDoDBcV5gBSoh4e0si3ZTIZ0mcbe0tlY6mxO9tNbleJ7ARzT0PPjy
fqYvWntrUtnRlbE6icq0FLEEq4OraHNeqY6cQURRWhjt2OFnb/xhrmwDAmjPYFOqxeqcAYflZGBq
nV2lL8hHZFe97gVIGHVH69NGSQphdjpxMD5J5i6gE/AkGwWqIV76JZ80E8CB72OCZLGP35oCaoTI
V7ahNNWqB0eAZiAxb7Zh2D1Y8NQF2UjTv3rFTuuBynAg1xBzK69cwu4sbGNhQNwOCY43xTHjWqkt
iLLkIRXCihuBeDoslNiLgutqxqZsm8hZaSrEs85fU+MpN9Q3QkbN3zOoCij9+6JWbx99Xtuz5sEZ
7SBa8Rj/NHHN6fM32O4HsG73iUaQVET/5WvOBXRii3SGqf96sXVD7w73apoBHSb1jm1rqGYawhaf
qxY6Gr7TqxAHNathuoZPjgIt12xC2mE29TGGxj1/uTWEtr4raG9N4+WH+jjeB+BhWtfdkJXormu/
eS9qB4rN3VF5OFiixBMdJtA0nRVj8stYU8cS8qySPoK7GUjlpEBksSg9k1VL9d2QxvSh8tgGZvHy
tZW0RC+Caaq3Mi4rRsYncRtBbKHmWuv++Ngny1F8wNhpHV+OKaE5x/xBf08oUt9GJEN/vcg6ATHA
r0vmdeHBy7manCAWMm/Ewd2PJQzrbi9C4pImX8OeFfazoLRxqhxaNL4PtIggVzubeg+VLijPEoup
kRCl5OEWGJDNpdzWwO17/srP6siz0vwER+1or581CpOwHUoU7xUbP826h8S3DGfPjRbHw1ujY1Su
7VxoeQvSt0TGckXxOIOvqZzNV3fmyqOIm9jBaFNqtKxq8B5biCnKCpV34RDRLayeGjPiYBe/fJAL
sV0LjoEFGnhCAB5vZ/CTQdgyX4sSkvc+zJjy1M0d62L0piKrnqAORfFejKuYrcNYOqWQb0mo33yD
co5kwf0vdNKmQMykWuTPT71RKnqZdguO2e5BnbnbgUA2Si5FfrqV1+letF4iu6pAIZqQb1I7vtN9
MOF1rVyWvrsyBALRw0wy3IG9JXLQqNp9EI5GwEZOM8WB2GWDBtJVM0h7O6UVUtqH4BrF9CIt3MKH
Hn5DPZ9HHwkljZvCS7CPn9pG3Q0wgSvSLuTxWHaOrC5egFQEL3e0mhGmbsRFzZhhOM5SBHqWgcNU
rO+XRa9hCKpV/ePRBNIyIBO5s6I138Fi2gE7Kr8vQ5s8w5Zh81bbrgmXlzsq1+6O9lU25Y5WfrBC
wlZ0QLyYVFhuzacF1mDeoNS14coVLks2FrO39rnr2qtvNHyNvmpFuyPPTEOxQIJKrAE80I+ZcJGi
UdjsyjPHA+4Z2j94t208GGooq2oQJVePLJsgMw8gvp1gd3oLALYVWJG6xvQ7zmzFdEijeml5wHBi
S0LvLRTH5RYWf4x40iHlWZwvAhynliADL4rrxdMFQaR1mosIsn4nQ7k/47JYHXTiy/pHe4/2mt+H
4JgmyqEZAAwzRS/g8gv2EYbq7uHb+oOP4BhKk7OFyV/R54cFteWiSx9EYpyggZiAY68Y3mTSzyoO
/NFOGnemhPwVQVe0nWQgFQlyrUuRZph1WKGYeS/wBC06IkQx6s3YhRectuks/TWIRAhvDZf5N/on
RKXBu+gaR0jLqdwudPIxByiK+xtcYvJtSGW5x30ReLSRRZeKMPF6+c3TdISVw36rMMnO6x5qzpvc
KZOOi5jyqipGDNRcZQVqdmQAz1MHAmwSb1EKPjqyOhg83qd76IjJkKErmRWCHCznKZs+RPgrj/TT
oIweLLbMmXcc1p72+bzjLzdQBDpHpIsy84rdVFfj3tAsCXPvf/rbuEuFktAcJxzN/Y8v33978tha
9GK4G6np49uz6HM6TBicIK2J/oROFI+X8L0QoIva5U82B3mnvESeaFqFXfpuUcaQ7vqGVgeRCZsl
3n7dYm/dzByHM9lg4CflOEmST4NbJB/XJMWL+p1c9zNBdQcYw9YMZh4QSQ689VnwRu7PBJHbgnkv
jxO8HeCud+KjfXH+MWbghzBSdubgQU5bwqozXNGYWPkMHvUG9qRZU0/f1R2vtwDesch6hRXeCLPW
aea3AHXB12/EDltMAQxkGxQcX29V+Gw3WSocb+hO7KjXtzJ3uwEj9AvHr5ZA3tbyXFAlZV8u44n8
UT0onkvplavSlumCNYuoxkaPMQAbo9OVWDNUMGmzdnkY3akaZvxVuEm3M7420Y+ZthPk+dBvYIND
EyvSXkAxgBMzbFWUlPpNdZsijnztuQwcQR2cR1C25fj4eoduyPIi3jRRVfFn5fmWs5Ws6/ZPAJbk
+ILg8AqGcbLDiNKcXDp+M5u1c0DdDmud/wsPygyyjfyxrk4hd9PdOIV0aGKl1FdOBTgQFvGVKNIu
Vl+JERnDD6xaliaqUd0A90zjrYzrIsUmLDh1H7iAb13lPKskbh4bXp4pOH4Cjnu6y3pb8M52G6ZW
0ENfU7F8jGQJUyKljgIdqN3y3gLn5GEb9LwBHJkV9d/v1hRIAiWKrKFzyqdUizwKhOo0KV8nu5/G
aSjimbapaCfF2CPD5+v6pd6iocwmKBsJFBqmEQuTqzwmfAj2R8WPKhKmcqAkgdKDntVf28SHZXyj
hz2skAB0YEW9b/XXj7lJPnToShVX/sbKL0P6ug0i+8tWfRY9OZFCd0bCSPiRbdL90IQOvbkTLbE2
ywmTZmqWynGu89Lyao4WbMsc5zwz4Id6r7c6Pssq6nT0fB44Ms8sjFU8j3SHlyRDkiG8T5ZCRYPV
8FMYTE1EFgKQnNg/YKUAvg6IXxQsUN6UOdQ/aByT6w2eXRPwQUcCpvYd47E3lql8EZzWQfDFrDtB
OK/7m84VnZhfikO+yd6P+/uFp6/LOENzx9F7QlSg7gWU6h1V4QXwjy2qlrje9ER/j3+OLdU7ZOMe
5m56838ubao94BcDY8FKtJbb9fvx4F59P8O1ELvm2xZJgg0/OH2q3N8828+aiqrcHA3VwGUObzIT
iNtxRHMhiHSAMsacmQsI2eD2+pom//gM9qU0uupY9xeu9qTv7+gvQS48llVSPJuvbXaH8t4NBrB+
/9t9rwewr7y7rSuBrswSjEIQqg4s8Sy0ClM/QCdPGRstoMEjKL1+BZOrk/DM9gcHvxeTzC0+QoQe
zuQKwnR8r44x+hZ4XNV0E1SwhUnG4yUB3VSABpDx9Euwn/IkxQ9n+AxEY3IL3X4yWha5MKJHaGQd
Gu0RUC65RIMWns6jhz8Ge6yAg2139+diHNtYCXhKm2rb83f+LSD1Krbc6HqT5sCTQ0Wyx/rA5Qug
C5mcSYWIrjkPqQ+V33yQPVYWJayt/jwzvN7ti3+ylP93av8muEYB42U89cttoz69GT5qPMgh+3u7
3AF0EiR2EKvHzMXraOEj6U8S9YFW1dORQ6XiDwu1S1jP9nOq35ySOQlON1jZgjSAR9FCPLLC1cme
JTx4zqKGRZ29HEIpKGLeg2LxVdnRPqe6BFhabUWYM5ZE+ohZhEcJ2pPA8ZzqRpXXQxveXOVYhX2m
oppS9DgUHJEl+gzMDLZtM/b2xx2qXYJ3ApipbFZToQMlHzp84VMPMy8anuq9rTote/dYg2HeMomO
VqO2qgIehn1vQGOpBPhNV2w/PCTYaImwYb9eDVffgbPj3Iesz9hK92h7UnH8BnVkjkj5trqXrkSE
ThoYAOsK7N0caslwqtfn+9TbR18bugd9XcFT1l9pj7LwWGzPTAzeAKe8Ce2/OfW2TiTi4nUgHsSD
pkbsDAmx1RUxIK1Q8Vq7ODuBzOOruTS1lry8/02C95FSDta5wFmIySgxqzofMnf+ScjuDHqWf0Vp
Flr/n30tQVeBazLXdmi0Q4FOMbW2C34jdZhWmhQoO5gwjC+lFauBbf8Dz55aGvrVtibblArf21YM
6hSSpAKsfzpFNCpzXX2MPM2hqhGHs4an8qBTVMf9W5szKd3HxWA3a3NOBFCs7qZbRJzr9p0ZJNqd
gBt1IP/vXwoKUF/K2NJ6qTAk7Pk9GByckZnWD4pST9sx/tRp3kJSNbasvtafzAeiZLzHj9Z3bHXl
D9ZgHYGEjrE3wdWWiAlB0VXJw4GtExyB5mb1o87YelhumnPZsHE+NhzUq4ObrAiKvDvYbi23pmPq
gWqF9qcso9XDJlF3dygyFw47cx0/MCMiOjzKbZZu2xKIQlw6Do8dEF7f042z/z863L/xTI3ZM0dC
/dP+BjI7fNEY3zhlE/kYhtqGweUtDTGoP5qlxX4cfzo45VC0mlnnhKd3WSM6PZEYVMbFEGg0dSrC
mY/6lXV4m3RRYTPc8EaltI4G33danPM7qZnA45/DAMKbDQYEL3BgvYsJ2upWXevEd+KXFyCdPfgT
4U9KBPSPsNF7rd8oBfOcTp1gwCLo4a+RlyrwVvkQjl7EZmhVQzVQaVkCgHZHy6B0Iagtnbngxln0
A6bqZP7fYBy8XfS882/ZvpADVZgxfoctOBVv2IkaemWtGYwPFIvMYsVcL8qd5ldaJmafRYNjnEo4
HoZHwBG08ZpVf+2vcKYCc5VSMiJ5IIWKDIxjSJD55mJDczVBskGomILzJxigi8KGG26iS2TK0oih
e+zdoUvH4quCGmkiIayfhYW9JMNtbQVyBUQTdzu+H07niWxZzhkdXzqjlVUvhM325DNL0hfJyGWg
vldxTGPayx1hT2NSCqkQ2XX2kyWp68KDMYanL8v3AgnoxfNoNiPy2BIgqkVek5ibocfC70DiZDY/
oyjMk0MyHayxoxwuZLxdgzEUipeAyQDCX/gt5jLA/+5EsKG4fQuChKy3bzMFJ/UsoJPZQyU5gsTO
H9f/ISi7nsQNr699cQFoNfYFOxNeUyVD+uJTMB9DmU7SKGeNHWj7jsEB0tr1p2u2EqV40YYeaf3n
rCclIkS7tN4qEll4HKvWfVs4V1dHyETf5SMXQ1sdkmArwqcl9gHu3mNitqdSObJ44Quh6GCgS/Qz
HSKz/XmQMgcAysURyumOw+NRzbYIySl3iPuoNRuUb+bYTra+XVUr3Ho0AYgsMv5iub3zNKi5QrMm
VH8zEQTZSy5x/yOrXTwLo1GfH/miBILK/p21EzuuiKirDV8H8HzRltVNa5iRwQtlpT5p5Hecp1cb
01sAbJgBVftuz7PlDOSWTEmv2oDUm4PuTTLPtiel0D+bKiXegzWVBM3ZhAYS7zaDbe1h5iQUIZdD
FkG0We5Fsy9XVBVtMNEmfzkNKl0c7DVfgxOExWz9Y+2ZffNp4l5iKE/o7s8nuFtxaqyF1V1zEqp3
/OL5bgVnEh09gE6Ra8AVirdgGpXA95yXubNPy0ehksPDBrC8qQ4DpJw85cyWNxySXgbWQtoLSb+s
CTtS2neCcrPtMuwIs7EfMVZoMESZluk2wXKp5gfPqbsMB6l+SPQCe2d1273dKVabGS3WcrC90cLR
pbrbts0yPwcmvIbyL6SVDzvvHNz091Ql51XktIzfOV6SvNb9S6SP4jOIPnHb+6U2tw2rstqPBzHP
NHQNiW+xfC6EKwamGokqDX6t6pLvl74vqGOQ33qRlYMvsQh9E/YqOOsAvtBYiZHjs3X+E3DrzZ2j
z4thkoaixCIrRNh85s5fYRiUTjrYo2sMLD7dWXK+BVy7Aa3ur0oDCs2ZCZw+TWRiPwa7Jrx+uC8F
FW5kPcr0sUTrMM0JhsrTvJmMjvRrYkhMMQ70F2o0xKa/ebjzw7w3ZpuDWIwyt5avux2grLAQILAn
IMOm/JcD3DOrCWy+0z6lBGVLJS/Ks/QQMBQ5Pb5ct5yU6lka1TlIkzB+HxMNrkB9tIvFyKdSFvKv
1N1epGQFXd26WftcFb5s+jITfdKe2qERo0zgqgySZRWT6NgmQUVlwrmen1oG3aFqNfVKDCyjCd3i
o+tBKgmgen9g9qGs0Mj075B1WWHeQWOgS+wqPjx4W3nNvAGOZpcHCEFtNGqFVsHUItPIpfJQDCyk
fxSfGaVpYiUeTNAgeFvXrK6x962nt5Lq52f6dmTLpyeRMXX6m6cj6E9jZbcWikhHnTWIgRSxqmTY
HV/rFt4OikwHdc8EDpf5aGdoZYgyjdsH8k1p9CnvM4yHJwinC+0fnbCcNCifoFzAGbllo5mVTdHk
FXfbp3dbAT5bL5Cx3gJyaD+VEABSTNtDiu9st0V1IQclTQdFtGs1/aKC3lTLrIKumciA2iGHWZNl
dSS7Sx6YzYORfdbDxFOKi3ooMvO6ShwGUAD0nZTtyypZpeIZbASV2P15ryYkrw7mTo7mi55QKZmd
yS8feK4Umazuc6vGxjf/3Fq4oVbZ7EUv2vstRaFzYCQFdEPw6rLJ65B+bUXSXvd7Eio15wPp+imv
V5uqD1+U+C54WVSObCz5aogpeg0aYLlxsjA0C5FhtnsBrdlKtW00kshnKsUvL1g+1p89gfX/pIF1
Jrkam+uUhHeqFWG5ICg+v+/ti8KBbw+GWLqQ8eeQobPkdmj4O8giHXFAmc+oOzKpLS4CzPVnCnt7
SaCfPunUxUoo2cgWEp/xLZqGM7pz9mPBD+LIV3REU6NYFvu8LRHpHhng0hwjbOq5N4EPw9CuqMec
jQNDK2eBACbw31s1umoZf/7xBQNp/7OGEr454fJOimC+fN14EnoGRFyCgwTnBLKtVyB9FLlZNfuP
NxrZm8XkGOVeGf4itWS3W6dLE6mqbAp3rMYeJ0bXB10lWwIcGPgo1PsLYeW286ItF+nZwQO8+nsP
uP87XhmlzcOvVpyhp0SzNGiVAE1l/94RHJcBKb4ogHTOXE0JyvA4d8pCWmTfGk0kgNhJpvyuqeT1
z08x3uHNOmbd1yjLVUYdtoUbOPcwqeIp8rXGNkVdiFNHuvRvxjCmFByA5A2m+j6GjAZuciupXxS+
RCxrR3bYp4u7auzIMHJGMCJwaikLVcsTVXC555AMtjUM8w3PY2riucu8vu1hmo53FAuq9WNhlTX/
nxvZ+AB4M7JnY5RQeBzp8X1bkF7grHINaw/lir4ocV5t0xbb+jjbUjvfo/mR3nXu+hSigLBxzjNv
h/9DGF0+LFmRzfy3BZMjo3G1FLa5LEPIfZEe6AmiqORMtmx5uo+rHXy6O7JejEFiJ5smBt0xufaU
cfH82plzzPXhNLvU/Paw+8myF3ttIPXYIzxJn1OKKFns3hwL8ggsZWT943VKM+pataH9rnJa8nUt
xnt6VjgvF8/EFT2Ji8CwkJkkfWqHr7AHSI8i52MA73HvAnoL2Sk3V5IIJcR+beREkBUqOB+/tBID
I0nmhK/pRbvu26J3qObH1zSvm1NOdl+EtHiMhqGPGjc85z9ftG1sBSfDfK6oAIGco44BsSUKSYVG
NZ2zOkPaR/vHmCEEmOOF+2sQKwBNxWwa9/kwn0dyDeWMQGkgkjAVHIvFI5UoCbHSQqTv1v6nA0nW
d8wFTN0HFR/jfsdvnco2AukChhxHz27buBSQfjjr+MxWgfIBtX6eu3i7DTJ0SIW8lqhrNnDb4SOS
2BO5xaq3Eot5ALCXQ/RIwZKeVdJbcjZhVt+k9hN7Svn62tsO14PgDgsnW0wtrCnarr4Ot4Yt0PTZ
Y9hanRfuKz6jo/yvo9/hgs7bVW4dHZQ1tHcnqE0hlgDgbYleLILfTKQhmE8+XmFNhhy+hBqOShQl
8RSFzQSp8qe2Jf6XAfY47BGCq3pnFFhuDfyH5LhoQx9SUNU+FkrLnP54kpgCRfmoHes5W8tzkzD6
OETaqHeyuXHuzqftpMyQtxEHkXXEM61U9F5C2Iiu+0sIupFzohhUhw0AjxXdnHNsQGMFGMQ6B0pX
lK3tbMsZqr3chcqPgVUrsmSWcQ2tg2PbJ/9zNs9liRCSAdQcy/6XxoM6CKxFGrmX9WYwpl8aOa/f
iK+BwXlUpnh1YtfQXFubf66wY2HjqQJlz8ifx4Uui1pCkJ+qky2ccRFEwBQGxV+uzne4tw4NGK27
WIcoibEnpNpt+yvwPOQopyy4ocpxPXnenjSOdr2IcO/RQbElxNPdsKhF7uS696VtVXBfTv7OPEsq
4SRpeaXpGBRJ2PPtxFMYgCgrAnwaMx9SrMnyr+tw7lQ3Wki1Pre07sVzZEC1vWCx4/xmfJpYraUF
rlYpMHnHr5gxtZfCblE5tpJ04CydX/0ljquDA4s7C26uAVe3q/w9o/v8r+9fc5PUja/QspoKqvaw
Pyl/A8UyVIKYc+Q0aJjLmfo6tai5as6e+CIEJjZ1CtOXCdlz3axKi7RCkzJktpYe1/CJsTVlCgym
f36w0eDhkNOfqAurtlsNoE7fIskYIj7tjGpQ7MsOWCe6wqEBovb7F4LsT0/PV1QqbqN5IQylYbVY
sj174H3gWI2Dl1KcMpm3DQztddiBbV8rkIy/usDWjttElYCDZ51hO/+j+tIOOuHjCOBnAAl3OCkf
NDL+eRKBzhjdKJmize0oJXsqjKAeu+GY0UPpEW1Br6uoILSyCHe8JSgNSIDiVMo4XiSEn+6E0I4U
T1bOJ4BHsfFSy96feCzt/ZzqlVoyu9BokYPRakwWvD1HuQd5YtgFgiHJAeZPMeNb3jCeud1nH31g
PoLbAQx8hVCqqoZWyXV8aiNX1epspeOiPaPyQjff0zxtpwcJRI4bLUpoWK/St8cek5KxfrHCUicP
Fh+FGKdpZgyYIaXWHdyGyXcUFfuKl9vGzLWfNBzDhIUEIGvu5BOdxInHz5OWvGOk+26vd68iFdJv
qtWK6c2o4YSxx6s1QFxO9/O4LA3P7oaAU90VavmJVSBN2GfQv5xaTsy4nzemOEJW1Xqg1HZyeJjR
Y605AliCvNVilVwQQyZMITDNmQTdDXvi6fGnCtOIZ+CZPdlVpO76wdgbgpbLGAP4Yj7oZKAYacCC
tePTw7xq5L8TinXZSIUMNFg9lfyOB/x82ciSSysrzhEGLZ6fpEt7bNVbVaUEgv2jCrau8V5PPxfK
5wqB8cmXdUAnT6YKAVT7rr56RKTVYUVcqgLY44Li0y4+1S4HAQGmNqSGnjM85Nfjxrk95SbzNM19
SqcebMU8Wj6OQzK1Tn5svHAsf0I4zyDL+nuISciGp3YNFzbxZAfcJF7Y9f0rL0a97RGHmzzwhCJX
sukT4YnyJLpu2l62XlTfttlk2JKey7fSayAsptu47vrWMGObto69af6MIvSfjKPM9yOF5iZZQMnv
tOJJXnzAnxQZ2EofCpZBekbbGFVR4+sKpI3GzVFfAEj3YADWypt4j+hXKDqyE729qwgTMpouaYip
OCtqyEniD/23dPixq9B6N/5edorVb3Eu+LIf88ux7+WL+ASUR89LwAH+jLaNVcD1O4e5mYtyUAHJ
VlfcZBuJQXxfNR4VeSZXr9vXhT2Pb2NItMYM58uD8nooNuK4PfVW+QmD2YCIDfigbMrWaNC0IdpU
sA5fKvFuDY1cV0v5BVU+Rm5/LuXkdxkyMw7U9CXyy6drzEytkkg282M6GyY10H7+vY0EHhFDgnud
U9pjiLd/8sJ7bRxS6f7k5PSUu5cX8TjEix19sZF4iFI8Xz2tEQPhQ9r895wv3nobPtZ7GYajDA+E
jOTxWX4zFds7+lsVzaZQi83gHRcOEVi1othB8Dkf78lRCanYGjukHYcmjkL4MJcY0lD+Kyibf45A
jooq6m8ntK7GrdZ1nB8Jt+hftQRJvMspylewVE87c3XPLv3o7KLNJ5l4dVC/cTINkP7t8A+kBTdV
YL2gsniU8CNWjVAh4xmknyFQsxfcSMuRYti88zU94QTE7a4JqM0MSQDqSLz4usSgmTx/eI2uoE3T
Izfs4geJnBtiZaUKS4INBy1ho5RBg2ysui0sd/RSQPFoBjbb2CEGBsuu7hq7DzcmlDhandAkvahY
BXg4YbaB6UutoYF0TvgCsnCF8LmRdD6+NhnUfJnkoDR4yV3BL1HiKRW6oOw9SKkS1Y87viBkumqU
jMDrK8nKvlVqr+gap9amKWsEzun3wlV11ssnbMxqft+1NwxiyQC21A3+qa5D9/G5LZqCrkDw0SP0
MBXjLrM7R8zE9rVWy5xi5KPqDr34lTFFKIqfRsnFSc6AVliEgKeh5XIuFfzWj6E1tyGVPotyTkD3
49OucMwL1qxQjOOJ9NSS0ZbKakNn976oVoqVMhgLzI/Fs9KMyRQhn1l9ynKzXr3DyXeOfcqksYlF
nCfsS4bp1hzakTfETPLcAFARBKLHRlcTZ4DcfelTL5L07sJvlM+qY6TJrUG9iA+SBJ/HCjP/+fLM
U+fyh9m4FsxogIcGURBjh4Vh1esQdwNCOXQbwDvHjskOwY4hZ6+puTaWQhqpefoJrDQpOtqgBvGc
4F6yJDPJHpezx9GhEeOv2Mm76LB5B1mCEqfJiLUFNJ7Ccwrd9/9nmwlSeGViCq5EmdkVCyAZ5wwe
0sICCRSH3EC+s1ru+EZfAvLjXyvFQQZO2I0JUTmzG91GGk30iEENqNIpuqeOVYSghXULqaMkh9lT
SRiinGt3/Jubh6zYJHfff7y/+m3EDgCGbGcsSSgd+1EhVUoroydQas5kgugw5QXAj9HAEo1UlzWP
xFgK/m1heGvSfJVfz+Vmvk8CkmJf50wFLY3s+tU8Ut45igGoqmLROdMvssin8b4og80LD14pmYJg
ofm1t46jsC4s1ftKPJ0nEVkwd6GT69EIhw3Nn8TtPIStQOC1e74ZiCeBQfsO9RiLYWIiKVJkndcz
v0lMWixNaAm/zBXBljOZw8bM3o35hxDkh3IQEV7ltGI4rMLU36Xxn7vuOMhKpxPLo0GNY1SjiSD6
hZMXo4riRJS7Z3xdUdyBVvCE859ziAstrXPJWXWSK822QnCCKENwxjbhpt0F73ga5nEZd7Ude5Ew
z+7IwXrbaFo2hLk/w/unlHnGU8UJ+QxkAZQRFvkT6AgxWJ/CmX/E1ZTN9efpFnLyat7u6nR7CFAk
f0C3qq18IFX8vNR0Ffc2CYx5EMUSj/p2iPFbRSSqkdIu8v0iEN17Z4exVv3Fvoh8bIsMDb0aklNT
AuoOw4PZpopEoKxmZCUcRS7680dQaPicQtqJqwflSMCbukybpJiGpAPkbdp94O85eXXXmGO1u7eX
POpo5kBSfgFv1oLDM6D1756Jg3OpcJYOg+MV2m0hir6voYt+Uvw0BPj15de/cCVP+umcWHlavklF
aRPhgRl5qmZajWp4t3D389DSYsgztNo1yCYY6VF62nq5L6q72Le7RxiNP0KvAskTEGe/33XWCtWe
/uYE+Utt5zAeDOjadY52vsO9aGZmRD1OdQHHm5MaozyKtCf1rC15NJsxjawyfXScMGb7er4ELNlL
bh7beHpyhu+kR05NL8QCfcIZpk/W8u3P9uS5iZsErRDirnPYAddqBm+wKVrwTJDcBvNxkl0QFwMj
83k1LmVNMcCIdhNJD3Mtwe3cTW/Hj9aSFJkm8wEilZhD6/dFjWbg+PLe5H5B2WIJ/BXpuCoKem5S
460BHfq1L7NEgmNAIodHPfDZbVRmTKZFAHcg6MpDl4yYPgeLmXjqjsRdXkFPIpcRJpnpSyiu9K2i
BOWExqXD6H346TriLlbPimkF7hRuhDR33w3cwsqbdpc81R0Z1MGxOMNEbqedaU/jyviTEUWZtQ5W
7CV0Epjgk2Lhejx57u39vukUfFt2+jtZwW4FmBCyMo7c98s8GSXmTHj9Z8lR8tBTOt6Pyn6st6LT
yXl1ezvgjiK8V4SDPEPLgf/e++7WJF1Ntf9vEfnG0qBkW9qzmcRteUpUkCqr06/koORTdCOG5ptC
dEOcfs8zwg9FCnXKz9qpXe8hBhOnUKB7tuC3xGTkMXX0f95Ti0LjFO+9FyU/Ntlvlxc2w47ybL1P
oGKjGZjPIQvkeMTPIyEw82qe+qCAAbJfkNHbOIr0ayupU5gfCpp1v7Zu+LP5b/NkVaEpfh2IO98/
BlO0ST8i0ac+N09cAzCC1QsOcOxJG9Wl6QiMI9DSiD9kWfnL6D3czoUPlx3QbN+aGhpx/QnGmltc
RAinlA7k+x5Zxh4vlEqoMNfVu5Gr2PM2T6hfHcuO76FZvVDFwBKwzho0mOCmYDxEO8v3KbK3oYk9
Zl/+d++3JD461Hg/WpqJFIX6vGp7MaPwYH0ISqNCdZ6mEvWSn1toQ0YCItjXoSvRnGw9uCw5/b4S
0GiaPXhe9TpcQjvMyyWUhwxNgopA5KbyERBL64cS41MEEbcuIssRDckA/7Ky3eM9Ka9YgfhtF08x
cl119KUuKwKQPMgkh36EYeV0S0QWGctj/Ch9MJVeWCdZzszaMGFsAL4lbyePVGDpDqjQEH+zlWlb
jDfI+N2/eiT/4jxSYAJkvfAAGIBIMMnFusQQYiWgBMoMQcZPQh+IJ4DHneLG+06hE563201B5ftx
8YOvjsQE5/g/omi9Hbosy+IAGDFXbPcMxBWego53eCEYMhtbt9XZI5NeXFz/YtZ12gYmtImdAWG+
BwNBPJ0omJh/pUcTpwsJzE9RCBxKoa12HY/1iCNUpIcnoWRcFDmveRYP3m1oO7YSOrQb12dVnGgk
OTuwqNUjus0SVTtuofDPbVTtU++gBDPqCFnlNJKPQEVxRR0U3JR/buHwa7xe5NAkhk8mpu2L5uQD
Fa1H05dUY4IiB9qW7wGq2AG3G+MtNYe7TqtwCA9ClYTgONsmvwVdyXSuytrPp9N5etSfmRjoT8AN
CV3F58ClkUHLS7ztmghX7Ht4S6VbAQBygpsDW/aTnoGdh6u0YlGhQd2pE4B0WWuC37Kxzhk/r+pa
1ZRBZWws/bKVzBpXjrpBUQl2m5KsE5iKnIVN6qAbw1hP4HMGxUWryOUp5lRx6tHg+ldDqHLMl8ri
GtkD/PPw1pnx0iKYml+Mkiaz1mLOXvZvt9/fEKDCIZymWEK9Mb02imjszkpHB3AyGmXtrSi58QYL
YqhgA01xEo/bz71Me/1ZXtfqLbrRrGMz99kqZ3MNBTIIFbizzEIBEkE/SB4dgLQjraUd/LPn1IS6
WdezU2M0oxzOX9RDV1HxhTQ9RyK79EDxXIrIOPwi3LaMdFMDSvlRA+AiPlc3Zf4UiF9mXWl1stxS
q0Sg5zzQku0ijNgJ9xLGw2Zh2CBAAKIszXXfdymrjVIuPtKCNb2tyOVC0zmSKC0yx+QfxgEhTGAZ
equRkBPvgFfom26aSPeEw9SFoLD1M5VF3+916OaEhkje7CRrh7vDDx9wjy1+GUmJyBrruzuzMbTA
24bpriWVe9fiNVxJqYnBBfBqToETOeaP6XkXkXyjNCA08SM65Ujp13J3rxYn58eyDwPxtSZxqIxV
2fz283d43KdoBHhIR/Aac4m//SRLhS2+6BwV0c+IWIC86RLY1O7RuMyR73JXfJnq5JY6VjGFxOGP
TF1EEH+cHSBgdtNOiEd0SxRF/iGcAS7cMFDvy0+0ci2TzJyhndBWrA/vhRnUnQIXBhW5IYkcA4Fk
tCbJOa78zFdJ4CusvwUqx0hNnUhFXvv9tZO9kjqmaniKPIxUkIb++ToBpF76x6SY94ZgpPJjKCJh
lDhs4wBCxkn/nqnuEXmn0i64aKnoAKC59Xlwk2NhDBUPZKBU3JVEqdwz/yujpQMF7M8YxOo9tOXU
8Q4zQHNOC0mUXOKv7fblg8ARucCJ0n3vMeHO5nxxW/ZoqXqvBvKZJzvQwHdAAmtNQ45YYxQR36cL
l62M4kuvFp8t4BxfpUzFXXwf2PJcxfiMw/1gVAUEpVj6HCODZuN6ye2IMpXVx6howbK4bYncDXoI
WNCixCnUSMvkz9GvJbCaRFNTbUc1w4twaSRaUnRP3IU+zNtwtHxrxdfDepp9MczRNJ1Y5tdYKPEc
mWcapBBapPGiAUN6GTzZW/uDzihfCbGUJArwUev5qVQvRUDFi2csbxzcZCn2YkmOGcJh7cqFiJVe
VtaXEd8B4h6+H+TvfkNUDY0j8dLxOcchUYAK7IqNJfcF9KQo4Pdkz2dKeMpR0CVi80NQgvt78Yu7
i+af5AhUzKHxkJm9/b8eeOSNop5nNTlguE7442G+RIEEXCfDYkaeE886IfWPMb8ftR0NZtCnIcFE
2J0NZUP+3YAvgh/KeEbctLRNIlljVfWrgA+ulQepgx+eP4oyrBcF0I4JDa3qvoRtU31YKg9VRWCW
soaekNoZDCojlsboFRpOASnWaZtJn4Tx85xfR3X3JgmRqq+2QcqoyxNSoc4YkpqaVsoCJxJCZ2K+
JcWALfojGc43f+AjpI/L5UqrQSjypdV6uNgk9ouMTz9k+EsYmjmhn+YoxpIOEoHwZwDPm68a5BnN
VBrda/YB1+gxlfTUm3OnS4KsBfRQzAbIsuDd/ej3Pl2W4Z7vdMU3JMNFUXZI57yw5EC9OYf8Ki5h
TOdS7/M3A5y8IV4HV614pklDdBFkvwtBf0Q1r6lkKv0ip1ROE0W+3SKnyXvQfdTxhgWHs5PFQxNL
rfF4P/eR/QwpClQ+8Yo6Suky6MBu/9oGKhO5niR6dJkYgM3+1tNJPjpu/Dg+nXH4yW9yJknIzNpJ
jJ5o0PqXLFD1Rz9LhJsZ5bH1ojxjvZ3CQ6HZAVLNG8lDkPVTT49G1+GF8Dp01Nb+3XrznGH7NrFH
5Nf1YvSEO/O1+U3i3aOV5VR1h9CdYW+ote3fU+ymKpJaoWDGqgOv1qbSOQEs4iI/Ocs3RYAgGUfg
rpiZghW78NEGGyV7lKAaaW8Y4LjgPn1eL3O0PNboQatfeuXDX3eagMHn+RCXU3bh7jLJbAdgidMi
IhU0OtdTA3az1HVleeKlAVRKGZum2vZuSkeDdkx4FiHedjYKe+yo4xZFQCvppa2yc+v2EppxuHg6
RLRMQNDENoEkHv7pHqMjHrxRuI7PWmZtzAvWjIs4JE2NHLe92FKsQsSCgzcvNhVtnSdOe27lPYMk
JFBRV4zYr8z9P5OM29xQmoKTWvNfkz3/8RVS8D8GtgV+Ukw4UeoDdoC9iOAwC86ORJ41r2A2hJaw
ZZdy2AQV+9gIg5c7jNDqpuPk/k0s0SlzCRbWyFXjQmBpVVwiEq113/HfI3NmwlFwGms3c9NLDUDZ
mcQVqosz1lv8Ht7P01N1m7cEDjejpzqU/pm3Ud5bBNp+PrF211raTtjpLYPbFTj9kIQFz4qr1lnR
8WVPpUKhPPu0qkFKlpNluE8OUa2NCjy4v2VCnBywLDS9v1SMAXda/2UAb6MBcYXs0HBbNBut46nF
E09DLvRWaqKv0hy6o4LJq1PCpmnnqJ3fzx2N5BMKLguN7PakBazv1s1TEqgiuEc1/r4UaABpVR2o
rzNvecaWA+44kE3DgPRgiMcdwGZMV0erVN8T+ofXZetwRjD/f6XRS0o+1xgaAtHK3G1k5m0wRFe1
uLV/Vz5q2F75LhzYM/1T7O3lwuEogXCnS1T7CueIqCfC3yhvEgtllqqCdbfVPM0E17mtTmcMiKsx
V+c+E30m4jkBRylu4XBuidJcaoLaaMsCZHybC/k9jjxmeBtqP8KCnmjYQx8EZea8nxCTrGqGOD3e
4C4XHcteg3lqNfpSz0jK1CskaZFClzp54JKx0wMjT7RJiVqt9SRV0XFqPwkvfpjlGDvrgVABRQXG
t3K/ysjWO3iZnRWM8UhH3fY9diSbuYnIISFAfbFAZUROSwn1sk72zLWGhDHofCEsX9ffvUvtuLs2
LmqhDV5zqe5qyYr8MITa+QavZQ4zYIGThuFZc28rBNYhPuTQ1OmhrjjsXO0BTanrKJemO8radVh4
FDegItYA8F+lB5Wa55JMNo5ISJBdkixFqUsNwh4QXw7KZA/FfyC0cRiPqqVuMnb1rseQRiSrkCZz
Hx0lrohAwyeYY4sjdpcKplLeEuxjpUrQZWp44t5kM1y/AIQTRtuOqlZWb8PwmJj6qvuxb+od7uiX
cMcH2hZTIdOAK5mg3ECySrzRWmv4+CZL1kEexl34ZJQBBxsdgW47cdiEaCh1rGkF3vpjf3JBE46K
8WjRGPuGg5xmx4T9uT055fDk9ULtzER5+yeHqd2Z0fnGnDXsvofVglPIfbk1BkKx/riituKsm37O
6CUmwT5As/jBsOvEtdMpt6fdqQRwzNv9fbMSl0kvWgVP6rG4tpF4j1HreHLEqpjPsmMWtlUfxJRV
jO6EgCgX4y+dok9Gp6lJ24S6KLjbY7aF85hS8ugbQWu1TlTVLVCMj3uidhD5d4OJyeLYpXBDu8o0
sWvMfkBBkEafQK32f6OIfaB8iPLCCkYB2puNgSvHE/d3DRQ9Jy0Q2KEbafjQ6xP6VbgQdCoQqVfT
UlPM1pxUyQ0VVG4jLpKC/Ki8ojuia2ld5u+83FEkO5526TAyq4MSba1YDx+d+QI0xZDSC2wTQbLF
J8+Sxb1lOhx/l4Eil4BxGB6aBWHhwdbr08HiMfHoJmypGmnucgpilEvJI+5Rcp/pvkuA97UIlga3
nwuCChsyr1bmzWGbNBbo9AOXgpMUTZ+2Hvzc3dKpx41FHlHBgNezktd7VK/uiCUv8RoQqYULQ3XJ
zq18nF168RzGreQM2xpsqq/0YICfgpHENoQW4//JiMQQSdNab2xA4LLq73sKhw93HFi5fhDBAWjK
1yc1mHRi625jy+aSURo31crDH5tkjLddoiVtqVNFVBNeiFCSE2c50haVdCdiuyFOYhn0NAmA00Zd
ULifmVPkYc4RKCv9mZt41VbzS8AZY4ufAY8+Czy+BIbDlt5oBDwOZeQPf/ZgggX4034vjrgXgqPJ
IWmn/dU03a4Kd0NQcixiftKc78CZNjLxw0MQLAPVzsJ/QBXfoGG6jjMaODexySojNJcPpSvJCqkR
VeLAXXQyuFVQ4j8Xrcg54HnO9aj+X/4RYk6Xx+GgznXtb5EfAXJqhKNNgsEAdM6Yo67P9Ms8XP2Y
Ia18ov9AQnCKcCN4ufPyzCWjJbN1XGIt/Ed796rxfvoJTV8zwwykl9MqxpIoMDFW113R3ydbdMOH
hXUPLZTUbTRuj4M9DoAZyHEn8l1i8xqbTwOQoJW0j5f5OOO2vxxvioYMIYmRE3ZpeTxf4I3bxaeJ
gill8GeEkKYbIDLOvsjc+UG324PTDYyPfhI7nsM0fd+CPIaqtAbLjwfvIJQA7aS+tFSBy0P5FSJb
Rh0pBp/pvhf326PLX86NJ5MnheDNqxPWoskIQbiyfG3sj9H5oYG3Kx0QOn1Taid0OK9fnCl8hAqd
4pReZmq8ukA87TLl4QXuWy7qdJ/Wel/qWFwOUvRD250DPD0K0EDUBaLS7LvDUVa/Qe1okBe/471e
mWzaUvhjBWC7bj9DB/wgF0T0lO5hLlTu831FF/0dn8l494qaz2tDr+YBiQo4+s1ykipo0vpvG94z
8jT5NO5ePfh1h4rXQIFuHqRnb2TV1+TR71+dXfr+Yo++e8B+2r8GPuZk6K4zinMVvHgromALR3tI
KTIdM/4UVV93Wv3ZIiLZDPS8SmnChxpCq2k4Qx/baOTaWHPz1fbQma6OWh4KkkAgkJLjAz7UAtNm
p3XVMKxcNLv9Kbm/e1xE3H3nE+jFAKZJMgHzlfzcjVB17/MEwrPREkFBSLbRrhwMgo6WAhVzvS+q
7hldOAiF5nGWBqnOJn9imL/gKa15/TSrZZUtVOmf4MK2ivXE+3s1ht1Xh268Ttgn8ylSxDWwPrxn
0WaO9vBueZSf71jhry3YDtarQrsrwGywbd9XEdr5Vdg8pr5TKQqRYRdsF2tNoa8Z4RcSdTxTlnvi
OtBfNJg9LK2U/3Cv0FqCyVwkTUYP3zpCZ4kds44LZuE2tUjyv0uZhYClFawE5pT9FD7DzqYwzBUq
WYmR9wV4xKePz+iU/UOGagbQuiaN3zqvlp9+/lq5MuBXCYWY23HZYr9T3iPuBOuMPtmN9/tE0S4S
BjhhYjvnCKU6iRalV6fwtMmoprYoPga9ZPq3HcPCpSstfau/6qugSi0YH5SrnyosEnCGvCrPMIOi
VdeAEdzoe+h3Dna6YKDAzCHLowjawFFjSNT3xneJn/piRFlY1X241VeqHLKZVL4KWcnWyLqmOt8A
bOy5tnqlJ2/fn6HPLN7doisY/lj+lsZewBttlWs7wc8XnG3vsJFvW6Vdn5eo3cplPblITrVTeova
+7Ng1x488lgHiSgOO7oPOPKJ+r1zej3bJb1C/Zfu3/E65HNY22FhXa6JVzE+cMQOssBnM+JgL64T
bwcAkua46Ka0OdhIn3QpYkxC6b43ecIt8tiPUQOrivuhqV+hDhtmoiHiTdKSnh90r+NGmTCK3H4p
OVWWalLuPblrpZdMsPT72pWVmzLU+fEcoZTuF+Tozxrk+7zy3Mt065S5MsWLW85P38pogWr8QOB9
Ss4kwCfJafG21o1aKdEUVW5pB3qJ+nSBOtsIBRD7ujtS6zZ18UMmro+UnYXvUt/fvcavYG96zJ15
6wX6gpY8bCDOEeEBK0+ywKBaOJ051AoNuN0nK1J9SVw8BZkDTAn3yx+a16Xl5IG/B6BGuXapcZ0k
nIojMK8lf8on++HIG/Ocr6eVNk1SIC4yxR/iqurMTYNOOfKzp9ETWzjpq82QSlZw3ozNMWycumj+
ZM+/eJBlPJvkMNKVu4Jys/BBegN62SpW2oPMBl54qhEvcx/1coz/mTWT1yEa4CtVbGlb6qTUNYtv
PM/cpiCUa/veSm0UkQwUTB+kEv3dd/YB06FDGgDibGZTtfInXEc4dTQOB/B5SB09hlT4muv3OdiZ
OkOcMSa8k06G310/TEAn4/BJsMPvOlw7zlumAcG+mD8qldZqAiqtlAXC7HbqIHIFs0hy3m+T0X3j
bsTqpF8UlQL8xmL8+TrOwqhoDN8H8Je4ao1optbp0G3bj9H+RCvVtPJzlvJnSDwg/D556eBPiIxc
tKReTOu8AYJcGHFyf/ZCurr7408QYRvePtZwN01MGdV1vL5hf3r0ftJ7V6UdGg1tycitaX7XrG8a
RPThfUuxBA4SvIWxI+IDXqIzZQt2BbWHDAAGvuP0PKgCTimzlxFwnAPdcFYU/hpFy+DjnsEaTBnb
1GfAK/78PurCNEkIkq7Pk23SdqUzTi9h41pEkn8WTt/hIasnx3NKQUOJwOqcigkLBGKWaLhr3No5
uHSRBcSZbGIghrOg1Ixo4+SKTnKY3yjJMqzRvQ79KmsFkHyOMKdeVqRaDtIVZoajBeuHiGMDyOfS
egyPU2HQLLTVXh71pK0VWlnbxYYJ73AATV7bvjXZsqUmuBYgs5hQzqmCEPqxLN2S4uXeD/2iEDIC
ExIsHL8n2mrSBuo1AtE3lhOMQ/V576DSvESXrzPtF8VUftGD2llqHMAwcRnqkgADprLwUbOr+i1T
uCKkd+MAfITnh3JDKxZ0f3Sh7HwaNVZRxNwGRep8RFvU81BKzZxtAaCEkIurDTWj/3J2ZhXGlusL
UtYRmvQ90vRiZM+SGXG7U8WrQEejCAWa31TgUTwBk5g90tysFoeHfROTDf0e3EPvYohbLBMb0Cdk
4rOkD3Au/5Ju3pFaWUHy9G8Y+gebm8T/pT1I20agxNnjznQLXM6d8RWly40b2TmAp29wgRryLmt8
oMoLOvPozFeDCQJsoeXIkEQnV1JHHKBeFwc+DXOGp9aaiCEMXOOpgX/lwdAJLybYd4qLnzXns8+8
gyycik611pofI8wD8Sshz8rCBjmfXURmoYnL/t03KvYy9soKfubNX+7rTL0LhfzgyHVJ9xLWaV9C
/hB4yB0L9Zf7PSPpu5uOXpmYW93pzYadW7Lsq5UECtJa5zQUQcIx1TYINTGvaDqxe60RPyGyTmtc
7Eq0q1tEFXBOpXw0oSxUFQQ+HNkqZJcZWCbS+kNEvKXca9/gVeCwlcKYkLIEo8E2mQg5qIpg0ldq
VWDo9vShmUpz1I7dxBuVq7JnM5jUt5zF/YNdEPZeY2Aw0iJGnukjDxRoU2ZqswV06Op/IA7Dbtoz
pqiimCUHWN4bozK1dt0wB68PrNso8XDsErusOuAFQ7cPUOxLDNlaNt/c+W6eAHGzeaZssy9v4YDL
Wkqa1EcZ51KJ+O3AOkOyCK4pC6bStkjFCxmwHeV4Vj7wFlNf6wqfV9Tpad7h5k+vGcXb+ydVo6MA
WCDF5H+K8DNX4SV41velV8c5PC4Rabll00kTIw38v4BSTTbkxpN8Cw4UFOHE7GDmdgxbB9uP36hM
bBN19lW9M5Km8qZsLzC5E4R25KJk/0uMM4CEVhmBtV0sh+FzYp2lj8dDjMcY2Zncp0eORDxE323i
sa/aMetnv9h7PQv38F/CIyoSZovuxym5jeQsi42Aak3ndSHc/+jKZPdEa6zbQjitfWgdZIfSgNF4
nJA2I8W64/9eEt7zWDYrxJWF0JKGAxmPZUPbDf69Qc3bszqqnFb119fPFY+7fp/CZZusBvj9pYXn
CItKPssTGWkaefycd0QnwbEVGWOmbh5UNmXWR+C5VML3dk0Trx2Tu1yB+m5E+xDU01sHpq6Q3tjX
TY2q5g1O2xtEnLdLdzcz9Bt9Wwmi4lPZUtqMw7GRVZNAAKspd1CuDf8rRVyCY4VKg7orbjwcrF62
I+usPJL9Bd7/91qo1p0T+6Xft/3Zb09hs338G8Wmq6y5KGA69rywZ/VYnHYLg+vQNBXMEFqmCdIr
QH0qndhmUWdi+TO8X7KpC/XOHaJfvIMTKJom6838dz8CAnyNtWXfT8djY6KTmKeHaQK3bo1u3WC4
nJizhcnOaaHj99Wx+EnBEG77JKbO8+NvSm8impuwbAgXs2TyKh8lYz21ftNBHKy4rPZ8m4GhkNrz
LM5Il1tKJfmDgVllzS+DKOj0xwVFISBUnxahUqpv5uL1hNfW43lvjzG75AUFJ/S2mHbOs6uyyHZs
H4hr8ZxVjzhjCD3O9zb/HGwyZYHVJfzSTjplnjV+Kd46zmEHmqlSX1tAIlBUhqqSMqT6MpkWx1b0
MdtKO10nXDOtE1gXPDmb7d7yJ8Vz8b6HUYHzAZzd18mCjgosK2To0+FeENSaMyMkbxzgClRhJ2MR
RSe/qmUhl2apdU8wmlvkwBmPiJe4zOyclVemfiBw+r+NdZKzNXqqSw+tMq4YQre5nBX0fWeGhj6Y
VabZUcVzQCgmQ1kuMGxeC3wyRkjM1Ou4JM3KPOgkHNbUzX/FyxhPYqSIzCjbwlUd1ZEpXevFzTpx
R/GQfwxCSH7Nz42A8wBMfyXF29NIH2cxbBDgjTe7j09dgeEKlw8LjBHp8S2jQGu3hjPqWXT1a8fQ
EPd4VPJbeiSZTP9hIiDEguyKVkEZnujqWNCx9t9k/ih+RvkWYUxJXE+e3YChO/A5mTJUbXNmV3AP
BZ3MU39MnWC8rxR1ubuEwuTirpIFtn8NamGCcpC9JTrRSprEqoMJXxOKyxPqOl8bp+GoMvZ/2UG6
FKaghB3vc9++Hy+5o0Fs9lfCfR+0oqNhttLDD53rJEM7wlWb0sZQYUktHyb6lWaGJm+YiiCwj2z6
LOwPEK9VzNO/PsE2kwshHQfCx6Y3otg+ce+zx49JenIH3K7fhJ/PyV92V5yIGfbXiETyB9fxGyFQ
aVwiyQMHk3Q3w+66gSGd0jfzA+Qs87HpbCzj7K6djH3BXKvKumIzJJNgJfLXXuMzArN/n0G+rOA0
1ORYDAeqlVDQoeP4ds1dgsA3AxdjI8RcoWDUd58YGeoBF/jOq4m6atD7vOV/datnV+i6SYpaCIOG
56CHjYXL4l5MudHizE7pF3CmiDaYGio6g3hp1lxdHIOG5h/X8xPya1mYyIt56RJys/KYJdLKTKgS
jPwqzOmKMURygmjb6yvdn2JoE6cQ+ygtaTeHBzBb4x8KW60jWpU8ldF3qHhrc/ziYRNHUQhSIptr
5JGmlcrNHrxIQoLiK7VpOcm3mTH0PqNoO05Pq7w9oF+qbGoxzQqW1+YXjm9jFlUQN2NYz4IZ/3JC
4gARbC0mzgDRwPJD2aqQyFSijeEudrh1IYPymnnqsfQL9XcaxDZOBbk0Xgd2NZIIdhNjgkUr/PmP
Y9yPlaRRrFCvFuAZZsMIQ8bxI8ah+E3KCAjX3HLa4xZ6ppULd9xycSzzWOiMDdTh4JUeX5lFF+gn
i35W9XfgOrLip11sapQJk1tkkMHZzZMZknjisuIyWAV5S/yG9j+5tgZug1WZu3gEk+IKZbp4YbLF
NWmunSHFhG+Xlq3ek7jlS1bjsgeg1m6mogTQXj+C+aFomPZLcfsBSEv31zhu2W4ApiVDM1JKahEK
c3n+1xglwSQwwT52UTPDF0dyeXoyZbAQ2h54Ama51YuJvbm5Zz0JMVVc/UQJEkd0/7wqU1hzACA5
1mZkEhDgQyWFWDiryGo9FknRKGF0cmiX9F/jSajqZfrT51OeaqBqYpuZrSwVLPfe6rEuSjK1gVpi
Xfbvo2QXc+4UTNVWp23jeRkzZsVVoPCzU4mIp17uPbuS5IaS75tem1WWZHURLDuWJcSux23++RYc
ufIW88O0m9kWsl/DUqHYFCl5yEmC7M/fL2DGGsjNF4lozWQH0htl3hNSCPd9Mgd8fuFacShjO3EK
6woS+mu8xoqe8vVKyWVQOjogSmnidKzb0UgNJIxZEWwH+KPcLezjxwmQrA0wjv55G9xf3BcW339j
AQSf3qh0mDfAgspHTLwa/3if/CTSQ6eTQBPrG8B2hyyENWdxCO5KBL/HTsjTD5fWlnWSvFO3iJSQ
CoGWYxqZ6v8YCCyfuLMDt/iv00whItlxU2d2ZRHXWIWakCNZ4wGdwioej8XX2yBtekbFpwLmxnOh
lzpB/EIf2Dw5b43vO9WjmbMg6h5EURrGW2pFZe5l+kaBsahgaEKhCILHSAcT3keCULao5A+DYBrp
jqJVx9uRSpXilEAVermUvIA/aFdXkZqVnXdVkAwAtGo5OM0W8Q7TgeZL/BWCG14KI8hXbl4myR0d
RmC8Hz2o6Xv+pI9GX/I7psMQsNH76tZ8/VplZlBk1zxv+ankAJT7HdgFtNSTpGXJCCzt0CqBFbA9
0CHaeqNzCmxD8YjJqSv9nrCXwhn2mTYnXIUa3R2IxMkFMBthGEXG4gztoAMvf/GCH+cXDdv0Mp7t
F6SnLWtocYUNojhw19QpGnjQodFF7dn+3HhO0uzzFEBV3GHs/cFGlcRrjtTaJQcYhngJPH3hy9xm
gFIfAe4JnbrwupkrSpL5aXu2WzJV7bkJrbiR186mhjfnc9bAXpmP79tfpEBhbtZdTh+dy1KlWnZ4
6W/tX6uYPM1I1HHGpsOZWG9MayKwu5t5bXyraAZs3kSNVa9IACxlh2RwiWmLWO3HEAFjH+06LFAy
6ZJZGH+KtwawMCLIuNo9C/Zs/f5AhSfNAYINXrhRiKF4uwW3YVFYJq40ht5bHQ31MORYSaxJGget
unwjRAGfTO5DUyh0V3+gcMrcTwHKkSI41Flka/PtTVJeio/Uc6Ip1PqN7Cl5Qpj6wS8SKWE9/lue
TZ6chHyNUbRPO6u9jsT+qxmJgyfsJQUiohMQcrWpSnYzaq4tnFi7mODYmud4JXW3dFc7X4KI9kge
6VG7OlhBrpaTAAdqGLisq4/0W2yqyf0ubo6PD3MvXhT8gBrho87mP85zK+lb1/yr7h6AgvVmDUV9
NYTXHbxVxnVVdbqzRVMi9Q8nct9MUv6uxtcftKQ11oT8kUI1b9pH8Yth1WCVK4Yg+Lew0TRVwZeE
sGXRR9GjwqNEjPw97r+JBmTfaiKKimDaxqZnYnJO/zPQ0MHEKDbVw+MntbKHhKdHGKBZX+mFs5/m
Vnw7XWyf3FRuq0r4DEs5BjFw3xhKlDiHxsjS5cQo+Lo3xoemwtEKFcVGZZygBPbKr8hStVCtKxCu
WJGtWA5UBNxTWp69QO0Ddl9TTkSoLg/TBOYRCNYSnWg9rld45k5hXjD6QwlbLLux3I2K5e3BddBm
iwszAGsgjc+o8fs9Cwmpyb730ygZgaz2bWM2Xn/lIfUd5ApycDvMjIh6G4Isc25g+gqxT5j+b2ZE
qZSvTR1W0zNnoAbGaw4Jou1Zhrr+3JVtrK7k9pXLZzyeUhnafR39B3zKpqAMMkPhUBG+tY54dvDJ
dQDVsO4N8fWlCDTlr10ZHz8lCyhO3icStkrldvCgKEBsco6XiYvgIA7zVTfCWrKVJ05jjOCMgAvd
FBAD6T3c1tLBncSMObOWepfyfatD2hnpKJgj9o9/+8Cu2YryKUGb0tPLDQmc+IFHihtW6duzcOwT
JG9BO2idvj1LivND0EqSZY40Nw3xmOxqxQ3Wvhx8/bCItBWRsGW4oPbfHhyEmqeYhdw4r2n6M01j
Mwdvsnpp0Jpdz+uwEbPDSNS7H+q0EXdXtFaUHQlph+VH0Z3jpFm/FBjEQ5Yc+2AspBF3O5Xkzv1Z
cDuceupnLSjzAO9+O228wYOVyXhv+oIpsXChWBszLD+Yg91oivDb/73k6PyAKzOTHH82zeI3dPxv
9E+gBC4hUlwP1nUnDpha+WUbzWJElW40yN7d/zi1+Ac6MYhd9duM3abfOhGFOAgXHq1HCrbdr3JB
cNwIYitKwGPo2bPfI1SIaDqvrefVm4sOdxBI6y+MlULjMR69ZDJUFRvoMPPLnOSr58KTsz4q/RRE
xURZuddYB1NvmD41VuwqmSJCvNU/V1Nsx4tSzRmbU9bYfS/Tzz/XIXWcq6TrTO8fnNhOXZqGCLnn
vIixbcVihqEfWL1DPoNDA/Q5KWXjXLvnlm3TC9ozPa5YQPov3/XJfftR7t2TDRv62W+rsQdNwzf4
n3YVcxpBqILwjvYXl97aaNvfdLSC4cRQiNIuMmuS5jVbikLMxJzyXxImMovgQxLhZ5o0DaQrHsgU
8Uc+Goh4O35QXoUvQdqFhe/1kpUYeDWTcrlClEi8IBSjOuZMK2WD3QLo9kwTqQ6sHfnJm98S8dt8
pvs/thGLFnjK6rmBxBmtivScaz/k1aTxgSieaoh5fqa8ktg9jJGJmr2xaRhwd0Qap26AELJR+CIj
PZP6NYrcKZFenD5a4mhhZ5K6SXlpS4PcPRRKH404jgLXPbZfHmf06ZqWTvxHqof+fk4JpJnpmiT1
6jb9NGdADX/k6hbBOIbUW3Wa+5G7jdLC3jD8yMWPlMPVJeq8mCb0XV2QXoYqHYAQbf4UTDtlBz/P
mL8WgPSi9OJItFGhAXlaZlOajeMjyKvLlcoyxYVzYgdq+oWCOCvRBEBYokmkTbWgw79AlKF3MMVo
NGsWMVENuVjNlAB8tw/MCEIcsnGf2vus3u90Baq51XdFhrXo9n+YfP2Hd7eAvKTgFYUArgcAsMUw
3MHQI7u5ppjdjkrvItWC8KQgWyufCkLryP+Bz/414kaMOr34vIj/5kCd/oYnhjPPwo6Zgui8MumB
0m21sWspLed9ouqAfx2TFjbyNuHuw82z9+XnTIuuVOdR8Uewud+deGlieTj388DT7iPGY2dZXQZD
GzhwHx8HCgtoxvbaeTGUz3lw4V2YFhhirvEaRrP9Vsku8WL6poaTR5twfQysE6oXIEVWUbzhLf2H
j0DhxsGNmtC3jqNTdQJ43p9BpCyPNYa8+3AXJkckhURhDBY3quSijaRiDsSGQGYxPctdjoZYXN4T
0akLuwPfjslQJQ7sLGell3yCAkkd7xQWCHt/G5H7vbGO4UApL4LalmosHHG8PzD90Z75Bh4s733s
Qmnfm6Yxbsnju8HZKh50pF3J0wzHRR96S3v9Lay+DGKY8hFWvtwlufmzuBPbBzsDmFvyLpZf1Yey
qgtsQx618p+MeAxXyxEDADrcwWAh4NqtRSVaIkorLqQ7MsjT0S7GOGhzEsXTkImp1G1brEya6Sb1
9ab0+0kv9khH3bXrbf2nqyijqSR5/HHa30Kj6IWi906Rb/hALsAklBuGk4wZAgsGMB1oxHs0U7Qm
dxudrUO7FkYOtmCtvGIV8RLpJj5Neerxwrt9FQ/TU7Fag3cmshZqavPsy/cg5bS0Hiy6eiFq4sGi
BWGf9q+L+7ZyIv45yEDs13hHwttfLc9FOSDJayIZ9FLPNaTAty2rGtg1nUq57oHxBcVeMbuKWgKM
veVktwxRKfBcUW0gM4mnZEoLvg8p6Bn34LyL8/pj1T+B0vee+ci3SfNSfeRs6lraUpBlPF6Hji+U
pryKdf4b1utestRWm07TnTI8ZtvIXM5MM21ZFSf+rsOql2osL4sw/1juYhFsyjoozeOSuY+Y3qWm
N5pb6AWHbtrc20rgdO6MohIPK42kl2SPcdLAy30+21RuJgoLAjAtBln100LLYA5JcZuGdB3YzS1z
Jiteoh6D5zYmC6tJkd2tzkO1qCR0rlXrJUATB1GArRrOmintFoDde7t5SmH5zG4h8aZawyxRb0Q2
HcdDX6t+15BYT4Y6TD052THlqPG1IRLWYMAyRDpBYnh8wonbv+9eUCCI+vmqJjBHy7E4jOV0TEdJ
RwgB/0SYNuQixMURrIY4s4ngjk3cHohQt6HDj+CYYkdAwtg+76P1SgDXLwL8luhRFsw00myCGMDX
3NBmWfcZz/LUhVqoxVSm3COGxq2c0WJtzYzZlVG3etzk45cvVAdjpS4RHef0Kjuqh2scmo+nzv5Z
BeG/knFaGsypLtFT5P/6uU7/K52cnzmb6adTLgmZdhqctwQwPcU0fXgHt5haaesKaRf8XRZf5Q7y
HT5NPz1/5TKE2NdV8D4K/JKR0M96TwUuwvl5sgoFU/mcJykSx0SUbh47UM2kNyF4TeEEZeeKVIej
eovWkmlRUsgp3fWdGccC6aybsKXyngST30lM5uriseAy257O87RpQBxOWZmOiUdrFO7BWtbvsHly
piVJLUzwoFqQwHGU/I4cP8dUMbrUiVABLW5iHRkLraG6tm1vK7k/ih+fnlnWXq4n39UIfzzTfEYL
Mlc+Pkx3q7dpBDsRO5ywXJIUFx4IQz7fyoMzCEuUtklAoQsN38XSpFuD1OUFyaXAbj9KhE84//Qi
K1Ub57fYR99eqPnTi4j9kf9/uGte3x50VCPNMZHloPaK9OYpaH5BxrEymkWHf3RguB/QdRusTCqa
g9jqXag8xV8bAHBaZbbaE4JOHZ2CcXrCY4hewpL/AzQp+Fjwe+q0/Wx9f0qPToIBLbCizj7/TDN7
YaBKNHm3oBplFvUo5ooOUjhPjAAldYh8pnEyyOg2+XRDtwyJRxQzEZuYuiO/ZxfL52mP7GHjf5um
O6jbt0VugG3NlQmy1dxRCQT653NKmisDPwScqHdS9G87u+L9+rhXIlujEw/yT4QmTjMKpW6EYSlx
a2p/jhdAeciVzy4VqQb+Z3Tv7LsL3yu8o8f3JlzgT6Wtp9SDDUOG7RXGA0oViSMOz+VNvEFC2cLV
zaPOiWeIUken/t6CvJFeZ+X8MQ47cmCqWvja8n+HKdSyojHwV4zmFn7oXxArPlI71zOFWFUL/8zD
dvSo3xxYvDbykJFM5CrA8IuN8sH7Fuqr4HBxUEozBl21ryCn7Zft6FK2E9lhG1CsdzTcX62NIN6B
ObXcANt/lkrFwyFjF/F2noZ0ZFp6Py7gQUic4O+zbpwhZEnvLtE7TCnsYk8uuf7OIOTMwjCQJSPT
O8nWD7UZW7qXC50a3AoJIYzPb27N7egSvYWHO+7j/tlDshJ0/VA43X0rrhL94coqj1SpxG3QMU31
F0aJD9S+tlRrpB5z9P4xiGUXfXBDgz/t6KKW5d0+yCeVoJURr/BYebC7NVuNb3oVgHaaFUsguniT
zDW11Q0LJjZFZEXVCXyj1TPlkBLyJRy38xWNyr/Y1HEg/gPrvNplsFI3JSqZ4/h9AoWDjbE+DGvZ
hn6ziHGDn0qn9inejppo340wrXI+BkYDstw7FJcSLqxy/PsZwsyCQWplz8w4yVzDHtmci92X00Zm
WRk0EBLYqLiS38QEjUH1ephGS5rBx7opdPY6DNOkY+9veoqzPMBUubGGP15dO0nWRtFzJzoBiX7n
AIBo12jvou989hVCjxJEm/HoTUyn7RC/RENsTIINvjv/iLFLuZchKp29bmU+qE8gnhtbYWmYYOCO
RZPr/Vq0x6BKCeeJ2dm2m3fQjZX9xvcqDDZ9K8byvQUpp3rtvVwWdBEAEw+hMLjBBBSttY60ChBd
7bBrmcE1FUUNvacRESqQuZzwiF3dL/LOd1l/p4SwkwtMWTFXVT5EldDWuHPcRPJC5Nd/f0V1avfh
ZqwtbEdRSZIZf9z4K6THL0L41vBfwmE3Hn/Ibtk21xd3pUD5fWGmroyEqgCfPTXTIxv9ueyg53HD
oOzrLi1C/cdE2Ts0NRorMAUF55gPMohcAvCSa0BifvqC7f0XzpvMDG0Ms3eB2MaNq8nEvaBKmTEY
1CnJ6UpV8HcLsby3LvfiIa5eyVViVH9jJ/Ol8b7HYB5Ue5Tpn7/VS9sJQSELVpnnGSM1A7FpjEfu
F6KhXD7w1DnxFynKvvFInRSuqti7f8E4hqVut8xvgWuM3plDrQ66ET3g3Ow6jZUUEzwNcMlEYq+d
0+TgRlzFVzTR8YWH1YksFEuksn7UM86ZRlQWpsBAVGf1945E5bZtz0NPcQFjSJaCXvDkLnijFZYO
TUEbJE8amJHwuxueI/Tf3qTsdPVEAt2saITByGhmKxZWy1oO0bHwvNornCBGXDoDUypmhfKNH12m
t2SK3KIkCE4c8ZR25VeUMc3ZexLDQAikLJRBFAGEhRhyQbBvVP5m2SU02aeJGd3CO92tmR4Iuek2
T6ygd8pT4NbLgAJ5eHl7VvQUw6CO3XrTdcl5hjxzUKsErCbTKTtIv3oEDbQ/f6uQ9QGS221w+/NH
8rVpy4S5XIAMnPfConFZ4txd57OkznEeXiDHuaVUX2CfcdhkKUIiXvTaH1CRfxhVBHsrDE17AQXa
l1w995CpxQ/HtwOGSwjKo497HUVsXGMRqwnyL8UC28L/+VE61ewvX84cMYWnkSoi/5OZPwRNHO+w
DC4vOWQaIAj7fBfVcS8c8r7qeW7G9ApRTrbmftgz2lQFKvEIz9F7zCKH+bxyrbULr0o+BDe/OwL5
+ai1xSJDV1I6j+z/wjRuBVloq2dcNQBgG1GSSrRyBKBuP1vtZpyWd7LLQ8a7oa7IKP/sHYQhd1IU
cBNeyiYG/oq5l1gonpbAWmnItkwZ+x0S8hIQ4gyRku5aHWEWnCiRgN3DNmtO/VQs7xQJoxBZxt/5
HLpKM66wwqMJgDD/3qvpHh5PnIiGwwn+xZY2y3I6Z8KW6mvdEtvTXeAJyFCg/gjzE4Z8aoBLylsd
LBfHsvBixhXYCRpB6iXHZxCBybjlb654rXqeKUeHXqQhMKlafwrmNrWdErxYdiH3vByUtFKsa0AW
20rSSv2+/ZowFXOgaVPQRTdjvPNxlonUyJv/IMTmlH3I0eFGqEbEQ9t93w22t1xejTwmwBUIwhhJ
Aj0jhOvJp6rObUdUWLcUcNxQKo4MJrIMT5KhkoB/zMeXQxmYR+NLXzVxDkd+ZemeSwU5KZawUHqj
N/2ue5/tuO1yqMSmrIywO5CUh/z2kw2w0RTIy3XOqngap5pbV3wmpPdBldnPWPl/ui+jcdNGMB9J
phx2Xb0diituPNe6Ms1WUmTW6qRxf2BDCdrnwm6ZVPZG1zzZhIv9F9RQLZHc8moIjbuQTew3L/PX
vl1aXfbRAe29fipoZsAx3p8HP6/8CiRkjUC2bwnYY5OljSaMqpr8Xg0k6udGGCpYFxB9WoWQj0PW
saw0tiWrndYHc2YTjcAyEOJsPmW/XjFYYOu9nCDv8Q4k08zdQN2irW2f0OImAIDHn6ynIzCrEWtd
XI5QwJB9OoZ8X+2+tKeqtbogBwEZNZgeOkynPjtqfts4M4zcp7jWJgbgkhEbEMGrVrWoMq6rpLHA
mJtMd9xrbx/JqYObJR6bfy3A1Y6e1LXNFbQsG6mh1Ki98ZClIV0yfXEZ5VBrjtjfEQgucPMYX14j
anGPKnxgf2wnwB5OggkEk0QyPwfE+wWsSS2lC/UW66yWvQ+1BLrW2qy0mFYRYWIEs6VhwHo38iel
Xik8gNDg0xdIa6zFPgfgsIFOiuOy7jNVA5r8fDp5EDC8yEY2zRtHHzbByNsWiYzNXL7eSmLlTN3v
BTYZpuRJi4FAhwKz3C2Hxnek2f6UXGyS4dfUePz8RpAug0tk665DD7DkhHlNLC9NO/UZGpi1cg9m
yE8J0rlWQ4ZRQRYmNzsojaMWqaLwuzVpVFkQRdO2s9r9+42+nTffVXUNIHw/vixYb4r3sDswK1YK
D0WnoqeLKcLYfEcpReUrKFqIiWCDginydDb9sSWWHp05+AGumT7LllIDbF5/CddVmnOMvd8ncEyh
WqO1fDKwl+ebe3VU5wFYbQScG7J05+LxbsPLBhz7rWUqudTWUS8cporHu+kh9KD8CJsmtMyxy5r9
+Zx8hQA6V5tXZO5Kt3Bo21MB5yUhHriTN4+RrhC3U8NKJPns3GuJMKIVzgzefx5Zm8ZAG7bNDZMV
k/6uFQ/YAkgTAR+8U089wZ/PMqjCkj6OX8B4wSLhQcJ7AsH1CkguzEW0AepERaePA0wB0nfbbgNs
m3xTPwl+donnPq5jHrCbexVRn5wsP8Tb1OMcpduGe+EC/lZAmjOnqOve4Rv2tKNjW5/P8CdJTZzi
RApOgymL5eSSf1wQ4WX2sWyrLSYSIEgefITMfQMKjbW6W0LVDusmjGyCHgLMU/MAYvGRyeM8rvcy
R6OSvdpTxkwx6JKPX/FyYYoG9pgeQLNKRFPwB4IrLQ90ev9Gn8fAr1cU0f1TB6DwYhwiKxXrZVAg
hhifHDG04JapQ5uiCPpvTNixLUu3jj+nnVhdUKOWptJVsITvHYxzu558tOb/X36o99rRlS2Tbi7D
xd3jCpyKm/1o4/7NJ7byBX1uceV1Nc+Onq8K1Geust+EiH3QTmtwGVHxf1ONJgBLcHw0hkS3hJar
gh0ERjsZDflLgGNfLGyn0wck/OGCyUfeGNwjosuFSBwCkQoBHMMkEqW2Y2e+ZPFdGaz23ohhdvP2
9CpvsPXHLBE4t37YQMNeY8L7aYPVUd90lvpovkEVfuvIvZBbXYoRYFS7dqKAJqT+IIxx4ONXnSoF
XYVSsEj9AL45JNyMbrlQZK0J5uoJgbW4IpR2UXGpmQv6JcfA1ukqiuIRrXs1H6bKm1K2+9KHbzbM
A92JWZhtL0lwxMrcZzf7MC8j+Y9OSkwcpVpmUMEQsIygq25tnWIkaiR3ltmsfZ9nQWTOvvluAvtb
FaibxYlsDdu1GoZJtL+LuLqds6wyFrZefMoYqXsAJR+dYxxxc1NzS1ujhm42p+FtiqOoYooYLLU3
cIDbfbKfrf+HYEcz7Kd4Yw+vZ+aTaTFOot8Yhc3wHQWbfAb7ZlhUykrfhH57TMVnnCHqVnpLGAPa
CGKWuWXUzzl2b18tPiAzO11dyL/E971pDTmcBKrjh4/Nlt01T5xkcPyI/iH3lMzDHW98Qj1W9ebZ
tQd3YAVrLyZv86GRtiJtyQLGhemdPr9mrn4Ely7zd3UuMBHNvK8M+nht8SPImbjADJRhAJpMAm0m
qyRIqx3Y+itH7dJdP4Hc7gkV2tzjmfQQD/9qymLrUfgvFiCbrZicE3iOShl65ax2SQhbnW0B/y8l
wvDAn+Qrj00oZTwLniWEm4jnYTXWG6pSPbj35vZNr08bNWGtUYQ8imw6+OX9iAvoOdE+NjyeK0MM
IFjvXoIl2VSRKMKXpqSuQxFspG8Rwg+aVFAjDODL7jnDlqtXxDYfLiCvFZxNytSX90VA6lblxdEf
vKvtVrtfWTWW8z5EnNyQg6pS4t8cysbLJgm72NujFaM52oRQfo3bCdl1kK0kgAy+TOQRo6/jIVEy
kLI1YG/GajnGtYGmiuz2JKX/k3EnMYfrzpuocb1LRVBa+O7AR+vTBLYiPaTXONJpyrEsK3TLJITB
4xNtanIbRvAkX02e7+SxqzD1/+2P1cmPuptIey3ilLSfv0ziB+duicUNdO+ZztrRo0mjIjsXnjki
2sggs9rbpQeN833pC3RgQEcGsmkniQWwIRCXFc8uAiA73TGtubgnIyAKNAvsaYxlalQe6bL0osiG
B0gADmdZZ8rVjTG7DsPUKPe6EkSHByObdfjx98+u1rk6dnVKZAlVt8kCxAtHTcBibc0O2TfR1Mc6
Qcj2rFU3r3GEQcSVn2yC1IRMs7CxETdxKibxaB1OMYXhupmccgMmWb1oUqFt5lwlk9+PU5WNkxvx
sj5zRBLZTjaa7/Yvxbz/2IpstvIpOyJgXlC8L05SWt22LyRiFrJ6vR1hC6ty82/rPup0R1l9eTQh
lfBB+IRF/H1yWHPeI78vbCxFIzozuk6pOkpM/z89SJ/5VbCXzPCD3jbMpLX84PxNkCiMX+T70RdH
plEBh5PhrWwMY7B4zaoz8maNZLLgalcOCWUkv6mYQnLi1NAkr+z2JrzjxtHjZbhDAm3C7l4UPla8
iy4bGc8hFSrfg2DlNXWEzXShnX8sFFXqnmwMcLgo7UyNoNwDHpF0uzXgeCsowVvEW7OW6+vVIFRy
9T+HZGxSWaEUQBcFkBqV/Nm8kg7N1OlMB87VAaOe1K6CqMKmn3pcKrRchtyIONVEVQ4siBqACw0C
fgH8+MIwJWbZK3cCeERNha+RNZLGw4dYJJae0mLMFxFp9Vf81XUr8/OzT2plLuSoioKAERllxPaz
Nz7GofTiHQ9iZ1Q+tL62JQ7q7iQWfLekuqG/2Xnmf48T9ssMon4SHecC+MeFOZR3yEPSNw8qepyN
i+8/v2I51eL1ESZBr+EbEXPuZ7YqGdHxsdcDJ/mpcor3QM4nUwO+1cT3qy9okHA8f3yMgRadZmzt
qyJB8w/RyDaBUgf88+3XrvFDLi+2laUSbUrYo2ofP9fzDS4Xv0ChDxY9kzHZZMYswmtibd4eGCT0
y6TPokGQ5+272ifjI3WPjyomqo6bP6yhrGkX2xXqaBBdr6WnxwaE6+ebFHpCCUMel5V7FupUOaxL
UYF2nRJBXU0+nItApsi9ZeO9zNH9fWi7dgnV9+H3NvMBmXHcl6zoVQM+1dhy9uHI6YrYqJcYf3K0
eJM4WcApoLBNkusfAbS3una0hvk+iaHdnKv9N55TAjQ1K1NULL6WLJWJyDam53Qgaf8CTYHJ5Gsd
9txEYlT5AIgSPnfyocV/7G3DWA3CIi9gG5S7LAJtaaR2041ATpnrcjsSZ7Cm1sC9nHZtUZzpLQ/C
3whoLlYYxCX17mhcEQBGzMFrvGUfi/oD8MVYHq7T68618uyfXJpN8FYlr04Mr4Xw7sObZzg/08/X
tUGez9y8YbwheGzLV0Z/yhxIcijyuRQhWk1SrT5k4XnyKye7GB5+BbgLZkik1UZov7latI30gB8I
NDLKVtwCqNR3rfyU1xHaR++L4P54RvQDzoKLB8sy+1Y62lQCwAytYdQlxer/SIjyKnm2OaifuyQH
LKBMdNcJBvCb2IlHQjfWgFMXKKGzRTDdUmWrJYI9N3iAbLRZx58T4nhrWcCsi3aIddiofPOEbouu
BByGGM5JQpDiqySUTazVaGiYqNf4I5Mt9jp7NAp9A6Zhv6GeQ8J7TKbj6WfHEYpGzukN4Mrjpm7B
J6xh6ioQp98OJd+r1IMdyicAtpfzWiQv18CvW6uo0/lpfIH5x1n7WLILQT7UOQi49vUP8FNkubto
XySTAd3LKFjNPK5b1+X8AvjCNKajYeYTjrWQ4hbJcMBgx07E0wSSSpM3JQDTAMnePlZbx3HhmWG8
6R8lk2z4cuWm4PrNhvwvOBWU4ai0LatlyDki7wWC+ikMBK0KkdIbIXYtrXtpD7fjS1y+/Xl3OsUY
QTbayTPEk9QpTrO2VVfvyWz6wrpPdaOwRlFI6t7poNTiOcTOnf4bZ+2rZTNZT2VFOl4DIb4Qifls
4kFX158gKZEFSrpooBKwY1Pa4tMDsAszkoBriQhdcPmHo4zO8CFSKzyEZguA8rDGXATAsqn0cRkv
z4jBQCxiX8JDDxr7589jo7oho2xBWUjulUtwc2Jwf68KE+MlX9YkWwcEvzD2UJFTYydvxrjx448t
EiQFS+tqfwXi4672ttxnNGZ7ynSXdPheTPTPpgqyYA3EdoZMhNI0lhLOo1y+Y70HcBiG6/8ps2Ix
rRlOqtOwsCsQtDLToCYU0hjO0lZw0ewYLwEuFAemF1yGb18fn2EfR+PSREpyodq81kW5/wFoq2ZB
9thWdrKuyjLS9MrC3ui1h9xlXMREMLklAXtYe2KjJVGTqStYs1Si79Q/dPH/0/Rq5oPfegNN6edz
nfCMT0Q/vR52/hCKN79rq2UsJp1Oymc43iPGnfSJereCjRnqtWTHukHz0rjOEgH2gueNHeo6MYKl
xPY4rD5krGvEJDjV48GVPS4GVLWkrygfFCoRYt0eKuezzYx2o2j6sXC8HMKsupgchT5WXCR1PzKl
+IEbJiMpEkjyUmadIdYivuKkG+IDIOS6dcYJZ7CdQ1lzgE5rVoG5WV7KPkLMkbIkAkax0/ZX+7w2
Z37MB5Oj7sp7NbNH68OF+AhEvUKKsh1oxEVHrwcbJU8PpPwTLRFYs7HN1AZv3OKqb+yDNVjwWCo/
oNzM7OCCBurXuSRFr/vI/ZW/X2MBBg+sJ2+WXOmFQAemst39jwsgqkOGrtO+TxCHJR4q3YCUswae
GErwygZ/Kus22ItgBFE7egdQJmQAMhm+o2/gUwwGSMnBREojvWWbrVT34FCCzPoYAfe9vnO0Ww9V
HF7SYeRbgSV4gl8dMO6vO1kFS9+24mGOg5bMShxH6oPhVigts1bK6nU9nLm+Z3wJbWSWYiykbVsX
ipnr4Z9WxrF/jx46vbLhBDHhcHsEk52XEYqSuLnwoMHz6pUy0OlnFANYTkGF270zmQoQul2v4SGP
byIbxgWQsaUMWcMS41SxbX2EUsk0/11bnK6cortpYjE8XBPD58EyImFeYNZGubmppwaALqLJWGVa
iyIjBeOlCoTKNzM1PyPWunEpjlIUXm4aSK8Fferg3lFxGnulxsA1gXkDj/IiJ0rmVfmeyLU1Xlmw
iUmx8pnrP/74wpATgndX2mD6zNkhkdBOXfr+kK/47DK3lKuUABSExW99qAPlijlafVSN1eM/5008
Ziz0Oug3mcWxgyh/u/46lveEgL0PklDVsN6op0t3Hp/CW5Buyu7Vil9lCvlQ/+iwLE7ml7BlntPU
YJQ5ng7bRVkvfJNj880/XgrRj+YxT7PJfkI8CvFYB7cAYYUPiz63PQ+0oEFDmsnlYvfi7fZJlCEM
FWxVzYvuo4hpRyHZ5LUnA88buIse1IGNHn3gDdon+1OMDxpXct9G6wl/0bFtl0OR1zBGJxWACnmq
tJObEbX7SVC2seunacNzX++orc0xM8ZByWsS+pbWLDxphOYPtV2NYgHtD6MSnnNWWBNAB37n1xl3
rx7vnidq1uXPENEsB2LZjwkEBkooD7lUzAa35tBa5iyhP5BaS6VlnO7IeMSUq4LsnRqLwGtE1wQf
fNNE8B26Jp9JQDBbi3pTmODNwu3zgBPsujNlD4lpURIomBKUtizcs/34EU/iHyRF63dHqcnQoUqM
DpNhn3Xbdub3xaqoSAfztFQoqq1eZN8YJOqq5UhxswZyjHElkzd6X92L6mlRYAzUKfldlryvILOP
MoTay7SYEvX2XQllo6QzWoBkvKExtvKBmLEXCsKRubDyuXw+Ylg6pj/C5TfPxklvxqBvotxN7YAy
pDWqgFJsWsfBd9JWDcZgsSg9gh0j0M1Drre8pWtumc6nHHhVIYPZ9BDLWG39oCm8LosGls+v2JiD
AOjh7paHef1wO2ejzb9doh2tOyKpHU9Lk/wFgVeMIqAbEctnyLQq6xrzjvtkyXiudaD6UPvq/Toj
gkT0IxtsydhFXZspZ9oBKkqWWPu2SEn0nCo1ggYyR+tllPcKqVJZnGjLdSVS252pU10wNkNShUW9
AdU7oMuCqZo3r7NOkH/g35YazzkqC4v5mC8/uRJQWbWYOlzm/z+Yc7HdppOaLFiXRfyDNMSFoFYm
U0yLcAPn85LxGua3q90KkRwG4zUnTPH2VpVfhMT5XypFCBhOVfOn6K1alqpL8GMMhYAx548qgavH
MwRUo1v5vl59mi5U7nv+UScuI7UVFkSDO3gJrXjR2QWpBsUUXkvJgUTd1xr0QJSz3r6zoPxGJ9MB
rH0dfYEyHra+klhudP8fSICo0Z3X2WZzwFMLPRmT0IMMinGwIw3GAkHzU+YKxGDJ9zx/U91DS1Ey
NUrQtwQS5P0lJsXeTaSU//KEsXpZOdqO3jbAhDxXi/BkUSKYoPaxCXvD3nFQXC5/+TDKEtEbCjU6
R7yAhtEaSy/0+eYWvyxXYnUlb2jS8mVtNvwsuY35/0aRSRmsM5jHBS5Lx6UwznTxHfRXW2nlAkFU
MGrWFpb+PXUXNtPof2ZDgmYfcsFRszc89Xl4lc69mfmQaXIUfcLlQmoQmIVwwkE0+lk7a7jStZfw
HCFT0dmw1Naw+3E4aJmVtgWQGA+slatW1dfzgbBOKrU/B+/DA3fA/SQi9th/oZuljIKpUtCrs+Oc
hinZb572eaHR1kvX+OxMlQlnWW5nYioUkXAKKLPKVQ3kBRaGPWfcFOauS6rq6UQMnQt6REU1HaAm
hi4OD1MKeiPuktlZ97zSDgkV2qg0A8MUcNaLSEPl+UWAu7NkiN9eDKFRwASSNcwx9kSe5Q8Bc6S7
W/cBm7T3P800T2rWuIB/rySpiZu3fvXgHWS5eFlXeHvnLBlJfdyTzVyYVQUiTsyJNKAePbA/UU+U
YMnGOT9464PIIKmbVSfEGLFcroL/DA55dpYBm+/BlzHLZZpT3NPIFAwcO9jRyxHfo3VKygaKn1dp
SjLjnCXHjDlWA4yB5GtJRj7Kpgir6Xcs/u08s8qRBs5AG6kXIsnMYnUIB97NyN6QU++XiE5RpREy
YLR4WsVHW5fIcAzCSmBm4p2pah24XhRPv4Z8VqeSSUqs+UPc63pJ3qLxQr/Fw7aWtFVdoq4iRDRk
yxbNCj4cRitvGcNgywhxxkp7ER9o7Pfga4HOVBmmMGN1p1uJEf1wXiMwks8dq9Rvno8fThU/jyIl
E1OfkGZN5ESulTB25aUS74QdZZ2en2UQmTmVE/ZDNiCS7hp9VcUfhGQ6Ym0iXvtZ5DMVsAevb9zz
xFP+JD720ZxS9Ye1kRBwB+ETaInzLZPvbU62X0jJpkT3H9v/h3hSC+f9rXTo7J6Xlezhf+//OCPL
0yySaT5IvfyG2TsLrx862VEwnHJzHOACilYvrTHIjrkGeKPpy2dsHgx4IvYDmp1z9Par/MRW+xWJ
OfOJYBECo5pxWbVMBflI5KxiZnD+U8OR6JuZD56AOHPpM+QeMEc4vpoqwOfBuqynpBreQTjXUSzf
I30W+vR8rNQc1kfv9zEF1Py+ymXZ9FQANf1BE6cqvw7EAuP8VqhB90BMOPftscVfBqvHb+Oox+5F
Uvwu0NRHG+y2J6ru8vu+5ghlIhOE8+Ba4f1BXJFDmV0ihEZlI6WVJLb2nC8pvLyCNMaMBuHO8K3K
M9sZosOrvNGCPE9CCJeHZrG4mtZfX7bh7m72oMg/eh5vCbrlVjyYIYtIyXOsjQ5mcF2rTREucIm/
vkdlIyvt8FB6VOUsMPeHd4/AMahTDu2PHekTUQGjUkh1/LFGN0dOsKAr/3caYg07gvTvKoAB/pIb
bgTrt4d1Pglwqc2LlXfMqmftSIVQwMZJkJvUY6DYew3mWRof7OIL4zAgxRWmW9+elKm6rw1gfcFh
MqjtMlMH8EwoCEHt6fhDwXcW4lG122SVc6Jq0Hm2l4PTF+XDMST4Je4N/kDD7MSBe5YEg2SVDSwN
URML5nMRt6QX9a56ERgydPyPEvZcfC4NNjiYsuOHsqr+jK27EJzdasUnKHJjt+ij0IDxlGOcQS6Z
XF0eDL89LRj2V9MIW8T7DSmAbgHhziAe5HIsSEnsmhGxiEGl878EubslNDzLmt6Uf8KsbnzO4fyr
vLQob0xMOrafZS3aDWpU+IYE292dyuT6gfFZ9RTVZXEYhV/mlrA8kuYphhCbifl4vghJtnfnywN8
O7p5WZwo/0kGKuNde2auQyZD+ftZ+cCdPJd7yqMBI3I2JFcJEBxUMT3gcypf5TMfulcgisSJCwM0
K6rCuG0YEa46rQNALMi5DC5nA/2QAhE2COXt3DMuXKtLe3flWO7IkEiM1dwFmPftZjf3A5LCBc7l
z62rcJKA7Y2+bWKWfFqZoNcdzoWKj0ay/S+Ij3fREutLYzxZ4AcK4PY+UzMDuCXmuAPi5rvASVhG
eHfbN+ArkIlLztLteNLaqIyVhYw/m2fXc5f7K+DjlDf2cFUcXg1Nve4OT94nGs5vmFpDBlxxNFwT
z6o1MOVT56gIJvB8XKXpE68jAnyx5L7Io38tSl7hA0rEePAI/pPe047VO5bNxYwPY0JnMH1pfHTy
WDxkFYWEWzZ7N0jAiX0xplJlf2x+7TjkpizrwWeX5oqHi5FX20QkMBGfafN2DSSoZuTT1e7cG6ni
6ju/6QSf0AS9MAR0g8o/FW659ckb4co7PKAX1dAylLbXPrMw44XuKdmOS6oj2p0VQOi1ugLED9YJ
3DdZhaytxdaaaip7egW3Ox6TqmQ+J4JS0kPxRRwI9+EGmSWL0P+IvCyP9C/mOHGsXqGUh95AxyNi
WtMVFICqLsS5eyU2XBErHniC6+SnEH3447dF5EN9P+mhN5hxAQOrBL4DtSB4TWfu09tKEKzdqzV5
9ORx1U+M4YFWKASNEIBFldfAlVVrpm+jYvOZu3+W4qhB9KGYpoNHWM15hw/R4+Ae/XqBqPezjuQp
kspg75acIC21qSOXWBJURkF+KWPb/mF4tzz2xjmoz4tibqEzAkSvdOvBSXpCpsAgeGF5fJJwwQn1
tFi8I6G2Rb8gBjGaMJIdwGKSltVdxjTvIGMvBi1Z9mzeKI8KrBHX6Ud9YaHvPGHMwPqpxhTGYVsz
TqNHGZUpTQToDel33lf7kk4tznKrhOuXRvAL6BcTxT7o4Jx9AnMqBsYoTlRsF71gloogRUEJcKuj
q8y5y76WVkSEMiGK5K5JTSB1xSTUkrRw7/yW5T2IoMO+FD0feX9flF5Wjdk/Ys3gnXzZDW356cbF
qkPjQn6SmlzXk/Ht8yX4Oa5QA3G8zSUAzGZnRCvBH6NguifggHj14NY2m4JJmtoVMY0Fn/cybtvE
U4P2XzYAJ38/bfx8u1j2mDFdnQHoaLxNgsGr7/IO8JeZcaYB/fh4HFoT7DaFZa43tPIIImNPHvZD
KwvK15a5bChmlcR5rzNXWRAAGmWJnNadqAPtl6/0r7TVHhWIa9amidL3zrGWsbhe1dmuKnw1ThQl
dqK+jWdmLJN+brxqdWOrvRAn0EpVmQHkqeezftrZ8ctxE+KFUHYZqCiJAlkMDaPT4rf1fUlxaPgO
lHnkrhsmt3mmjNrXaDrPkTIMfQhGOsLRDGyC0ElwgsKMGttA4RDtU7iDRsQ7ulM/6U7v0++vWnuV
QD1rdQ29qy3p4+7pEtJUBV6FUi2lwo+kxk2+YiXuNdjYjicqKi+aGMHcy6GysuMRORnFynOFX/0E
N4YB0L49orF5tWPOGM6V2ukDWYbU+L9N7MChWuMOqV9PDbJCNaLA4Ry6zWVxsZZkazMJPyA9Hy2D
/Y4mVpDgklxeHIQOs9HRcfeK7C/Y7F3wJT3U7HBd4IyF2Uqoj357cx72xXLdZ+lwhWnlahgj9HqT
5SknQsRUHkor5pFHkL2PhiwthvYdf+4TL100KUJx0KPVbpb5rP6RqKs9nIEWsWqm9eVnswVHyNSf
VdFFbjAxHGWaB+Jl6cSi2nDLUwuzw6V9hLVine2E9vdDomEja2+JHp2PfCoiXjjdJ/hxZH5ssWGL
VCqDBJ0Ny9jO/Oy3GLra4iOZVhh3fZJHnoM0ysjbrysKFcAAIaRNpOYSlTbdMz/+tSXUeUCsSS2C
lTkYYvnLFiKa/vFf1Ow4G6QdHkvW7EG65ADlmsYk9s7kWSw3waul4KYvpuRhBM8ed0AN/e4Rc6yK
MAGLX5t38CAI5yQ/aGpPLPwAMdt26iD5JlNsyY3Bxb/R5rzBuNg7WaTEkdEbXohi7nNHiBg0GIst
VM6YUKzku/J6dHyc+z1df/3dMdNnYmQjHa+q5A4q5ssad0URElPpSz3ii+E6CFWPVSaPH6jR1iVQ
IU+7jJowZc1efOJmr/yM0TBOEj8zcOqDlrAC9y183cbNEscd7IQWK/4AXsHlIR7uZl9z/XGIBfFD
+2LvL7zoLbkUfXmVYUYyOejYcMSul0aHHiJpSkRKLL28bVY/OcT92Fqkfz7Z2/p1QJ5VeLdoootq
yuGlcSJUVMnLt0lOoCXOTOkCcyWMNi7Vh3UwOVGcCiXX3amFuAM16P4qqSiJxzY/d+B1esMYq/ej
70Vj3b6/qgswaGq41635G6iRO+ODRw3Qgeo3+vGhw48LXg+RFOhFpWFEBLK79O8Bv27+HpnPllMy
q3Zv17iYye1+fIxY+j1Wc9XSkimZMUILv1WaAQ+bgBhpTrKPPp0Am18L844k2dMWf7RtqZm/+usX
L5eUrNnxpmMlV/VOzsENXOl0793kJTvwdiObijJxJyjESoHjTVhBIIT/f+JGfS9skkJCnFmFHZ+O
53JGCBAVVITNz+uxXp+qvXFj/TjMlovyJ18TzbVFh+abkg5ggnoif8suuGbz5alZ/5HIvwxNXoSN
0UMt4BvLV8Qgq79Tf87Lr776UCx0t8jl+eIUI58199qCuLnm/v/4EDtn7LAI4odeafJwDrKNvp+I
CCcG+U6zx+QQ+nv/Xa0PhkR8osu3AOziK9hnwhcBwxjr8v2piDD9vWVq16oiW7hGsJoFrG3A+Xk/
K3GraKtnsOEdJhRneuB1opGO+GfaPUP7gDI6Kye1yzKuPJqmcHBoMLYETArLTZJll7gZ2XbwDiul
BAWdhHDbCyCFhpRHQf1iXSJqzw0egLXoVocvKIOOO0nXw4/Yd874VzqsPWU0MM0ldx4BXJuUNzMT
rOhw43cps78U6fhcVRYSYJ3vIrq+dZZEOFC9ysC75AIj/3bRWPCpE67bz4hLtAdrWNwga9mttGtL
swvbkyfQfsvdSiWBXfWAbgiGHECXHd4k5z28WzzMtfqFc5QzfFyu71wn5XgHabDPmXHf7SxjVeJ6
IQxxzdCvkar/hBlL6K+FNoDiNRD1vPFrGifO+uJomt/VpEW1kK0B6ARvmTIbxs/9pfWm997+ZsGb
Jm5ZOc3/MTOi1CxYsmfzu6/O+0DhDl7ifsLGhGovgkZ96HhK0h+OZ9GueHL0r9p+N+iR+bvaGgM/
r4tdFwcIN5He+FwxgIr43WkNHHgmGcnY1ztcf6NzScwXrkJiskdNiM3CVwQy/6ViPDJS/IF74c+0
NLUrsPrgiF57Aw7G9lM196UFqWdZVkDP2AGg8in5mbhkQRsA1Z06NQAsfN4AD4hPn4Ank7K1rZKz
6vK0vd3oVW9cExKI7TU2J7auoVi+FhyvtOP0XGJtttze+3zpfog9xzzNcfIUQyyIr/fjAQ1l/g6M
2p88MlBfG9bQSlitiMKboD8gIjhmLIXDvooRVwPgOfnkcPEaporeQjE5DmnzjL0pOV/vRyaITGbT
b5v5NDbvacY53u+h1Y1UNugv4SQhQcfH1kSaEA1w9IhG+r1IIBrxdd9ofDvdGPlhsXGU8j9dM5Xp
NWdEnQQaUAgLLrbgWFmpDSjjcSSDULrd4v2GbgI6grW7kjT9GCA/UmM1PX2C1CrWy4ipkf6iCqAD
nsXQeN7LJHSzDJfqm13mdnoewydD9T/z//M8KGbGz7pIbIEEpp7Fd/pnNFE4IE4S4BtjfRlJ3vFl
EyoYb4IBEMJBXgf5HBLXacaPAl4kTlwq5xt2tVMmdipuYCXU1WAcC22vzYFkwgZMfBZTIXy0TPCE
fEgjXqxsBQs4TGBrPCJhehjP+6eU8IxGtZcPdcB1Hca+VZYnJ+Fwi/cSQ1miJMQssI02erU5S+SY
t8CDCBFcggeaZJLAW6w+X9Wp9KBgSttr8mhKCnck1dqv6xMmTLGiANc7LF8cnAb/S/s2ySHmxXvn
ACNHwKZenxl6Fz8BVf6VS9Wfq3eRLmAOt3WReu8iyxER2c/0wp5Q+K4U8xN1xr2XLGfVfJBtG2HE
JdMDwa1gMnYn0eSuX7llGwN0HO0jzWP/HTb5JrwrXsqSgxKJXtF/uzExU/FWwtYwSmtoWeDUkc6J
K5lm2pa3qadrEZXxew9odw09A/vnxoo4mP8EzpgfAxDR2c8fiq7yFk81dmghugU/iEGCiva/ssdJ
ncjY5cmKj9ydEbM7EpFXq71WtxAWjLQaKnEqHWxfQ0BhxLpFi6YR9J1goinNTD/xGMXwDZKAnVte
37fgi1vJGjaJjkr18b2D5jaKYNKJkmkPHFJHWeYmboJGgvbcdrds6CK5el2EUhKbyGtLO7lo0etY
S3g/pjwwLj6Geja1sJ5myUr9cjRigfE3LFtklofnEmICgGBlwdrd9je3PGPCycBx0GtP182eed+4
LUMleign2jmSNbZ3pMOZC9ZhNGpQB7q1F2S9l9oMEn5EbxC+w1gu6qO2HTV+L7UftlHQmWMrz0lx
CtpDtr4xWcXBng0Bvh7/o+qNkAcIXu2nFMyG5RbbFpuvUXtWW7JqokFBMOaoTeeZ4K4ssWUe2yCB
rlK4GEHEX7eiBgDxhMDbKaRbwJE4AEpNQmNMrhlRJoixBhRGoN6VL7Cs4h0WaiM+k8k/7erYRmmZ
GIcCtBOlfkS7tnfgkZaSJG7+49NlvYabcB873+JHcDJDhKQNGOxcvorUVm/ctjtTwMDBcNvyExhT
j/R6PAjkmeMrzNAKPHKxNarK4Tw8kl4XmtNAdakBF4JNk8/lRJAmPxQORfO5h2IkyggQyfSY8z/d
u6bZuUnWNTdXQT3+NzprRz7usM+eZeawukAKXfsiX+3XturaUOD/lL0FUqB6QeHMrIPuHGoJ9so1
7LdOXcZX9NbsTbHTk9Djg0q9OOh6S/yPDHFMeWGeJtU0y2RrSK92aFLHyJkp0/9Yu1oJlERTsKLF
1vBuMRweYc3J0Mg33GWva+e/ofbcB66rzJ+b0AY8HHhnNMFCh6Gxvm+Z5HYLedxd+yAkNqxtsUVc
7+H0/YQ36BzS4Ua6EXRy7QCdLlk3CulTCaZMfKU/HG6oVzeKPRWYQGfs4QY7IiL+fOwDbxUGvuPm
Kw7oCGdQHX3oXphFaCJn02/kS7WzMSbA4njnZwR+VrByqj5OqAyZHvv5EnWAPyxf3qdaOlfR7wPf
nLkggX03LeheG1CjOMnL5CQrKYrLlTiOo53lfWeLKQ46BrGaIdedxgzrMnOLW1J48R2phRzi4mLo
D6Tjv21SerTSSIgmsLsc17JK31qRreCO05Q4kWSNYm/yF2o2Fp4mCNFfW3E7kSo0qWu62Ud8HKeu
Fv8rJDWBCYqyoBY7ZcM68xukji0poRKKoIaxt4nJ2dS+gP1bHhwEpAcCWuaC1PpKXCuAwsV6lEQ5
3qFvSily1kOYn/WraJ3v80Vjf/md4mfTH6aLhE2TuNkeJFrFcqgZtQnJbUaeCyfRWhyvYKTnU0VS
ma8ybxzaUYywhzd0Wg3vh+0CE3c26Fczhrh9oj4GlGXg6hiLdpBhYOiDIM11MKauQU8jmATypzXJ
RG5DfeK9VFXFhEM/1rIIkEjRUHGYq650Etbj4K6cOMAEsqiL7qmCPm+5wIhHeKT7paF/Nh0SZsP8
9B80unh4d2gQOk9iuqpn6mMOPJfISUr0n/+30rCEqUsE7f1I0Dg6aOS/qq+2fA2R7nLKqwgeENR+
wutR3R2NItaIBMfScnj+fgmAjCQPia06jSZP5yEXcVqH8GTxMhyA5u6I7IsOgGNxp53tpghhCmhp
4qoLN2QyWChQHQhsh9a6JfnCtdk7gFGM8A5EEnEOdHEB0vhFFWIQXMBsC+sKhzKoYq4Z54500lm9
i6R7OmENElA1zOkce4WWQTqzl24S2JJ2DCyhOz1Fj1n4kMEBV2EGagciGo2LcZezMXZ5zgKaiaPb
0IQoC4XVEJDwoqavKY3U5fv286xqqnGDlGSqH3JnG9Udxg8aOnkpDzqxvJmsrX6676cZ652uTUmi
zCu0xugAeofUEvY78rst9kMnWfFKgrZtNS3QNFW2XRLWsBP/tCLIJTwcelBfr8baEhYMM0AwjeyB
XeC9LbirjlH/5uyNFYEc+7uFNwb5EbzLdOSeM75HFMqzqQwcNfjjm7/BkZ7yzd237czcSGndpH+f
MP+rIhiiEeDDMMOdtKBFbZp47M12Drzz0TZudWZ9IpeNXiNV5r8bqSYpVjl3aI3hR+Pj87nvuqiR
AxLH/vV/T4fC0iNzP75WveLLs5mYYLqgge6beSUzdWYWoaHVf233lwa0dQnRpvDnSXEWqXp95aOT
gbS6ZBvDE1hPmfObWdZHazKKMcFGUOkEP/5W1l7FxhpsdV71a2tHNkmoOi7FCyFA0v+/rvpmG2FY
CrkowWSDdzXhCt/d7w6FYm0byz74nGRuplCWAKyi6vzskZtHg81cZuT837XjNjhcz5YxQChsdVmW
jpO1lnrW0x6sYJwyTy2tC8WLO7BNCGZQfzQAdkp/nSBi6JLZoR5EDreilZmkFOrmUDdT5zGYdRjU
JFj/8fAfw1S71lihQ1qnPcPwedrNarDBKleAKokUh4SzND062ab+uwkU1T5WOZ/lo/5yYFUi0760
smb7qERunESGcYRGpPpjnlFZYhrH6xqX9aLcODcOparT9iQ3D3XcfFnsZJts0lJAzoLFLpdb4+CQ
gm614QjPXGoqQix/uJTrrwlbW/vCe7pmWY877zEJ+UFX9yqyjFxZq9NvpC2+9bSek/V67yhrdyZk
emQ85e759RDTumudOz1HkiMkMQ5v133q/uFQNoNDTXpnSaSGoR2rOTUkp5HUSQ52wmWSDPd/x0Fc
RNHRbcJldMlnxJbqcKN+CxgxPpB1+9ZZhbg3Uxka0hee1Qrl07IfYb5r4/J8WaBQc6EQyZxtQuvB
UbRCzrzCZcLGjAK6sqKJiNo16z94aAxybk61v+2o0CrvB6kMYmWA0GcTJkosqHM+Ixmf81zBeGr6
JLpTPv6oP3w6AXnt7S/0cRHX7LAMn5S0bu3Ja0Vl4HfEj4YZjvIWtyHMkjndVCkWtwBE96SNMs40
fO4I99xNj4AHu+VKxUTi83di1slRSev1vGWPAefQtJm+/RnwZPZWOUonANaGQMCAJc9mZAnuQ3dt
zo5bzkHEm5pcQAgk5uJYUaqbpmDyfjtU1r+XA8aHVaSMMsDuArhBkVlB6i+Y1gVNOaQeE7EMCLW6
pyQcjy5kuv3VEhZCuBC8C1XSBrk1cg9+O7w6gsdhBA4UvHdbprVNgYXtKA5EAGzTVW5SZml7gnmD
Ml1ugZPhLUuXQdJIl4avXsMRTxE8HODFFM8J2fJ9iJW1ZpYBAdKdLpi/u0NnCqpXPBa57HBeq38g
FBOxNDbzfm3Rk2SxKVLJqpoQ2iygBETgOk6MPM+ybK5BzhAVLcArYvonktvOmWu7iyDQIe1fVbwZ
MfZRnZK0Gt/FVa6rTW8/nK1VY0jpx3aIwMl2MBKURaLkgPj/Y204WjMWBQXiyg3qVYwe3hgpBceG
d0zmsWW6jWITigiwMs8CntX5lTxK6KN9Yx6lQ0tkIcD3/6jDmp1jx44o+dYdyhjjjgmo3sttf4E8
cpJBkVLaYvZ1ND0PagaMYkNSw3YiEVaiWfCLgfKFoV8IWQsYuwVuXzcNjFmr1lLPArljYL1IjcuM
LrI5ylLxL7m9oiLqeQoYGc4VNZhr5imrd7iXyEPDcPgJj0VkrNl4WnxUXUeruhQn9FxSygAWJFi9
JQR9vgcYf2cMxIrrm7f7zqqTQN6PxzYYqrw/GXrQfCbdSGWOfIxPDguqYx6OaYXN1B48bipKLrMK
P8kEOTlvhx6E0JlDmWIRuP6I+4PqvIK7MvDVTGly7XMeIXGw9QFF9Dk2qwFiBucLHoQeelxNZ+a6
dI3oPybC2TsZYUOg78fG7ZRiD1V9Hob/B7pkRnjrteNLuY9/QKi+q3umUnjXTB9uSu8qgpF0ThVh
mvau43Q7N293tlQnoktSGNChJF+6duAgXI0McPfEFvAJmtsu7uay1pFJYoyBDeCzSbn9YZcYwnzP
YV0IIq6O0StjRlffDwc4Oav4KIzyJOfb8q6Pm3g1JiimmEQDnC2S+ArQp/o6D1RKion06QqgMFhK
b+lTrW7a1Jg1c13ULSOtSqjdVJot91Y9oKG+j4eGwGoq5zEvPprpxCRjnmtlQR/7fD2s1Ya42U/b
o6P5vMyjXvttsjtWGmEm7CVIA4aXhYftjiBPFfs25rHH3ANDqPT8zVd9wNWAp39gYnV/fXKE3zZP
wC/n72ayBTvCnc7Y1XFT1LRFub6nt59yiMd5U70CqzRirKw3MQ4G/9p5i1Ffgk8DA4VDcHX404sx
8jqnUmWythne3lzideixRfDBJwEtIM259nWzjl5CIeXwKLm3rfv82grDYjFYwlh+g+8R1o+bQLdO
RyIG/gW/4Ia8XIvF4JkfCztBV2ZQ+E+rSImuudN/syIcH4VAml7g9t4N8iu+EjfXIcVhq9kjUEIJ
/RAixyWBE5OvT2vyOY7+UZZhVKuqeBFCFZBa0i8lKYYMuI5NAakQUvQptI1CzpdB4I2FKri5DKNV
9hetD2uI1HWeHXE+G6fz+QYUDckirWWYV8Q65r4PUBLhhawlZKUF4ZaP2oyj2FUJ2c/1foIr4YvJ
DSjx2QsMbOdfnHeJk/qFW9t5Emr2Glxmb9CfN0wLRrGi1LcLtET/ycCsUerUVSWubJuRjULqOlc8
Z9FQVwC0lqKzUI2u8Nzwu/w8nM8XIErztMn56NRruBObP6v8aUAAuEl167EMaPOr2BTn71qlavha
/fk2iJTITmC+0UScwsIt4wGgPFbW4Vz0CG/eYdZ4WMmFOLCK0B4/5B3TZDob+GwpPyHFPOS7t6FV
Nd/ZZl9IzQZsXtmTCH4JXc/1pO9yq8MAqEDXBtYDKVLkukVQ7w8PqUN/bPgWdWeDGb49HzsWMNLl
HnX3fq7eB+DScnRRftZDFO3Adi0xxCx1iImRe2ygJeSqXIkwWwZfdnzQb202CbTVScQAo7AgF0W6
jYqnjC6+ADsGNSTRe9XKYbnYruJf6H3pjYfcXRdw7tuIYnyrliF+N5aEfhi0ywahEldL/WoD4t7T
nVh2nA77EZqA4k5jUmdqPOgzk6GBrhXUcuZCi0Q9kxfSrF8zS6Cs3PTOSldP1XqW36bCJ7C4b+9s
cDqmAu7/VaHrQSlzRIRtqvaxKoayrXqc0ABEF0l0BzNX/zM2ovbo49kMZnDodydqsH963DeVCsMs
rf5dkbzMiakB/wzSlIAFr33KlMOrtudweGtZvNQvJS8PXmcBrnzi8YqzLaLYuwz7EwTG0WHhlOl4
OsfwXyuBg+v5VUMuSpuasNsPTa8LN7J0yRl76uM0arOPdhH32RwmI0dX8UjNwj/TS50tWonRkEvL
wPoYsQKaFB5rwj2owMMjAR7l0qyQC71xYH9IBcLkoPztw2oaGIIfFcyVC8BAB7qfXXV0yWEiPKne
1991WlxpLaewA83hFBWKB6wu3WhpbMSFYRHG4NNCFip4Zlq4O/BLAIVCk3IErVcU1QBPZn4a/4sg
aCmzY2tjWJ78/QdYx3ley7qS1ta2s9HEtodvdCgzKe453Tgfmp1B/pyeGxNZ5d1ugPDyIhJW5JND
gEwwEmI0KhNuQDFsiuf/mICJ02PfNLv0XG+BKwMy7QJ62sMYrQd1zZVZ9hD2aQTfPTRgTBslIdV2
dPuXx/qL0kdfKD9UWwiBGT/QFUIqHA0+7n6J0SzE1o/IKsZrdy18H5tz09sopgNE2Vp0TovFYhm1
mHqaNdn0OVlw0pSo9yGQR8u71FZCR1bWo1ia8weu6Sj5iVzq6z7Xqn9VevQueeX9Oc/fRe44+jHR
YaJ4pwK1Lj6gCo+k7ofL5hVnx0Rr/WMIeO9mPRvRQay03ITpC32TvgezeeoGIVzos9Zd1S7f0e90
G2ZXPsT2Ah4Tc8MB66OtMXF0XZ2dePa1GYBW9xtiJOW19CIBDSPXn0h+ZdKmHMuKoa4cc08kXd4H
5Gm8ShDH0toYQ2GsBbqgGzX6Gy63KKYMlbz4tDZaTAaDrB4TIOaDILHY5ZE/FLtfNSTXXYpyjq/U
XXGDjLzvI//wVXfGNUdP1bRnfGLsRENkZLgWMpettFjmiohJRKPry5fKWRzrYc5V5dLiah3MAr1U
X17/lhJB8IIjI5yCwGyEFmmGWiOfQRi7VkO3nTMZllzlSI/3zlaWDOXGcvvFvasTj2kwn5FTMxn8
aF5B3m7rboGLp1yKQgS+077PGfiE5CM5tyudyxXJ6MzN/u4TtZH0jYB+PkHNOSUgtiKtZWtgjqdF
qJ1sx1z6bOuOzSPgP6lVsyo3GyNxKKePaPHf7gdGqXLxmwe3HWBvit3evc13wxSYRVsezKz/X8bW
jYxPdiHkbaVFSFH3NsGoDP/gXc2sWGNy/ZeN8S4m1bMgG8bUDENSe3jGcorLdYo4CTRD8i4Eriej
GPhIe3Dld69BtEHEIrAJYAtctTTa86Qe1mXINYEUXx0H8gNcspbmmffVuX/rWce26P7uGCo0iRc5
l/DfHhJVYAxnoYTo1HXZnzfI1Yn+FDb0Fo+1G/9LViMdXgK+DSv/cX93mAMDQO6jrb+4R+lWPzg1
fR4I5/Bwi7e+wsRAgbCgdpJ9nPvO8xxKl7VezNH/vsGCZrI/tOFfDUSnWu06Gl7B8nv7Ml1bNJHm
ptF4OM5/GZ83Q3JzHBV1+SM/5bGQT+/F6OygeD8VKahsXA1N6A12MopPiAc8pKvrgywiM7BV8PoM
1W1FUaKg4VCo+HJ2F0DaZYvctWLtxH9ehIIBuHeKrSFTezjmx8dnnkIaXXHhpo0OqylK3VKTkOUU
W4+7hpP0PDLuslWbn45hUbOYznnvaW4xxXVRejHPEkr64PDTNBvuKBz2VdgJ9s8CxFaivYHirLzY
k3CXgxxyrOlS9yfxhNcl97KPxqBs60DTy72J5116BCyumci3g/qJ6s8WwBNWZGGIibrXBtFxDE8v
WwZqLbrAn+Algru6l0YyF0yQqP46cigKRBsCTaA+9+zfubtkyN9pxn6g6WMvJVhb7dFgYhaGpf2V
6zFbMvCUVAv2j+/5wlt7LnOxD/nl0VMZhebCXJ8x2RWySKBqsewLICGMxwT2mchU01Hl0jjM4JsM
OgouxUPSjEL/jVzQspd4urRpg/5UExH09aT8ZLuBrXqV4CB9MkEnCnWup3xDtFcnPplyNgUAdO5K
bNIgl3P+cgKRKaSbtCM1NH4+Y2BRReGI+K8QDNhPMIp1Z1X9S7uFuULmG9mPHhoJGIeB6hii8Y/2
4jNxyEaLdGONu1QB/Lwk/VI/I1Y4xBtvfQhgg8cdUdf+Hhis5F/AIBNMjyN370OBAqNgNnHCntHH
wLwdhTRpoUFPhoiEAqftzbUo+BqCYIkQKZVtgi9KSlSSakP90P73LcfNlBU+J0kmkt+f5uW7isWT
ljDzOhtKaY/lkqznPh50viZNNewP2+jZBZOx2+RCLApvDZKbQRtKgR839t2XGqI1jk+RlKPZfj0/
bIUGhtORQePyqeKJ8HydJeXfEmvEXtBQQ17x+DnWaTymzc1rzYulvmbjzjaHVsPjl8QqOXMVBx8W
eCpMw+rJvspaVCyv2pqxHNObJ/IlMPYye/yB0j5fT2TNvAhxwXD/962/nsNBJn3X0iEM9SJPbLlR
DGvvgPjKstFVoGPjWnPgAxp6l7EyvEQ1c4XucD4MWJuWS6PZ9CI635PpfQigwaxkE7nWLlEnibme
mFZTuHeeaMAksEwmSTCkVLOKgIP4tqKBjn8cBsWLWYXPJOMYfl0lZS+ow1QCIOZI7Lzg0w0SiSFi
1GUfVAmKFnBy0LA1D3LfwFwwmjOL3D+FUflTl6+wGyxZfNhGJoC8G0h5UImTbWFmZ2V7G9AMYCHG
idFYtARxKW5Ud5lJjKbgKy5D9U3NFYUHwQG/NvUBaDd8Tp8Zi551psJPOlRrUyFhi5iVptgXZbZr
b0oGYmebTkrwY2TC9Rc9yoQIrLJ8jt8XFqY+XcMAx+tKzTBnFdzYGBs1nWvB4LQKm7FVWt0Do/zJ
a5TNk8YCZHxbQJQEcW2aHHBRlrszXJWeDOwD8tffTGNK5b8yKvsCUzMoNnyZNrIt3AF0jPYBZUaz
fhi1bRvSK8Hp6a505jJr2FO+nD9DJ3R1HUS/yV8fHCo3fEzOwkhvTj9OUYSkCrlWnHufQ2JxvrMn
DfQ6d9qksK0G5poaKgoWya2miIVcDF+gf07bG80E7f/ZCk2DZQQuLNVaKeD8VAbFkC1yRLUp8ZIn
o+3xDesBuG5nYIxk1HwoJz1YLPbPdrmalQ4AEhsCQ2iY2GFlMzEEBnNRvmIUTLtrinCJJQTkM6ub
zqAd193JsGwNMFG/torgqFH2tDWqzEjb0jU6MkQonhPwbp13+U6h8uGQU9O7xlrK1I2N6iE47hyd
FhuC4BbTGP9cPc4/knIO9PhJ1zPewwzpna49um/9N2CTiZGTi7FTPVdyL+rRowH+y0b3WUeYpR1t
s2nqCtVWLue5wn8VjhcRAKP2SGVELChPw0XjZRt5N+rzLCFqyCp0bbibjOd23e1+BvZge/f0yRxf
QijycSvZ6BtDWqxYNK16j9XLy8i6CNcBr+sGeMZHHSxu/e02N+YKxEKbZtuxj+joBtWvCARt/Faw
zvrPGpXh6hPqMIQFp2uOf1oyJg9wbyPS0zuLnF3N3J0HEOFDhdBHdBKMVOW9XG8IchnxfV/FZsOF
S3vFTJwEkCcG76w3G5bFjs6wfuYnhrIOgZajXU8QA+PKsIExpraJH1t75+kA7p6mPFy0P7YZe5cC
88/MEYviVQ2vdkpcOuy2HDN6Q4JRTtliUUYU2QECZg7D6bxPZZQ3p6Ym9+eu7TS4Uwl3Wzwzjxxl
SV8HDBb791uwOjF/D2fu5IRycbZGzV8YhB3UxmUAngqjh5i/EtryB1fovvT1gh27Ny78N23XGKA8
id2UwtqYJ66OseCUfa+p7tXIjQ3WSv4AKjhppa9k4WkSAQGLOePyM5SaYn+f7DBQRNt6ooBitS2x
OKg7EacLC/Xho0Iqh3bYVDmVcm9qRziQkevZhHx1/AAUpboKSqFnwTtvX7Yq+/p6fBSJkdw7609z
kBqck+7+lTnZAdiCWEoP7u2F3rJ9AF/CWNL2MxOJgrUDexCq9dV4g68+oRb4/G6ZiV2SbrIMfuk7
dQW5q6QgO90YGul/7LvyYObNfcQnFBRNfBEQXswUIdKP2wRowehGrQIUM50+QyW/GjqKT+l2CSB8
/CAvtApRWL9XfscA8pyJ+1NIApI+GNm4tfX47JNE4qiGa+StFpbhUSQ2gwiBmGyFjdNYNgevfTDV
c0WMY5Ue/QstA39trBTTCDIDi3taXO/+4wEzGrArUbiY8lJjjnCov3nSjNuzc80dMl6JQoZ0FEl8
3iTfFccpsZhUkjzafCVR3UW0BKyMueYjfNWvrVzn0sk2r6URWvawrAE5WXCBc/Wkit8V4gEFiJLg
qJg3pblQvDAnTVO/6ioRNviAfFhemEWHzUlqyBBtcyh03NvNSdCPy1eQRaVrF7mZyrAr9P0bg6Bd
ET9g9osM8qAfhfwOjgtGr4I3k9rdp2CGtLjXgdwV7d0klhmKUVWXQqodxcyVvmCyF6H6o1NPeH0O
9yxMCPuP3TpEduBdRZKQSNU9+Ei9EjVxJxVbDGLpy7JDqmnSKFPTWqJbqcW4i/Kojx27nRWtN3lQ
Nw4b5MEzIKQrAA3mR4V/TiVEvt3jL6HKbLvvls+fgdGB21yU42ttl1hKlV2B/oa357FbYVvAF2Ey
1gE7Bo0ILzVvdAKZheG8UFoYs9g2LJQvrZX0mWBpN8wrGLwDJSforazVuooiemP/E9MFLu5RyDzX
TXip9hbDWrIgjr1ziNk8JR+3dyedUt97bxkL4I1e67tL83ZHtswn3TxdKlHPJtN8Tdxdo+uWc3AH
LQ5GHKNOmTj0PoSysa1WENxjoXfCOGKXLjhvh+dzx6EwXU8sgDW2u22S8C0uRZUfDaOrUiqvP783
XreYO8OxwF90MrFdKghWZCfIvqFtwW0XlJ0f43cBYVUhEQMudaanSOVrz2AAB6l0t6adLQ/vLMTN
QCusfJhEX6oqUQHR2N+PBpCHC5TG7HroW3bwb+tr6rMEE0diMs51KMred2bPPYSyQQEbOUuBLhwo
VtsBYwFzB76ovQ/1YI77QRLhATyyI1eznV5pOV5/P8hqGVpxCOhp5ahzsEVEpJ8QJOMe7jb2zkVI
siQ5ulAvcEFOcqnu8mx0KhM1/kanCOAvpePzFpyQ3FY8Yvo0I8McYrelrTJJ8Xh5EcneI6/9uXK6
zOVF5kAB/FelBHSWz8CAqoZDwfpYHPg5WFK20A7WZjW4KdZGOaM2yP6Ei6zs+mn8KFN69Qu+IRHj
u0JcRKhaCGqt4mIQqE8EWV13GpNnHxTIusTp06l0jIzDssisxXsl5YCp15H5+RlSuOlrN7qEpUCy
Jv+iWYQm0RQ0KIwjTHOu39Jl664TZ8uFYGNjoMsgSJWtpETZOPutDmbgSDY4YYE/zv63eZR1oZwZ
VmzcMaVKR7jsOsUmR2THKh3Z2zCbrMwZZstR+S45JAwHILeCT7Lcs+e1idnJUPDOUeyqJnQvuldV
y3ROIFhueCcSfLcGOp46gfIMK7xLN5/xj9dYTd5pf0P/ndoSP11KuUuapk5dYEhO5sTayOIncfHm
JChu4MJ8QGGqEfJfEqgWXVabVjPgBjP6iV2JoW+YLe3S8n0M0C0YAbSzi7fqfTECddChz+2Bfuxk
AOeK4wE+rFsrpQkqareDxb9WV1/dXHYLEkjORiWuooL54dswlEFkon0iFbZCA0onmtz+gtDfasfI
4zZ29EkMoLhmnbZ9U/MI76lTzM9myXRXWbM5qd4Jc049GZ89YcmR0oq+bU3rlh4QqWxLCsTDC8cm
4+H3KoSb1W8PRkoAcgWCIRIqpcZNkONJJhJ+nUFDDgT1V8seF3685qWXI6MbaxRb0thS5d11y0eC
pPJYrUQG0B9A7mYQOwaPLt3rdclYpfoMjQRCvpZLK8EKig1wg9b6zRdRwLMRcTu7fLDW2tiwNS56
oWyYdBLOUTsFsfs0wWg1TNgWhoa3qY1R0J2J7CSXE6tpzlVpT0Zj6f3OsbCF34y63d/2W52VCEtK
P4SPD8DJmyxr6apLNARPxcJDWr7KkXj7ejwH5/FtYxrwj22rvyT9OKwARdRvIvuect8MH5nKDUmI
bdqrBZn+lsZsqjDH7M2mBunc3p9hcXlNMGU84qxreIso2Fzj0hJvQaYqYMtTGPBrTyf9lZO/6D8r
9uNUaQwhxMjLJWgflBTtSc82AYTu9MiQYO/Yg/af6BoqOiz4fS4X3iUTILoHFe7msFhaC7+12L0M
+mZ8bX0nG9+37u2TiWfq90JZ+gw13CyCNF3qbEeZZZRMFZix2CyIMhk6NXqzc7r79W3Ih8DzUNA1
iGMaevlc5gq/RgSoUsVzJZeK+X/vDT1I1sgL5I0x9dj2/PhoCRteGAcB76ibvnHIR1joSznfr73u
Ng+vjIxEgaMwXy7+VnW1nhpLn3b+BXXUokI3fb8RjLgQIVVvcHkWaZ5frTJT4znOw/nueuyFBYQ2
jYENoWkiLEeOTTvySRBGr5cO8bS8TmfVeeK1Zas7zBcT5iv4DY45RMotv5hDxksqWy1cukPxgf8c
HR/arVuipLty7VWe3KpJ50EyI7kQUWm3Bt4dVNXyb9WTY/NwAAU+qivg+UXqv0Fg2rR9fYCYsk95
z20rAfTZ+plIxSf/KuALdqmgRV5OxDYly3+US4ADnaKVEqJ3hxaahpuuFs6/q0Nv5nXGlgUAqffN
znZLZeH7QEZ6tYlC5YMMH5mVUMv+1P64LKJgVOBUH2mn+Rr2zWnWrdJBflpgq9AB+Hex5KOoyHqr
p5CuozuIOK/ZpfBZdfZTTS5XY3nNhZHISVYSiN4aglzrPHDlYwJCNxBA7mM4hbaiEBwczlPDo4/y
smnjw4CnJDtkiSORsCEVcn8BPyTSwfDF2R/rMqkr2yB+5oEAOF8/B8/aO8oODunPYul3+hypTxQ3
p7v4+JyfghP7EV+vr8d/G0/Z0SvOQ3JmGeEWOoG8s7JkuWxfkHyaN6KtMoLpChCU8km43MEp7cg9
wEgOg96KtrEX2sP5IFrSBTIidLBMY8/gW+N2Zbz2ZXhHmoqjLVlFvol5+OBSuomLMT5Vbd5Vjf0L
N/VbbQUKgC4vltZEfhwiuuz0++Rzp5SHl8KNIDEbHd0RlnV2oXPflc2QduVUrIjAr0qVx3Xiyn7E
1CWXumAOczOeMRYVZuvA6FCzU7DLJiNdKci8SDPFwfSmW9eXTWNUYJ/z+6V3zvtfFatKsNXakuP5
9DIgJXpIrCHd07qwhjSZTr7EO55YtEv5qwyWUOqOaRell1MgsIc+qSbSR/fL1lPPV4SkeBmkpIus
zdJybcaov/bCqPpZV2ptKzdCTsEcKAAVakf5hDEUq6OimhIhSo4kP59GFY7TFibQpD72TJviVGXr
ZISNxexYNNgk+oyvW2G7f8E5TzwBpPY/833kUvFluHCtaIaB4n9wNmDsDZekW+bD6iUwsyuLyzeA
5qW0T2j38i+c7QNAgyY3kmLKWyQUFVWwMTBCLyiwkDtbD+EF9abJgpIvlk6Qkl8RCpczil0IQTYj
isG8X18jIx768TGr2Ah5WxERnteexW84l7HjL8boP8lwUpZ1Q8TwDrw0OmaH/mMjXDZsoXN69eeq
DgoPm4oS2agAbFy/iHfVyGFpYG33thBKJifKdjAyR8QdTuEL1h4Ik4bc89sxsTWzXTJXnAlUiYdj
kGm9cbMT8TSW37l+8krrMLLT+rvjCLDrAtiEoQCQgx/ez/EcovOauLHPjkQWA3IiU/yqSk99TCD7
yj6NP8iuTo3R/QEwI/G9zglP4cHR9+twJSAgZJLBwPQAUCxvI7qvr7/MdUmFlVN3eL85Ketxlyoo
xiJVI8UuU+pqtvxsqtkDnJDUAgITr3s2Kp8p/GPqStLsiIcCQsejkOHPQXO/qOb0CEqUJkCmE8EY
0C24MnkGssvjzIeT9PRxaR7HFeXjJpGiUoObBku+b7T4WhhbbPRRMY5DVDV/R0v18G5k4paQgfm3
wsYkccaJQD9stbq5uFGzJs7WM9AQddQMDF7vNy/HD82OxkRc3wGrXoYiJbiD3CtWPwkvHJpopQkJ
Hc45/JhRIfMUZQbGn4soTsLeap2YQHyVmkwxJW9isDRQYTMf+Zt7SAnrpIaRFtAfnXjsqFkwlilB
gzFhgOqeu83aue7OCuVTsABTBmCxhj8qIe7EM44nvCYt/SEd9vEluHsCFBEM4YJgbRkrdB2DH2J+
ptIokSZ2Ja6m1uc4rUaLSxoQ6f3zzPs9GoafppMggfnM+wtiCX+oIgXIXHsAb/d5F7BG1Te2WVyT
cTLCI8y6CcZEGRAXtw+kYCn3BSzUSCfUWjPeMLls3YUxPb7qetEHH4Lg7BCRqhz7yunAyWZV9Aan
Dmin39R4GG8yUEQPrDKJOJPZwF9CKrJ0ANXqeM3qKvzpx0rSRfAfqlyoHzxJkvCoAtENwa68HbYg
yuuu3o7lbfQB3hhzONsUhDPK0Rsa/QCbSNgfOHXY7Drg1QcSdqI7SKV5FGuHq9275p2kcFxFzWTN
AOaxrmj86JsYZXAnX94YRYYmWVUhzunNDG/G2Hz/p2AanIjzpQxcmlTzucy9wYKvOV0g2g1zTZMh
vEJdu6EWKQ2qOgUN1Th8gFd3FuB6+VZgD/2BjuO26umDGwXjUHWI8vuHOXf4h+k1Z0VRSi3HrLk3
M0pOHGXZoaCapVIfAJzGCT51pZLgKJ4EPvhSau2eA48TmpeW0xdyx6qBVhffriSnB4EUqJwbHfFj
/SW7ufwYryc8lPasBwKnCeq6L5S6MuboVpWv0UyMHU8ZADjnOMREfSYDY5QD7B5arFR2qGf+9Ke6
T++tKkfIvVVV1aUEZTolrXQigdtYPGTyn4gpCBL7CThcjq83d3j4KClpVXPDA3p4gLA4OjvitRI0
3DoTuE4//XxlOxV8I4tcwAXyWT5Rs/9yyT/qZGcoDzLMIOSLay65VR05DowHx6c9hwOa1we2yRdP
mnYuV0zYxikRZRd20TbmtFqb9GCUDI3v5bGbJtd5hlW4d9Qc/6mUMl6YRWW9FzEICPVeDPUGpJGW
Pf/aYO+tjGEaDH3SlNZx1i85R4p+4fXXSeAfYUKem/Bp9WoUOyHw7J+qqnKJws4g60zooQ3JDBTp
nml6fpvwWYpYIOwD7JhWinpc8+qDT9R4v4VR7RbYLIya/wQCZKOzsETL0weBvLZ4I4wLthvS8myU
Acy088ES0F6IcnDCqzeUr+SuKpZtYny1QiS4QrXh0kUoLFXEENtHKB6t5ATCv+m25NOQKGm+H+JY
cp6clXyFWROBP7p4YtKkgYFrVJ6XRMmH6EYLSgu1lvI0gaGuKaa7F9sJ7R5aq5Vtq+TUEz6lZ26a
Xlzm2kPnXHLJ3O+7p/vg1rhXLTECEFPYM/P2e9nv7x3dK95s14qC9SpIVblB2lnhJ/VV3yrAjVLN
DZY/J+CHScTXXepkv6XYWPFSfz2z54mSiRDXFbf8i9PkuajpvduO7+6pi7Vu47Axc7z0Q35ct6d/
tCFyfVK4++Bjel5t0jS4vmWjQfc+Of9Oa0nNGJLH1YFvXgrE7BfJJJPq3IX6FroF3w5cKwj95KPp
N4tLoPRijSDbhugRDis5vRrOlhnsveGRfMTApmWbdrGo31mJFoB8nYVVsk/ifEMW5zEEFmfmMLOx
fMBicNw7hLsAcD14KU5tATWV/DL7NNhwGntxpENH7HxTbEd6rrEY9afgk9G46iBI+7wx/pQzIgqL
4BQRieZpmGzJNxnFr5OYMSs1gE9dgY84lkiVvmZtbbjqT2fiWM1paxN2OQGB4cxD5SnwcOB6Eebz
jdi6kYwTYvK7j0JJ5+Vz01kVIF5eHQNhT1Q8x6DAVM/Cy94FY2wKvU9Zgf4mRms1SlE7t3wpFwa6
7r4F1W6od/gIHSVuLB3lmV37TvGV7lwebzwpAsiNCukJ8rc9QIb3JbPUysVZVtCikxaZduMCXxGB
AHos8e/7LUiOoXpIOaf/QbThggvds0ZZ5B0qRID+J399HcD4daVVPdgdY5h4o0dJNf6BoUZmD7jY
waEQncRrEOzHBtaul/6LWvu9fnblrgVUIA0JFvdmx6mqUg7CDELIy9HNniOhVIsbfNk/8PkvQ1Y8
AsJUEIioBgb9okQv13TRGYtC4G61M7ZKKgUUYLgX4XS4cfBznHx0uMf0qq8UuhP0UacDwfdRhF1u
5v3n5VqdDp+UA252F8IQQE9xR8vpf12Mv2V25RHbREIn0lA2HYaAlQLNg+uudVbRTgaUBOfJVwLM
dRPcWy4VQw+sQdeB/BeNlv5aglCJl8EyY3U4V2G88rLGmUsjPTW9qFIiPy/7xfuOydwcIwfH0Wn9
BjbyUrA1pX9PbF+vq/VmtA/2vfEkpqknUcxX2+tKdhCj7vU2UVV947VuxqCzYqAv8FS+9FAKrg+U
tu9IIWqlbzojEuius+901QuHybioGcwgmciQ+2NGR9EWsEq8K7GdN5KdEjCjAuwXl+2uTCWUsvp+
raEh1wUy9CEy1ANaYBxGiXJji+B1Ybi/cvGFvmxNsvo/iUXn8xL4cBCQgzW+RmFyV5WnQdpGrB3C
+cVlyrt7ai0u9cVfdOfEgPORVcPwClAddCqaTLgkOdX9wXyqLk/tffF/8M/VhrWY5w1TXR5PN71N
rZDpfhh3Dho9cXEg6suNxHuK3mlQ9vtqUyGUlygugI1c35xdGI5VoIHNhYuq/F8nKK7Q79pN2s7x
6HR0uL5S8mnWHE3pKOEUy+VM7QsL2q5QF4mZC5F+a60PLscn91vKdzR1jvBH0o1kP2vD7UDlh95f
dXf83GrPii2gKegzDzaos8e5o3C12sltsVCGF0T/4+Nd6bbqnJ4qrkUN9NU06x+WkvGH7r87b4g2
ykyXM8wYJWsryjXaQS+bgbeh9AD/12i468WFKXQGxX22pOgsK79yA18Jk4SCzxTDfH1MdsMZMspo
INPyqlsRi8NMllsx5dUThQF+vlp3B8aNQ01a+RQC8CcMwh/3ZgG5tiQc44o1VcG+AOL9RuWDmTcL
Q7AgiOCxI6QqIRXNH93qPMRdaKgeXbywcmZ3tA06IGloJq0iFX1csMW+DImo0qDCJ1Yev193/yDs
C4PLRehSIOC1qtwBHIt5o59t39glYXdxeEBoZxwtQKbgRCGFYgpInnUfIN9gxbo5mD0MoVoSTgUV
UwEJjjnCOriTeQas7RmWk3BysHLdCJILT/judOGBchQSFUJv+CP4w8dB4zJq7EjawGwMy4mrBbK/
ZOIaDWvr4LIECax6GPzyFhMTDSZXC29DithzPktmgraj9dweCAMX96hy5F/31OQg8CY2FSqkRF7R
kJGMMiq2EbNU//pwGzs/spdoWjHiax5rPSBy9mwAxx6dk6cafGtaZImG6Mgg+YLXqi9OVtCUsjuL
xLB0/J/9wtLfY+W8sggHiqhtdML0N1FWIumJ1lCmiG8QUiHs59nJoTBRCZXuTmHhV8bOUdbQdSEm
0wc6n4Lpz6KGQNFymuFoB9TLTMI6+6FJFEWUMtUxzb8hxyurChVtq5bKXAzuq2ye9L9ubSnB/Yto
9fpPLFZXqpF5y30lyaYykfOdaSifuInMHy5NOEfCMp3pbk2DbQj0JcRTsd6dXWRuXFRLz7pAntFr
azg3/I1DjsLUqoel8/tmxYGkrs09nRvq6P9yQIPUr3jbvdWS7cafOMCj9Xs+fQfU+awodMam6GkN
Z+QBiUBBuUZFGty7laW0oPCTbTZoDHclnsU9KpxnJl+Moi6heY9iYvdjuomAzPEEoTS1n1CgvQJe
mKUxIjksyv5bXsQjpjGAYLVLsSLH/MKi8v3Jpn02Am2pjyeF0V1mOAeJ71v+W/XCBWYoyuetJzvA
UEQbD+a7mViWkWNa8UhPN9box5zu3yFoytK9ZSWhn2gXXUC+7FSJoOz7UAYDC1Mz9IPyb3MOqY0n
TfYFdRswmdre8K8s7w62uSlKF/CkwoC1A6C8NJF0oCRor5754cr3+5a1EHjM8X5hQyryYO7jN1Ka
wHuF9nY8lD/KLVXqYoqf9GEaYOcHcKZLYYbTNPSUZMCzwhp2BbJ5yz7IERbbTgd1/4DTivRrUQDJ
eQaY9tbsSyTTCtrbxZV7o2JH8JKALwj3YHqYzNpv9ELOFiNLf3utH1U68hcuzIqx9zzij8fqjvr9
GlZdFNgXJ8uLIe11Tm+23JUFwvvjkcEZPPf2cmAKJqIw6HgI5J81MYaqdjTRbPNGG4MzTCP6NaFO
2ka4A+PxMNqmXvIOyquhCYuDjHGXElOzjp7saZfLWuKcXW1Th/f4ipXvjVHvQNcnPqyZNl6m8DGf
Dkg9ILVQuFL1MSblaR2LfabPtZEWKimDgvLQQ+j2Ez/0iyf2JTyLnvawDq+es56SNlTSfDNIWAVM
bXNlI5L4nH9M+mPS87DjyE1ZAIBfta1txVfrD8ehQU5PqFyyn0YtQMGMam3alQRDATF0XPaE3jqt
La0rx1amGSVC8yYuPmrO+g2g9WSp5VITXcbDeJCjPncEb4iI0K1fjK37RzoZIGsPqvMyzb2Eu8nH
wET9sBMccZbcbiL+wO605/+K2ZA4MubP42nVpqfV9djfuA02rh8Np3kNgPWkKL++QKLJlceSsO5d
NclBKbtO1/faGK1PEAr1FA/xJ6as6dlbn2qxHEzHHe25/+XA44koe9gFubT3R3650xkrJFBcoAll
1Kg1qlKDyPDAeionfD8W+81XDlgeR4fpZdZyvCKOXPfmRxRAWcBNq5hzTXscnFT2APzoyYOl1C+d
6PL+w42ij21DWlMWrGoj8S/B+uPn4K38Fmj026flgmDnCgRMkBuNDVvDTogb2zAasUCIFgL0Hi8U
SI/h94YorxKaigThiALxjw97YxT/uWcjCYUXFWpTh8pBdMnwchQvq1WuscPx1GHFSadcKNwvhaxG
GsVeHo0p+0NUNMGkNovHZxxKhzy6x9qWlKXMuMPOX7kBnYHot8yGWrd20FvlO31ZKxyff+hoxdrx
yWSZWJ2B14WYcRrznUc15eiuewSnah2rtATPsuYh/kwSqLfgCgyHCTZ4boOyLh5umCHAFP0cXRPv
8jTgLNoOOL+JMbekgRHyl7xv/nnnACymHapeesXUBpB6ngI0Eon5MNrIHi6F/5OoMgbLivha5jJC
ra2ApDhVn/i9An0E+C26PW5MwTz1ahtKA8ANvhoMkhisIFsrxGGIh+j6OVJ7BOSN17KCcI8Pn5wm
rwIZ9CwGTn/79cUeiFFYZyHfmFYNLS2t1pX/WbYeVZM5Do/bhcjVOSP0zv+kyvuBPxEZ4AQmyaUj
kMH3aLYOwruWjmB1cjYIxWEisMQ5T9DLWLijWGzx9Ahg+8JnBLSjrRER5JFDWPapYDSy7mX0KqkN
rVd0K6x1/Mf9B0DlvbX1ON5deIpB0A3eanbTgQm2Qp77o0JMt/+CtKL4Yj0aXcD9Cdln6UGaCIkD
IKaK4Vz8hVwoKJ5R4ni6AD/wKeXqlSYk3cFZXMfntAu8a93myz22Rn2U1GcmlPw1YMVigWreKoIn
qN0gBukQrbUNA2qMK4lKnmqMUM1vDrbsRmNmZsASAv/yPNQFj12OmskktPqtklN81qzzv3EmH4XT
hN5P9BjFKRjJsD2inRxTduzdwv9JLb864eYL5Ya8xm+a2KgQeidtrCCFml5FoEUE7paokh7ESn+c
eR9OD64rCT2hEilcb8I6RrcOIS7OwCAPFr4FDQnzleoDmDmqvxoRXMIJnhnciARVS3Ab0cwY9fsA
A+bl2VOt8VI2ucqxgcMF8Atu8NhMxEH4v+hp2LfjPM4Hkidb2inQlNgzKxp0alOhrOD8W8NN8mfp
mLxQyCLLywHHt/SDrlD1VlKnL/B1ufM1Cr0TTq4gX73nwod8HwqzbqQChxqUd7VES6xdEh6LkT8E
tQvrWcHs0hlB+0r7ZjJuG/jDnX7Mlyilqav0ZYJLEN68fm/vOWK4Sf8WLS1Xw+dEpnmRLPxhS05S
QR4abRG4B/mmG4fVqIwWOVvgQDhDwuGHafxNJMq5sQwWRiWJ/aftilgevD7OgxmluYjssFOKNHXQ
1bF+fOW0RiUmcXyvFaz+jeVpFSFHuMVQX4iB+D9oXNm6/CfOSH5pmB7qv5wnk8UtxP6TN2V8tJp+
CXTH7+q2e5dAfIca1zpD22Irelrj8v58EHqHOM1GEQPon/wnI4JS98b1JrX2ttpWVhmIdGZj/Cxd
oDE3TPsm8GWZcff9FaD0MWvtlaRfjoAPYcesxCqR8ocgNMkrM8g0+Gu7eLOIlCacUbzk4rp5kYZO
ypxmlbBj4i0qThePHbfslAb+YLIB+mGg2kU1WyO8JMI0A3VQRDy0yBCeXoZiWDqcu+B6eWC3xPF9
B2oLuklv858xWc2LNtSP00y7/rCz47puLXmhPAQj29WNpEsUuKMgwgh/+DNVhLLmipgDpqoP+z5c
q1JjYI7CjEhyqyd0H0WhWbT5gTzDiHnG5DR1fO1RLdPmf55Fssgu/ni1a7aQmBk65q1HDDuAX11w
omvqRXPqA4FIwzM4HbfuOBtBdrm9FUbDxg/TIqZlFUjs3xRxKASEmHUPAdXLX4FV4ppZI1DQrMjv
GXLX4PLJ76Xv7byrWLm1K0PBc7yO/vJEcvFnSdvWtyU6lN5pX1FWqaIjtNH9VDdscFGKlh2jtHVI
eZr534hsaG5Gb177bcLxPTIQ2o8vmZHU9oLbWG7tEjbbzu++ln5O0L9mSS6Wg+Ty/l0iU4Zkzqer
YehRyQppdQ9WxdgiOVUcMZz2o0zLfTVvabylkapVnQ9bG8th8mxaxmHvOeJnnz1wT7RsiA93bxtd
cJuMnEJsFKi55xjmrs8o6RI0dqnGv/ZQFLR0rGvm7wtMMF+cIro0KCiN5NQJzAnKwhNXnyszhsnC
XfgNnbB1QXm1vcB11q6yhgA+mxPEtLhRANpEjabYOSW5hN2gpZ3bPxv9vTXtuffCoOTZqb99Sely
vaw2fh/bXrl/Qrh2qb5Skr34coeIrD25kjD/DhAfEnDBM3OAoDWBSOjvnw84keri5vDs8uRmnujn
Rsxp5ethu1l5MToERtPQA4ph8PZ68WXq9CUC9fRoN/RFaMh6JoUIRumN5892eAZUI9PPdQKv+cbr
RkZWEuN4bRviisnzwfUEeNnbrHx1C/JGI5wlrWtNJox2INtL3YfbMKVkDVw+6zJ5/szrrDVxCp58
sWFa05m1PRGzQAWKFJ0xnxO/jLk7Eu/hIZGomcZ8oS8rYaV6vR5mherRQA6JjzAUXL+RR/+QPTAE
7fkCIv4n303RCqB1oYWLZYDnrARj8XRO1FXKU41blvLy4nqcNWbVLicyNi8TPDETWUmmBu8gkUmd
eZAKGkH1jln7jmZosioaK7rRnWx4JSEP3rmhtcpRdVHUOBaPcsegEOMgVxoxpDqNsnZm/YRqz08J
cTmgbpYkSYyOfrJUlRjiIN2OrLnKwABQ27LZURfZ/JmEdyoXg/KFRyaOvpJXv1mu/XPX3Yvfi5Kx
LCu4aSQaDeEMThEH7p0dx9CAhMwqBMykUFPb3zEzI0xIrdZ2TDW2m3YtPZHPHpNieIj0Y0PNuu9/
VsCfyDJhe6xDrf8IGQTFg++G7WwpU+uO96UYdJgLa3bjeADC+VVsLuf2dryLb1H9bfbyq3aPaacl
8oiqfhUK+O4zGxXQLtVjzjDWRYxvymncsPDpAp+kHkKUapEAv3qEf5j2MUxYljMs1er3m4wRGGXb
Cf3J6eaYYWSwZpUlWi4F+kFnuDRupjvS3FS1RPqCLW1PLcNltRr4Awzhj6gaLVN2htkd9H/xnlGG
15q4Tw7ppJ733IgTBXoePvRm+nh3WUypLAoumFlRrzRK/rjABjYWzySY06BoyH4cWJewc09HGWAJ
JqjQOeRrR2/sZz4QEhZVeZ+dYL19D8Of2t1Sov5OGg0+9E4yCBU5hTYEecx10F5JnROkXouzAY2D
mjBRMqESgsrJfdfxibnmxNktyGB/7oGB/HLFCJm2WWpCs7i9PPu+0x9Pcl+V9C4a62H2n1JWkLqB
SarmvuIfjgU0YpitzAqUVGUmYxD/Q9j1qasNFhEGGW+6A9UFNmM7W0qBf0vGCFQigFoHPtMtMMjd
Pa6C9PyZ9ZOsreishGD65bo7hRtIH110vmrS70Gbu/hPbWu7QH3Wa4IbrP8DE2ykDKnjmWFhO6pS
BSKU+Gio3GVzeBmiAh04eyWlkGplBL3SO8UX6Z+k5160RMkZ8muGIyhJz7HqfEGc8HiEXAy9omqb
GY6NSyUEaXxjWnsylW5dHP1pfiwXgIREL2fQukwj70r66qXyDPcZBaLd5MSFplv3Gu9OQs0MHtQV
HSqognXs7KhhUdSzcdi+bG1pBdTcyjO32U8qzewoMe4xcQTi8YPVwBRkCTMsIcmlTJuJomVR6Cv5
fRBxyrCw5iPwBAZ9T6QQyv7ijMnIABZAzcezIdE+naENtv6zDDij9a0rPnKovZHwJ45bwTX3DqCQ
+i6YIx/tgep0oq1hCcW7BXVX2yNFkuY//P9kHNnVp+PsGJO7y/8HClA9eAYU4GmOeMxwmkaIV2oJ
bzbxQjJXGivLVmDtRuWZA2o51iP6SQHqVKWPniP2B/T9ucKnlubvjyGxKwoUx3AoT36hnFE/nuTJ
Nhd0LBWza6VDFWadky5GMaYeaRiYc0/RlSCJ5hw67eHOMwuakdgkdYPShOjYB3BkXwX0/7k6QsC3
Sp1UHXMvlnGPlRUDzua+Va8uU9ALBestNH/46SWsSDfmEPqIV/+Vv+hv1gu9nDBKe6itsyGUGHz0
uX1dP9sSs+ZF26WlavCO7RGtHhoRzpHwHJlDVmQVqPsdxlCJt06CQVwkNrHMxLwgnLBKRybRrQbn
6gT+G6hGEhox75N5QqRiXfYEebbZvOmp8TGY46OLSspEsc5AUx9ATkFTNYrC8tf7f2fYyNqz793k
jHxqwYf16Ia/we9bYLYcbWugRd/Q7Yp1gc3iD5I83clxjCHrQcvZ9TTBbQWGbWJnNRG57TFL2K5o
h17DteASgvoPAtxBSuR8w8TopZ5VIVwVPthrQaaS1hNP6Sf9bTAzrN/97DyO+hn3MgazgQLCJr/r
38qH0CSBTAqEoDUuYH6lVe1YgttTYkHjKAVw79emwYUJARwvAq0IuhtFSz+cC4KPg4UdmYw5plfE
DPM2BO5eFA5Ir+jS9FVkqZgmDp8zqrVB7PoIbm4UwcFkE4a7YKljCAjuR1eVLYL+Cntya2htbVHc
UeD8v7r6/rFmHuCabNk/mdQ6BfkCI3EjG631+r5JZNkYX1UH/LH9NQ1piLiUMYqY5X1bIKt8WQqB
NdGHjfiXiwoIEoVrPZ6HGkA9EEflTHqLqURGu34MwONlf2+R2tmAel0Lg6wd1RjZjzlA6KVxXDCC
zvxEi165fmQ4h774BpBQKtMl/OxetbNWQpL2kDX8ACvV0IA5MucAb/WI7Upg0EzGv3qJWEe9xafD
9Y3UjrBX1MXbWlB+bGwIeUM5ESoAXB0QOv3B85Li5NiDz8q1aRCwIUl42sM8TYsLJP/zibcA0Zll
MCc3OCahjJaOgFYcBAEZNGyG7L1WU4IvF7gFonmdXCU8YC87lFm1omIRhkazRF3sqZ5DkOMZgLLA
0nVXvyKMNh1rc9uXioHZfVpusm9IVje1ddo2C4iNdkyQ+yn5Ef40yNZbfsidfboTCp0wF1XRfmEl
LR0xIuzwCv0maBpRhe3NMmPcA4SZESRnx+iRLSu9JGohwO95L416HN4qrmM+n42E8hz9AMLU1ase
hmyaWbKOonRrWmTET6JDPmM+HUtRxgeqv4+R26lXiH+H+R0R5HVHJ5x2w6pDUbE+rumEXtHXsMtN
/QLGHc+synfsdptyMwf/s5BZsIFt3EFa8Gnfl7vngcY8tllDSJBtkcu6ZGECI351Mjk/nZhm+6eh
yh+SRbq6XmiKo48k+oJ3Jc+UfMw272Tix2pjepyjBDx4JezstHBePYAXUy0WHqkSv+89Gl3Kz0Lu
A4y0mjkEowwfQ1y0U7STGncUO7hzZ1nlpRY2+KE7dPQ60ZMIr63brNZPA5nGPPzcMEqtVfrYZm1t
yNE/wXPz978hFk45jFCPWs4TMcDGvIkjgL/Oq8rSs1lIkr16DsS4pAuB7sP/E8Ay5M3gD3+/FdEB
i2w2YzsTr6imGGgIx0CswmqZpj2DykP8qOcFYNLbgzMw8Mroa0V/jsiF62n/3O2MMT5XU5Nwliir
kCTK9byOmrvgM1f4NnPER18HY0U6XpGfX8519ziKNAOuwh8ozoLSMltVSz3SA3oyNSnPVe25LUgI
LlNb7B8o7eY3XZ+kDUOl3lwRqT8339zPVhoXvrH3iFIlgKRJvB8Zkax2NiOVbnxGAnOCGURZjJCV
BrgbyEx8TeGCU4SPx9TkG2AnUNaNcLawrJYuNU/IrbrQl8JII/W00EUTkRWAIMdd1wHfhFoXSN5T
5eu+C4M1nTKV/3VZKKqWNvlD9kx8IDWeZ5O4Ja49Ga3D22RMWmYYb9wV1Cqs+wNbPYevvDulgbXI
GyXoO7XfTjR/zv0tlxI3KUR5Qda+toskeUoBQDYmJHfGk9hT0LxXQeF+WlVN1CrG8zqTpRVUjY8P
JmM7vO75oqxtClnDzaZ1YCaI3nsp6wqyEgzGoPrW7jXFKnp+By3B+19vJs2DQcenqs0Pe5oBz7eG
UgobsyOPxxLkRYnxcdoehY7PfxS67zR2yHwrZeaOQNgijO9Nsk8PH+6tfK4gjYNy+7G0yeAxc9NK
vQHf3HvKA9ucivigP5gvJ/0WXwXAjMTyaBdl86xjdBAQ6ePx5iv5TCw41/hF1VdJ9waqcJxwtJoO
ZsoQ6wo4tov2jaPHFyQ/tL25AKwr52pKXfusrqsTf2o7TEfJQ0P65xZfzxbFnT28wGsjTxda2kLu
SZvr+NvaMB6c/c/B34Q8L2NIBhZJou7877tc9vl//mzLgq07Eagtl5KPzuC71JYZhtAbLagJaFzX
hQUAbWhinYpzXCRoLvudSWqcSLC5sWFrwu2NKxRQ32IA8TiA9YFhQJ3Rqpzx0yaXUYMJhrdW5ZvQ
nC9Oah98fGw64q8lfHUGAkxeOS1EmzzuJV40VaEMURMQ21q6mQp5UYeSs3QK6Yy+OA0nL4zgiPog
E/CV4ZizT6tlazYTohCKWuGq+lp6kpLcJJDyNN2lKFeon5EU0hKbU7XEipMx9yQ3b5PBXMMWKCA7
cJBq1IgdNdjRYykifUcHU/2nboXt9aCPeV2HSVw+EQZCERXMMIiONuCStNGbu3VkPANT3ZvOObe+
wASj15xYCIkwvRob6g3P0gIuyGml4auVDNlJ75Z1bRaQgDwFQzid0ebWB7EhDJ9vW6adaO9ovsXt
gFh26oWZIgJDra2Z9HIR+F3SO5/gL400zeD8LKpY4whonI/RtEx3q7eX4Rj6nN83CKo0UXkOyK94
gciBTJPC+oL+mIfy04KwLHmo9lj7izFeSwsVAaSGznnNgNEcWEul7eSGWik0h0/nS+0BtomLpwsh
vMpUTMsKyxR1B8lu22cFnvediKVPhas7Yf/DDZ5Wo298a0ypMEwPfMecgzpukZ2IenLMN2mcKtuk
uZHOK29AQVy1kv/UUoxLkDR+0C1LxRaIcftKlKLCxe0ORpT1qXdpj2QsPm+jjLaU8uXoITzlqpTa
NiolviFq/yVZVLDRQQIHVsaLzlrz32IN30FvaKJxbx8zxsvMtpIEExC+rOKX41v/xotrAVQ6G7nA
eGxwlVFtsVdkMlp6afLjy3eqwTSWbaX+4BYZnb2dWLfRtOJPixBjUbW9vlwrhm5EYYO46l2Numju
viljTB1GD8oupu4BO8exGfUwfj6Tvm+wrPt76PFlrHDV9fLe/vigFlfXgMqPUntgyL92/NV5A2HF
EjHwDgxddPQ+p42p+9iL8nR8nTBaB82b92mJ1gtKHK3TJGFeGTbZHqeRke/LFTycH30OS/utzbdS
sbX+kLJAKZtkCaLllOmAV9v0uYKcLl4Aw58Q7PR1i4ylHGB1yOWdjKz/GJmaLpK37ZlxnIXhv51y
wKdDjdprzlsP0tevdzOBo5pBLU5YyUvavBUEZiPM4nbMuAUvQVujEcrBO9459wEwAJFGCg5QMjif
shKdyLC5r3OgNigZ3RDNlBgJxA4XM6yPaMZM1V8YYIN/ZudtKern7eh6CO1c1GSviodbLxfYkVkv
zv4Dw9yxC8hcisoR5Q8ZX0PIc+8GmSe8UnUtS2CCRsB5u9/SWjK6xOJiDfeSE6zkXLsxH3kSoKlM
g+i4opgYdfetkPOsNjnyPYlw3FzycwNLKg9JkI5TtkxLRBOKS2W0uwbpq70RkPrVuMydDYWQX+BA
zVFdMKMd6HMPA8+GlplJDbovnJxOcskTck3dMsFfyvl0KAz5XAUqijmq0qetVZS9aGHKvTODQNhk
zO1XQnn6tf7vk6J/0f0tUhQoWGZiERA0jmP28bRxcU96Ud85+ZyMd1QdvDR/hpkVcCZXpmI98pwc
6K+2xpS9JsW8aeGDixUbT+GlAc1mYzJGBqBJQT9QpNsIGX1cHqQzabnC2ZqSdGs6jjvfFrKJ+eKD
vrnQVYFxml+7yD23qM3Gsv+CMB31c77yUT4/diA/NNJpB700lYF/jQmUquevxKK0FAHwlMS/JhmT
3ciBBZMbwb/FrezDw8FAEjpYHPvJEJSJhrSDFZxCEo0aBaNRPrU9sgbA8Z0R8HPi5cnSiIO/a+I3
SwIXoqeX+FvuaxZSeI2vQqFOZuQdPvBohq3cTUOmzK1a/gjOiZeecRdnl9DHvjSEOiy9fUqvsTLH
RpJXtsmJjhKv+aKrsNOKjcLq8o0sM1nNw1PrRoKjjyA11uWnlsk/xpOP67WoU2k6gE50zXDysZy2
jWE3NUald7Su4d/y2IXNwdLLlogPgRAHs5/R01jSAq+CBT+xW83p78cVqPhE0tGixZnGvpp2PiQL
y6tiVTPm8MPHRO/EJpnXn7XtdPhEdCifTkjUC/5E595QmD4blSVeLxVDZVEXzJDG6Ad+3s93Nui9
WfEa03hNg6bI93qrta8Th2tUpJQNibOUmRtke694X3EsXlukGjUTf3k/whMHKTdQ6KroijCsGY2n
vgW8XqFWCYnijFwsYvxACGVgWQBlTcO72+jtKnt1toCQVeidEUiex05NBkm8/Gt93FkzI9DxdOig
ZJ6ZIHcm2v4Nbc66/LWdmaUhIgSdajay4pQLhhLhrlSt0hfMVitZ2iBlsCAQB+1ygNveCwvgdKmV
SC5ltWVpfLAQPddSoVGjohI+54euB7AyxvMjIeMMwLhBIIxTNMJh55kcRYqF3gj874YDrs4sMFqa
3cHib/U21EFQBz9xrF3n/80jTBcKpJhih/s/512SgmNwVqDhji/Y0+jTXuBaNjML9prRq3U/y+Zl
awW/7GrhNGzRQmUt3Sq8PHqRkX2O8YOe/3wM6KQ00Ct1KCTJB3sev2beQUASeJ7yEb24cPQdfNq6
JSEMzojbm1jOYpyfTm0YaeE24KS+FcEdqHofPAyyhlAMdNYXFdgTiPMcHYsGdoa2zg8k0BzJX8Zu
m7UQBE0RomhP
`pragma protect end_protected
