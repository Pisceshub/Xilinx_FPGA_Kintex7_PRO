`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7216)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NxONQpWmaioFGzw5JY31JROm4p5CSArg0a7
BZU4c5xmxSJJ0wmyjegkSDMplKNUmG7wxeavcDKpp3nDiyd3K3hxhwMHyt+Wm72G5CehELKD3CEm
6I/wISK113PiipMzQL+PDzNWekLBeWhNeG/Kq6pEEBqU9Z7e5njz2TugjwecqNvOMrGhoo01XN2f
UB3/esxiTI4bZO/PAXFXC0S8vS0Hf0vCscdGxAhjyWnewoVYMg+Gf6rK9GPGEBDplHWOa43K0X5D
z1Ucgpl+t5DuuAgvCeoWedH4zNGCKcjAykWPb5IV3xAuoEDcbZqjNtv2kTs0dHEQTbUrIFj6lddw
GthhqYvu1KK8u5TrQxQak5VgqIoKwMNZyClL7j+yNxpYH9F8qAMMlH9jVIkQ7Wa/glgwq4abv5wP
ja8HgaG0hMxkomK+ib6E2mfDBO9+zI/SX3ErEpt6xz94i3CYmtT6P+NPpOTiQcy9Taf6yqvwxN1p
ZUhqCjii73TAG3XBhrckW30Nrki2gh9fiVCnZfAnxP23jpmTS9zRgbsliujCQ0IQu7UhM2nC4b24
n459KqkmcS6eIZSdoy+KaqfQGT99qFMWh6VwdgYrmnDgbW/MgCs6JQmbJlBqrwlKLqHGVpNQ8Ww0
ejd4+0oFtGWVPFfzP391DOYlpnNEFvvx4R1lv5amVj9L0Ko7qkUoTBHkGgdjZKuRurkh1+OgnHFF
6uJrqX3KLpd65uugp0iHcmZzopd/dBkgact73GnlfGP+w1bp9vEGI0I2nrfNpVB0uJRptpfO4CEd
TbCgc09Pd7F+9izle8BJ28hrH3l5hswrl08bJ6d157PaZTfZE3tk91dHjnMGaH2FGBx/0QWFanu5
zoS1UsUA7GR+KxVXAkIQQbKw3Svt8uHCWSXwHhvHsWPYzgqZbevOq+W3tMDtLwVjTqZ2yAcNjkba
9/172ryWBLiYuRsOkujJhccLGg8KYGWmmBY3wxq1v8fOcz6k6/Q0iIuMbXWDXUdnS6XupiWS4RH2
HJD23By/b3VwGqXggAhzcxIyPUyt/y5a2G6TNTIPUP9wrV0Ku6X6xUmhHvETPkX3bw46HE0Rg2kq
GU7t/pvn4hWQyqtG7T7y7J8NjFj5vUx1jufvt8xZELAQy8w/o8ysEoXPkA4xx+EMP6pP8Yc0u4uJ
q87SR7SypvbX9NvspbTDPiyqc1nmrkrFcstAKgeNNykCGRjeSE6CnEDJ3e/0VPFQGzY45DrSUmn/
E/wmK/3/N9WgRxGsJ1xeR/Fsvlu5O/Yc1xlSBHI3eQ+iLVmadi77oWbiapif2hIR6RVdFiY1pbnU
X+UW1MtFwf3YbRpU9Q/YPnCWHiXXaLefHLgVgmsF2YGAqJawncqTC7iNaQUESA/+87W7EBVWbVSj
HRXKupv8F6cLynwHL5j1nAD/3BT5SbnFdanzwuESo42gYxhEQqR38DC43ob8Bvcp5oZa11aPZ/oX
e+xdUEf69/RpuIYG+h34RXtq3z+J4FgQEx/grIl0MPJpf+wWo6TJkjxuVQEri5xDGcPWoOuAxwEl
NEia2pQ2JXshhxnRM5wmypHDk/mCLx+1rFKHM5htnxqyZ/OBS1uTMq6x0K6pPGcvZOvHap8qCVJH
9UdKx8TTd65SjKMwS9X4vnF8HbIKQ/P3FyaA9YC1SB4fiWJ33YoeLcPSOfyRfN1uRiNJbNs/DWPX
kv6Y+eb8WVcb8UFZVtzzEXyaVJjyynlKhM9nO/r7CquH8jKzAE+ms6orb6YhtSsNxQV+PdY1n+SV
Hym8QGWUO0ZNijREY3lIvrC4lC/P5kOzG+VnYKrfX6+pSDSbmoR+z1i1tMznPQGNRDUb3bS0Fe4O
Q9ia9N1oTt6r1tlGjrko7r1QfxZ4SCdgo7qilNIGz1BqffNugincZy6laEHUZ2BCOoGKHNHkJvnW
V6EcsELDFznhwrNkuo+b6/QkwKkePx6n2vnZGFqZe7WFddXUBgYWMNtIvHClFxFtvDX5HWfYhQe+
sMtb3HSKFODPppqzlD6AOrzyOEHafVBRYFhRmVi/2bGzHz/1x54Xo4I+FP06raBvTUyww6O5+Gje
+aoJ+mHPXnsNUvPqT5v9NKNsOFeigxVuwkY9QAGEHchD0StbiMOa5QkogAZhMSHWdyAuWRnafrnn
UxcjY7W8MXdbsn6agL/2Qam+bH/4eBUCHW/pTPSZwcILq1XTZf3brV53th9m5akyvvu/dj6Xd3JN
BdPh15i0NV7JwjIvxywHLXJ7WY+O2Bh96Ereisdyf1iSpUNID9MvcgC9puqsJ8SvNfkAY/1j74ul
hh6olU21jC/a0pVtWWQjA7EpwXGmOUUjnv4k9q0MqiGFNE66YFFvcHDOKXbMk6besk7w1+CVbU5L
m7yNzCQmyDQr4V0zR+69jYAapRpaA9p32S0aUoz5GBg/HOPvCmYU0oDvx1Wqjh5YS41drtoM+mIM
Wfh8Uhm1E/rCrMoaDzuSUjXRychXYMjzCElI7GHCJScUVI8T9S8jlKN2rZ1LBISgtcLA1WPJpVoA
zSWjEUHU+BvdHSvi0YN5LZjvG2971jyizF/4swuGp3u4vmagC+il44QLfjHu7uWlI7biYvTICCpC
Fldo1jG/do/Q5eRVY0MUs8D59jwuJwir8YhXf6BZPHsaORa09E3rHxPkgbRmiHodHG2E6PFs5gfK
9gPFD6bXd8L9VDBNmXH5qO9dndU8elgc1/a/IYaVy5E1C8LQwNybIFgWgCa6w8DMGX4bSF6z4Wju
pI80RzJYzrigGHpilvlKzwKT+udsFAkc3eEAgVzYjE4PFg+TkHo4IHaV+MbML0bSTQpEKt5+8j/v
XTGwr5D21Nfxy+hI7IkgB1WnKNop5jkzsDrwTr6cKqroUL4MqTHd8Td7ZsCZLBTl2nT0kvYFAdNf
XzkcgjoS+82oNIQvGdZn4u3w4qAlKwIM2mHag4VmW3lml5aA2t3Y7LWdPrYCR339Kyybp4FE/AVs
5fkGs6IK3piyc/ZNFXcwy0tzIj94iHO5lrshoKTPJiViZ88wAGoS8POOgHINDUV2wsO0wKHncM9R
SRxtzwJcAXXPT38kHVCClru5tNa9PN7ahS/0HiP5lU4ILrlZ+SQzcY1dHJL/LgPA03V9fCA3mu0A
WvYjWftf0Sj0Y5Zt+ryreAzTkitaQ9ZTXWa8aE5tQBEEhupAvwgmgomisBhcCzT7Ey6NO52M0l5n
eOpfO7n5VtacQLGL3Q5QuGTtkwpO1Um+rXKl5QKIiuSOdX2Wrj6ezHXWmKga64Xk2wedwCam782q
0ufVpzT8wk8NA6J42fO1zFpi6v4gu0CtJZI3fdk4+G0HXy34BY6yTthWmf3h3GY8Yu0MGw9k8SNX
FJzkvvvmyWNuKgS6FSR0PWxch3QnBwsM12qPtlUGE9OHz77UOlfCuYOSnCOkG2OGQcd5RjSTffR8
w+LBaipx/RKCn1NWP2N1J8WzSvIKw4TrHFyZwsRGRR5S1vETac75HJDUFKwuFjOFEbb+5j17DnL7
ZD5VFfZzFgrNtN1lBxKxpzZ+6d500HlMLuGFBFLUMwqeII71ghsR+G2SOBbyGeZo2oAcnpf5GcXw
YvSl3JkWaeYQFAI82pamCRDocbCngc+NVCxS1TVtUWfMSW3BmSCXvCc1OzF5kS3Soifsr7bMd99j
QtQRXC3lU6cadMwPjVcKGuXxDQn40wPbMfqUrV7VT7D48NVLH3Fmf1LKaBWOoEbjobh+KS8cBWDq
Gn4S173+tlP3fRI0+LtB/Rbi97ScASTSuZMPSyRoIHq0nKUH4PVmj6NGft8GHTptNe2Tj1231Zaf
mmkZk0JrXWgLg746MGlBtH7ezeyKAa1MYL1Gu8DQufGKApGh1xA3pehhsvuzMHJnGULyG1urrL9s
IhBwj78PD4U1C0F9nK24iDzXA75OvvyRrncn52RQBA1TCFpuzI8JnojtOpBQkbuP0ffTbY2HYim7
93/ZXhKjLlrRLCgwS8wd9fzkYmfUCg0BRGLS2/snY0Vssdh2Efrpv0unhYgULkCN7xAXeailRGSb
+rOoguG0KemuREHdWmGzkt4biBmGFF10UW7XukuJDuqjD4vVsK1AzGpNnt4DxJzJ7GIDUFpAbjSu
6Qgy+wVFNhe/mz5k1ZoFzLlcRvY4ySuuFo/FDo4JuflTbv7DqrKhZWzamKPRdDe+iVcesyZiRhc6
yk8b7TaTyojdqFM1bu9SY++x5ObXnvnZqj4sE3ni5DaOAmqGDEjk5YNAt5RnlYXRikZfAb+Ah7q4
fhxbZvJ8CGwLbwf650EUGVmGtowXpG5tM+8iYdi+k18zTdRXXI9MSj2qm5o/FfTYfAgt8j0QWuKw
w17b2ZDHzbC3ahH12hu4kd+LqYh2dWgpIagek3HffqDVfgSYqbXNaeT6thKnhnw/JNS2dArAsvBY
lj4ekThP+RwzM5whwa8d6oDwF01/IDxg4+0NQzxbD3y10p6ryuX4EyE1vU8xr31ICI1HLmjMxWXj
mLwhtSn/pMkdga0Wbp/j/jj7ZTRDk9y8fhDt9Ko47SywH+zf5lJq53Ssgt568h3ifXGpablHd6Y+
npf0+4fUpZEs3rw9ta6TB7n47wXI6llnAgX7o+0rGCYb5uLCZ8aXenOU6TsA6kxwCXCxUscHt5mx
3I6VPOTCYjrDYGVQsVLwAMxPsvmKpPDp0M4VaKzIpliZr8/onRcmXfnH7FaLuMIq5zmxjsn00dJL
sS52ewpafQVY4n6Bfe6O8uEUnhJRb9wUgU7TBg5S5AwG1XqCy9NFF7ZG3gjI6gONC0vlXDSl6hqu
ww2jukyc/ZWhqGCGAhEHCby8RSMDglca0O54/ETwhBJZuqlvQAEsuaUrw/ZQfvQV/ZqSljcIaC8l
LStkzWu2TYs9p8w92LS2Gq12LMMnvkJ1FqSq0kIy1o0K5o/S/E1lFko9+i+ppBppT9yfzcp8zoSE
85QVJOSBHithre3Kih50eegeKdkTvhZYbnA5kEFi7LSf0lTFMRpIKZN5cYEzjDwgOX5Vxp+BKnMz
N2ODS95jvkrOUyFaURBWdGaMQLex2ZLfwTsEYqfyZOtDwtzdfekvCan8AYWVnEkKfwjpEggI7nlV
Q0tXbYhrUQVP2oH0WiKrJ9WHCAWlM11Mljb3xdKhpHeBrakGlrEL+A4irwDcV2g+BQXLt3B/O1qG
zmn5FDIApwpXwxmJtvDIqGeb9OQPdiAH4ywO8hwdxE7SkXNlAx1Ypx2iFlSZKgHnvtXKdR4ZuHmg
zqxprjrJ57I6Qh/01mVLmpPo7MV9YEIrcKTq5xWXRWcDzRICdQ1g6yaJVHf+1G9XHCRS9rtaDm2Z
TFVpydqKG1THB3ItFIgV5Z8Vw9CabBM5rVaR4H3PDVWmU7o9l4Wtv6t4MDJnwfahb7W81BItDmha
WqCSTLdhTbIcaub3EeVU1PS4jX9pft6Q6iOtKBYj9IsMYFw60XbvBQ33Ud8KK1/FK2kIpEj9UXVk
AW78KtYZ8Eg7SmWXFEIxSdboplwe2SvvrOV1FTwZGyvN2noyyMHt195H9/U1E8vi+FokVZwAC0sF
2foAplxfzC7AFd9pK3fj/xDke5hMzFIc+qqJtoXAKv2ZYgdEUB33GoQLgUj+Ew6/NzTC9VubjH2T
azqunppmswfKU4mDtiwFrYgPyi7t3q0V7MrVVG5TdmacTINFYW6/TQLRTgOcOCTWt9Lbbe0IMBHK
KCvC82jEPAr+OSOx5PIXaUKlUGzY4vBZTMiSIrWW2JWQRy7VpOjHid31u8TcsFgCyXVDRkPmyuCK
CxzTUA2BqOVLFl8b71S4JAKnZBgioJHU0PTtmh4nm6XeK60dULe6OqG80mDZRqpigPk/OgpxCMrZ
/TwiujZ8/uGQZdImqoOmuV8WjnbMRY/iQI2qe0hZBKmTOcLtdjBnuix2FSzICyNIEEmypr/osvI7
fiNocOYW9YMebuq3yue4YCa5xT3RPSfcxCKTIXap82G7pZHM7to0ykHAGSioSiiY1ZILVCebBK2P
637mxkor6YNUihVtqLfh1VmgWOJ3IaeOHHRhB7pkz9KOrZMc+ZrCNEYUPOVmwwhyZDEt0HiVGV6g
3z0Qc3tpRJ4JJ0D5+kkQ+YPCUQO6e2wfgl5L8SHUGLK+6m7HhsR/Hf1+k5820mfT7Gn3nsOWD495
kPOOplOECj8sYpKOJJ+TFWQgjzUF/viUmnzAUtHhNIlYzyBdSdTOp0UJ5rGjDhdCCOvNQoRwVtXT
ANLSUOfHzfj1sko4HjWgpXqgzqCeouPfijqFLjVfF+dvaDOSs1VJEkZwjU3jfBWMVvRlHEDRIjr/
7T+S2CVcYOPk0GfAJ+27Mmngicm4Lo4kk6xBvDhRgfpyfuTr1K/KGc73+6SzEV+nKO454ytQ0NjV
/ot0jl3gJTOb67YAfMEoytZkumB6MIP+8Jl92nX/Wa+qlo8tzsBW/RRfwkgMIxzG2qLbxryz3sYp
zmBYKE/mc57QFxFfxtBo6uf3d134r61JJZ2VCSPrH8zO3z0B/acutm+E7VNDT/83/sYNMq8oBZSD
xkTIpqJ0rUNzjd6XqF+FcSOqzyt3oxIh1GSfFRU9OFvffvAlsbgftzL0BKMzYJYlznXk6wnjQplR
r33I/MpztUK87Lf/7dqyTO7Eorbok5o3sw8NJoXSHmrQexUmytPt59uKE217018njLd7DUepWiJe
Uj1E78Mbt4NTqH+YdU6MoALs6tWo6xGZnpgCP5JiblQ8pc3rQZmk2KmHxtK0xGZN5sXNq/nD7iiI
hxJt2AomXOt1dcQyh5kGWSnOj0s64ZmDe5lSEjofjGlVDHEw2FNqUNAtxvvGD6+XqyPfG7C3sMRD
YM3pAmYWYs1jq2tdjWjJPih4ccXwR1cmPeky1Qqs/0yqQKNzgxCe2WUIAJy6FkM9J/dsW0I76O44
cqSMpfOVxX5hc75ramMRkqFub/3zb+ZJNVVdVJ8wE8aPVp+k0AFYOU95nN5THJEJhXVGxifDG+/h
SM1IpLMMCTQ34X6TitVh9OwlvncHQZlc+D5FOVwaj8JYaAhgBiskOGtCTchYh0IIOxNr3U6iT5Xa
+xMKjMw663tupnCXk5kXV2ymxn0du82kpTUttlMHDRd3IuK8of3LViqJZyU2HactZ1CmNQP4NAL+
nE9sFsbCHyzrfpps+ry3mblNLNDOptiKt+cReTnIrvWBMPRE8LA8Vk559Y692DnhXyygjmwAB0H4
MBAKkmrmCq2Ctd2vodG3GI3I6W8SyLwK77OOSAkP43k3Q74NQ/E7tVTijPiPvkmXGDJQMJssYPWE
PP52WxH51aB09FiJGac3VLtMZKQuF+AapqqX9cqHKw3XcLb4n44dgXw7zi2VbpqaLYKxYQZvXwvm
wivlfnDPlyCovJKM2/oMqKSEK3Ij9BoCKqBdu1oj6TBGyzRHiq80NTgkaA7RXrhuahZwhMHv6bl+
0j4E8BEiyIflrluqx/xq6ByUjj7Gqfdfs+z1QXZxKHyhRFlxovzRGSdGCWRUBAzMcnjBDRmMW1Bb
/1bJzuRmtl0jW7PYfrvLVCTOPwhehdAkgbBtOjW7G6l9/8RzjdAX7XaLLHPD2w+9LVNAjkxe1l29
s9dIU3aHOUAEMTxvCOxNfqu6DwzVteVINvWDs5sWTnHYpf2VDvrWrO9zLUqY3RuuB4I1p3abg/pZ
C+/auFXvR7W4UezVpS0hTLYaqKyTSW0DmlEp/e2ISJf/vYyniWQmbkZM/G72eGxFd8b2J3TeEg0I
B+IMZMEszbwFT5Brh5lpGsc4jwucZHsZI9wu/BCSkWmozrDiDzNMSXWGTTtXpPwt2Ba73+iROhI4
CP4zcS48QmSDSSvD9cP4e4XyDoBuYyZ69UXWTcEqM8lTGOXy8L6861DXXh5hEBrABVil1zchozty
zyOLyaCDn0LHhdCInEg8Zk5uPPskkfu5sLmXuMU8+4hQLBCG7Fl/wNLAOEuqyWQsPaaeaiWm8XzN
X7AlmBEUtMB8ghIjIAkpQI7yA8FOi7CmtQvg35STW/1EnuyGm0pF02jBRs3NVk3+Z8LNfLcblX7t
6oPhg1aE1RQXzG2cHsBEqXiyvU2O8nfUmj9KsxKdkDKyf1RN6GU21NPN34A0yaFki+dfBEe7iIye
imgVnXPVr+dt+7dxoksr15AkXEU7G3xLYo2VfkabS9yhjG4Bzz+C6Q4T/scsT23LO+0W2W3Nf7g0
+i30RO6FCNzqu4ZxCIcMtua23IQAbR+nqKL/z/TtMNqnQE07lfVvGTBRSxI6zibT4orT2r44h9no
bzdvMMFEEUD/uDzpCdtu4CW/VrXJHxDI6BEFXMGyULd9ccNuklVbYXtvTRSTyCuBW/3jt458T0Cx
/4037+B8T631s/0RtZsIYLcpbiXFkokcelz5+SfOGIP/Byb1NcEkredSj5Q2iSBMtgyQ0Tjj7vj2
ZacAV0Or0+HXZVAI6FB4wDO3hd0XVxzoleKvrQmIsMNhqs572eJ2MxZh06jgNTydw+MOQ337U1gB
H5Wf0JhMbtVftZSO3wuNC7LprS6EQhyF47jt1ju6NmZTM7H1BC7cYs7FFkMNRCOKMOQA1a23RO/W
0KtFynT7OtBagPlcFbR+88GMoFa7FZtb5dV3ZceYPzPSZK+QQwwDdP5JXfdPNnjkw8glehZTEgZq
Ug1GWJJ6PL/QVAIBQth4Qz/Oy27QprCW+H/GC6Dt1LWaj31adQH6G0rUfpztWyq/PckiHfTM/n+M
czoB6N8q6uchWYSu/nCVrOEJpAmbIrr479O/VbJMy61f4+De4psHNRgimbYtI5P/OARroFwhaBAd
zuxoSvWLWZ8twph2HllmINI4UhdDJ/9svNfWCc3Pjy3KmEDDqrj8TIKGxMQjoeyiAYcPjB5wmMyr
XLCEv2wQpuKI60lYa8bQbVuMP8rQJ1UAgOGbXDPCBt+miDD/rintoh072UqbCfWA0TagJ8oCOYNK
K1b4rWA7owpQIHChRgP7DL/NRaivGPz0qIy0hNBPE8fJSykrnvNMRVThbK/drY0q9T7YPZocgyiR
qfo1YXucVNw7JYwOBSrd5UDw42tZthQ3h7iULzTp7Ze2uGHzvzNph+ZnCp/B8SqNqpP6WTZzVYwD
E1crJtIpJ0FIXvJLtLfZja6xXRnq9uBh0k8sd1GDKpeGHQrTTVRKScpZsL1Nn6JChtfFwVaW2z8d
+19ANhxBzb8fF3wfYWGlilcCeOWAAucY4wWEWzIdNPs7+PuFPMSk7sb59055d3OR3dWAjyxdnIEY
15uIxNDudFrj+zu3RPCw4PT7zEt8YgVBi6oyhCKKe2nQgE0qZUB+OnwrScczS13Kl0Sjhkx96sys
5bKkwG1D9YZSJQfX7x4rM4D/wKN+cT+nBSesWya+4LN6FW7OGrAu4pEGZnCV9A1tUo+jtAiv4+BR
nDMiQAGJLeI76U5TtO5Ihdasw2bBBkbbF1Xn7hXMvpvDwKaJzjGrYRirzv/vPkLy+571reKtS+DZ
gcgwM1U9tUVUsLoFO7zeZRvjjnscxQk9B8NOxaaUUDLc4Q==
`pragma protect end_protected
