`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
3dBDzv38LYSblodwRBnvELFvDdbusrdJTfgKFrtmuyDHZJqY0n/3gCxtINfzRjq1tzcaSksr0Gkl
vto0VpHB1MYe8V7cg4tQsMYUauGz0ETmXnLEhL1mN7GYsFqHyBHLsmacwbDghmweTAc/SnDAzy78
GS9z/2HtK3o0eaLv/xAzX/wBE+lfBiSvu07LpGa5sjyZLvFZudo8AWGBwZwU0ufZLLOWOAWv7uqC
BTvsc0DbNQ0iW6iWxB+UW6VbEgJS+fY02tiN7GK/PSno7nYzADSXSwk3K0Rx+Gxtaj9jm+d1b0ju
SiXqegtmCTUrt/JhmG29seyUbSU9gIU2Gtg6sUUmJXXX1u2FaXBmMswOEVUIj0uDYrK+GLz0DZqn
vNmGMTzaEgVjkjuzYlt4TVEDeTgDYbmJ/kJChYXtXtiFiitErZproHtYrYYAbW6hWsh990HZaX7T
5fSEg0w+kNHdZD+UN5eNHCwk6Hkh6Adp01jAOPt3gqhT+Ula7iKuI1Ds4yIQzRhfZ65+hAJRHKLq
5TfA4Gt7yWSGGt2bL5EFB4PMmYFry+3fPm3lV51EwCi4tfDX9k5r4VTu4yBfNfPB9MxLmLIKMzDS
D4wVsDqaaOYbd6qemSAs4UqYwWM7JBbaVZVgQm6TSs/WRKz6fFy6PBq32a8FPoE1u++vfQTVZRAD
+FFW103iGQbR44u6MaA3ppbKbV0K1dgG13YxsKkAycLx89f04Gsfs9ydLUL2hjHvBN1Hjz11Ohna
73SSJZxdWoNDhrNalYiuamV+daObSRCv2toFG63jKVyvd6gLOWh0Va2yO3KD/xjldjJ+6em6mr/L
Ff82fC7D+71U/IJEqAZlNmQiOVGwa2bZJO3hxrwTY7hNg7QBE8MxtGe/QZlPBUuaAgnm3ds3OI1Y
s7jSipsXYgwUzvvMVcsWky4x6Ad91U4T/kxoPXTz1V+FyrCC/Bx9yLpifl/Ab5bXZB+7p2dBr596
BSnf4fpIJTjv/jIexjNIFiMujtGpLAZ94P4bEhJNw1qjASd5t6v078r49WzMhX6Vw9mUfkTWc6mT
Q9jPt9BoNGCeJJTHd1ltZTXiVDlc037MD0XDZUzmaVcdr8I5fu88KXZV9tVQxbmuIkZsyZvC+Nhx
kpaL2CnACQzNi12ok1mQItmfDGIYP+HlMjTsARNlMG829Ea+IQftuHbMXih3I8Xu20wrBe0nbWBF
NarmQ1qVG3gOTCguo1BBF0rVfl6PRo8YV/HV/pP6Ui+NmPJnvCr+VD9F+vmYpfcxWfLIvoC0g7ZR
ZsQjCyPW0WUtR6v7+GAaW2QdXvxyXgUP/yqzNCJW2K+YztgSjAUGhegRb6Ki9jzlF9ybXjXzNqnc
bguF/tGpCQ8av250Iqq0iUrX99NvWotpdG76wMpplrQn21LAeXbvE32wO/vDxd3+IG/bx2W6zkwl
lq50ttGjNwwUrGWZHkNIyorZcnD5p+/z/9jiJqjs22FoT3AI0Jt8h2tNViG+f0OZxibc4wyI/7G+
qBdAlx2KmGOElNI7N7O4VF8C0fJ2zvusE8xGiGmWMl7s1QpBWAec3/jrGECC42MjcxUasvkoGqDx
E/78GbCI2/iq+IapGiiC+Lt970JDVG9cl6DMss4gZyFBv8++tg7r9PlH1gs48P1JEATMQmifC/jj
tn/M3SZe8G7W5DfCyLCfsRd/s2SvXoC653x90+idA5iR/vCfVZaZAmvXogPYtBwEYEUoheIliMoz
3Oqe6FbUkScPUdSG9nvEHi9UFqSKnYSVpGr7u/o7qN0v5hl27+iPc3XuhRLhVIfPraDtxOXD4BL+
Gaw2YEUCUfW5IksQS79uPunnRpLkmTQkCZo1prt3uEc+R3SxQFxrnz99hXwzYRc9q3lcRw7SdMK1
yEKUfMB330wEhHDb4upQ4nRiTOZuvwkCPeqRUVZonKPraZXZWvj+OHEV/fsg4wFN6nlf9Gr8dvKo
QOtyXSPiakfEaMybl6N0x6kWM/nds5v6FTZE85RYAPK9MQvgLqDi2l85ofwxxprWKeH5vArxOPxp
+LJqLIDWYxacvDDh2Hw4eGOItElbf79ud6EjzcZUOXBiciYZx4zEuXpqrL8E/nB48eVvUfGGHBxl
XNWMhi7tHoe6jJsXM2GuH9LFRtNbYyKgpGgwALPaKfk1r6lHtHDsu8nLHX9ubE678MMlB9bsoKir
LHR/BiVaDasTz81BWAV+ZdNr1/9I3yCU68VCWoDhU9OYLLjPqYVP23SYDSGEhJTFKIrlQUF8SM7Z
5q5S1389aySxERCD8+oimW5r41lCsApUnhhlIUQl0hsLmwhh1ANHHqINMWLf2jQzfpPb7IPfUcgc
9hveNhekF/Y6FCTo7x9WevvtxC2z+yl8TfGHgVJjm6auJOZl2ZWKm6cQwNXNKxKnRFNbvoUC5ZMi
OKHh0Bh6+W931bbmXTAsRjUMkorNjMo3r3sXy3PBG/zI2BB8iHlSi/KekDc9daYp20UoYbzSLp7F
FL+abO+/JCWtr0srNqJ01DgEY2J/ju0thtrbB6ZFK8JAYMwFwLUxMcoxKplRc6Qov8LL8fmAYNXT
0xs3TI5KZFk7dbN2lACaDVft2PJmH0bKe/F0vL9w8KEdCgkPfmHiRAUTHW3KrDA90pJ8jG7zWVNT
lR3nongCdJelOaP2w61nP4roxdGu2DcQDIaV0nxvQ2ZTHKK7PkTK9GgF/LbbMUssO1pjoA6jfBCV
7ZMy5DzN7q+0ifV4MMnMfP12gJy4WxomKS8zECarenJyH4pskYKasiF9v+AQFM6H5Esvv9ilXnJN
0JS3Ta/988TTikx/zyx+ur9bcBz/MoM88MZZeirO87uGhjk2oF1K8BYDzeycEYLgnoYsGkb0+TiZ
ciUGx/3zR4BK6K5KZQ1D5lM+QjgfMUxELWSJ+6QGj1TcotWUdbjVZJgUXKqx/1TEWyHCnUL0c/JY
Jf63GIiKXsev21Yf2jhto2n0myH3DkjK04FGPii4bN+rUqfBAJS/GLL3ZdoCU1RRrwn3g2Er5c57
6uWtghtktyl+mu1AJvKMw0aXOPZryh16lt3VsASHVp4Nh1P1cgw9pleqRFyw7UWT5LfaLq0L8j2H
tiecs8C48Wu5IIqQB5AJm5+UVLhpLNx+KeOS7LRIlonv+dA7RZACu+jEwf6HkttAS4Q4DkwqBqM6
86Ja++sAVgy0pJ6u6jg7dnFKshNk+EAs/9kbfhLDkBXrEXvI0ap/QO8VThad803uLHQS+Ur5tAfh
MwYJA588ozMxfVxV092HZXrbiESjqCmNJsgoRx794kcT5ZGCC4hTRUpCyNC+Bn3XKeh88cFet3Cw
FSCVzWLmM50F48pR2a+WeO8S0GfI17gCB6l7lyL7lC6km903a/bQWfMr01TfzEfdWtK1VT2egLxT
U9vLdGGAvC6E/B9/3cJ62KI8eCignp/GcqDiicLMePcWFQiZp6TzGYgJX+VIDh7BgqdihUG2cl88
B4RZkxocxbPX00IGn7/WkjNvUj6A4SqIYTUCYcTWNb7ozTCXOnS+Z7BxhFEF1xhwJVvvBFMy4YrM
whFfvRRK29jHn6GPuRW8BdhQTp6U4/KJQcURm9Lrqnx68dP9Dk8+TCl++LGz8Z07qsBhb61mGFUM
7FEPCLoyI6NFIZRWBGFwSHw448uRu6/kVpx4FZbFooKKQMW4MYz8FddNtaI8BaKoShorgxrykh9T
rE1Rqbxg2Da5+I4LWhyEzBSQ1O5dqfvKtQdgkKbJV4/6AM5C5YUhXafDmkk9n07JRNn9nzjC43Pk
qxfa+tLBtmQAZNI1F21A5acP+hn/EN/6GXD/8tOy9xBdiYcsBrSp/0MeB5lu8tIuPGGaEBPCBa8v
Z5t7cKDmoOhuio5+x/YYsLPIRrITq0yto+vMCsDHBtnhE+f0pjt7qNUtGO6i6iczEygErsLl01Cm
U2KYDzrxVcvj16HLoeGDnz4v1vtX1aav3zhHoSDsUO4aOaFDIvjjgrLXN+j1bXngRsj6/dhQzhg2
DVm96EE0PwSXElAKhwxHL/G1UJUn6HNWilVkCYOw60Z/zrL2XawxneTSXUDy2gbYI5fm/ZkJemle
biKuuUs69b/WfZGJ20828JyZPrvCS7NjFxDTGTZu0n/omj9iw9Z9yUB/2YDBHGQjuvu4C644g9uJ
qGiwDp3m5XM4aDHp2yorqizQPD4XZM83uXccQREwONJIzCGEFa6RplrM6loqC5qaRHoPeHTF0NLb
PcIg+bJD4FRucO2gVxqT1BgnVqOA0N06FfCz0pvNep8wfml2XXrNERFCiiYFkB6++wzPoxRQFvBa
BJG691W+B67FHZxI158LgDSKfIEXE2zuLKLtMsp7AXLphf10XlJse3RAaXHo0XtQhMM3woFsDFdD
XPjCXltsZ9fZWbwUhPDUWf9RIrJJGE02IxVddQJCh6yEyQBop4k/8bQzMqMovVEluoL1A5MgD/d2
zB+qV+4rFx8r7tTmCOjkVCe6oFinKGPMkLNjmaDNMdpDLuuX3t/+qZNDdyczTL/nfHFqaYdLpg2c
F7JdTCnZTFtvm/+xy+LnnBbgC0anq/b7/A+bEwJ5IQHUFXY+Iui7duJt0VXKCNkYCHkzIPRf4wyH
jLPSDxS3UtaFyUaVO4lH2fTaCtFIOocWMXSC
`pragma protect end_protected
