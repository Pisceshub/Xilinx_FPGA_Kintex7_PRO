`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 86912)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9KNavgxBjecblo7CHyC127uYEg4bpN1lEdaRTtpaTvFL41f/BDAr+Nan
E7Z0/cOCC5sb8jC6NgmV6HNu1f5CHuD6EO1hv4Y/WWgqvJw37EILHeD2i0i/NTWl2OOt3DCve0Xt
hlomq6y6ScCC1Dl93+tJb7XRLQVfG0kcfdu7lASEfDcv84P/1IWyaKxuamzymx8dC12oxLATQGON
fo3ReItyF1FJONagvgkEUyRtUE8a1/KmZR03ymTQ1v2RBz2JnlZZ1jTdIPAikbSTcNVRS0yDRNRM
HCzhZ49cwZG48gWFl/0XhhpWxx92bnNk6P1hN7jMHveoAirai4A3iC4hrpC7unl8GsBz3hJ4/psE
PGlNzC+zzc5QU/up02CkPKGRQXQ75lB5FwP4kMe2pDysJFL6+9vJOF5z6MSXUv+OEKQVdodbBsSF
JuiRGglglOMY/+7tHMzZkmJsJ5415FzneDZpRuc2VBaw0s1kI1Zm0AlMJ/bOIGBrFpUNdp3xM1+3
67/PpJrSOMLpR2peMcOugv2aQHyf7bxQzSwVckpJzCr8yeT6XRNuNNffCUH7nZnZzxeVlAOLRpch
6jBl/u5uC5Yog0u6Xt5fg0p4a1X/whsveArFthuHEJQcubmvebjxqSkp964sK9F4wmPoW2RWFKxj
M56vQL8hpSoXdHduQpYNzHtTJ/iVx9wvmbm3zlxYROKReWbDTlI2Rd2VY0xx0djo6/ZfATJWYGAI
QV8X0M1JcfroDeswCYl9f69JqjIbt1luNrtbL/gbc7fpP4WAwAXZPOi92T1JKXETgE1PIB1JuERM
K0igIhqvlcGwioBqqiYN2gKqRyW3PZNvXHsSgsXlsMABKMjPB+c341wcZoczwivSco8D6Su4Xm9z
rdoVAdsQrGxwloIzdN1ZzUj/cPKdnlzJ3L8FsutUK+BSWzs4fSLSbB+TFRib0YC9o3xuo/0HD2D7
pxTqcW1gMUiMN6LkV+xeCAeW9L+EmkImyWBfAhfoNeE9LeI0iTxJzbXTpOvg54zWc5QNlXBMUkR9
FSlDwfm9ivFM4ISEV79Akg1qFfZkQqf9ZSZiYzlxjpWm5+gyN3tfVcZOaxUT66UzBoqkrMrZfSmi
9VlFeuY+MtzVRADIpa34aFLocBHhB6A3U23ghupiX3NunH8FKkGuNThTtHMkFqiEH5jsmJZz1oyu
FQr91cU+LHxQ1HmKg/YOQAqEYO8NQ5hXo4hxgzvuzBRZrJelLpY5P64y/EErfnFWTyWGLTEwb5Bg
CH0KjLlh4tCJoG/3lM8mT7bHEerB5kdb5QFSxrkofjcavflA+6vCLeu9ryRJKgKzAgL7sbnN3GG5
5YmnVoXzzvrEjzYowrOS6hGgW3osLu/zHnyLRPP/mqr2isqYY33JEPrpvoFdAAy/hHdnOms/DEDe
wV5JWpEmDGg7pnegxFDT53zs3PwWg8qfcFMSnyZ8vGWN4oOUHIJFAsRK9nvAYS1A+6rditPVZzqF
lTiPuRGkrIB1Y4xiLQIKCQQaH3FPIaEDPSfmfAUNzWDTGpfvpV9dcSKwuWddRgmLTLpGZS0UTejy
USz+5U34JgRoPkcUUkQ+LMUujNgLayRZiK19iUP9U+8LN6aMuX2qJ+lYBZAfTbF3y1R0IAPkdOi8
u3ot7NJFEKJux4nU3QmG+HMhjWn3vgwGNPB9r/hdYRdf7ea7AKVq3y5OdeyOsGRd+qQQGdyhHodI
yFxdyPqikWnbnQd47eOTXCpxU5zo1nZO//HPogLEsEgaUAdXyQZehz35agqtuOba3/ghxXdE2Rvc
iAj6yojjaCgQWH2k7Flc7eaw3hhQgJyOprIvmCyXXKfLK75BKRPOuJC4jjXsdPCGHZM0zatZofIm
p8wG0IV0TURubbdKn+hOeMOI5wq39ha8qUCMr+xjV2xBi+tFLX1PX5kt0mqMFes8MtOg+fxPCOuc
HwSr6/Ooai8k6AoOoeAyt9Kdm8hrd11OcRZNbxbcSeuCF9AZLx7mdT1/WON1bkrYdQWLrONgX+Sx
nXEdV1mIML53ATmiLw2roOPpMnohAxLQmpfmnWoXsIIJqUBxGpdRSZBOjF43kdyaOn/Od9qeaHYI
X2wSXxaWbcH28PIDa/bmyxUg8rHmJUenr8I7J8m+TM/+tenYISFzFsv7ocsIR5v4icbVm9+avdaj
G2SvLTpjR7xpqXNEogXYKjs1UnzC1ho+x29OUgZf9CBZEGiK7b7X0saLEHXTragQO1IYdvZt1gNC
pRuilauGp7YL63ziZldJeYA5M+KPoUsBQ84QQWxP7uYaICwAsvRE1N+RSd5Uem3u5kDinYdJQQju
1gAKP2CtOhVi4FIVOkHYOfrILNH821eUSv2tytQBM13e8UEA5W4lmlYzQbbaDYgMnZ2qb/793Reu
/C5xzVJLwecjPKFAC0c2xWu5+/I5ons6x7qgFlSVdNFUtuhZe7LYYv1nbag67LtmZDtzxhe2JAm8
EQ2X2/B9FaQ7HqLhCDBmuLVrKqmAb8vNvGL4HrN3x4KivigczM2Hh0xKPCzNRdq1C5ykbstABKgI
J6tK5XlHmgIQcDa6pCgOWIHAsWUZmfBKUQDUy+KSPAFnXAbhj3HUqA93fezcm5MdKRJwOcPDpU6U
52MZRdoSFbFd8unTRFhp+P95W5WROoEQBfpWyuBxUDqFW7qfCQX05xOZQzz9VwSkwVrFldErAq+Q
6NNq4yjGNbGUxHM+0NqXGmnl1reebxJJwpM9GULW1PDkoVTj7PIF1/qIBC5+xN4FN5NIGVt73Qzp
sYXCgJf70j8uQXePP7rrIcqy4hW2SMjbLpJyqjzaXA2Um8mZlzSFyxL7RTLjZA6rXJbar8bI2GxT
PfgnZrAHodt+x6fD3kKdfmFrW6mCxEj6NYU9XEEr1Gv6K2OnQG/0t1cuQ9mbeoiXOOyqfaYMgrqB
qBKvXDyEQShCQLixNRUkiJFhUDGK5/RM6PD59PDmgAXbdmZZDa+h5iuSCrh8RCsQmnx0R6GqbwfP
K+0gzY4XAVLl5Uwm/7q3YtbZssPvj7OYLDj0Nq6MfqcLBvAEHKZgnERSHwOmL1BGoJjxdK9RI4FZ
hpOqLDyH7jBXx7vTdXjZjp3ccSUm1sTvAeoCPTyBNeUmAfd9LgRBYpTZiIv/yt+SYtnxOAZbXcdr
+b0dL2Gp2rca3pUAYRCcPOVmnxlbGcroolsesYJfOrt43075Cp6mJ2K4CvXBcM3DdZauU3LM23Kh
eCgVVEa39iR5S9VZ+PjWRy6IQPwkKQIQ06/Qu9NRQA+P45klNkn4Zm5yNttTJyzH633vZJT6dm18
pPqIpQabg3CN7OLrPj58gbW0x5A/YCW6tKD+ro6HBT8JgZDz/z8xSJ3vfmHJdIe68kXdB54PkzSX
5n4WiwiQkaWK1FjdYdsEL8zO2PDH4MIZPMFOiTiun7gIzkZdFrUa3be14VmOWl85d+a5nymJxuQD
IBn+ccJ9oIIqytFyTZDiCFBx7sbXO8ZcaHK/ZZBfPaUuNNj2aIHnjpJ8srW4uhKHYXGgp4/88CAw
+XHyh4Lkd57hjfrfqDWvXuz5frNpVXo4JuaCZRC0rFqnj8aiwDf2eYylvGLtxN2ok34ony/Qq0fT
mcTx90z5bawMlhA8oyI8gkFMJ2B3XyrNbUb3tNq0HtwiOScIBs1CeaZxFOV8EBu/wSN/UN6eBp5i
WspCfQ1QPFQP2llz6Jh7s3ZGPTNtceWyumXjv8paD2F91Kli3LXwkjUQioB/Kkho9mnMI7NitLhk
++SrtVv4OWBMaUHwWLhVNXAVCfBdrxeFDHAoyHoVctIgrVkb9SYuxDZEEQu28AjaIUUyDQ0rSg2w
Xd/nYpeozzUkdwPliGBN5JNc1RTuQZO4NLiEsgaEU1R/gTUBHZzBRVom4+qgJRu1fKlkoTkG1TvJ
kF4WRnRi0m16e5F2s22KOg9KXwLivALq7TH9CzmZZB9NiY9nY4sFTQ+VvBnaVZ3ainyZBPES70a0
9/reBxx2kK/N7ov9z7vOpTPGxmHWq2UQT9jvyUFWvER2L8Es2G94ZMtcIGRS1PCp0Vh4yjMl6Z2y
jV4o/BEvJMHc5bo1TGBe+5ithl3C0sviTTtUC5hlegmnLzWj5SNvuI0D3DQOg3UemtpUWq7Gh2Em
Ro/Er6446qRMvtlJOnvSGV/JjtXKZilo0D/F4qdlHRd9WgwED/b63ybMe1ytf1XNhfB8JI89gc0x
H64gGMETa/CPP9AnOj02wG4FcMFExx6+nfmVDRtUyC78hBSzSZJMCmKdaZsfvAImAT7IazTN+bbw
r4IXZsiTgNy0UPdD5sEofLd1DZmDHQXYGc+RYM930l8WsYj6OaizNUbvyBmeJqfafh6eVG/imuE1
+udrKggPAOlp92Haau7bLdMtKBEI4WpkSPUmmkoOdB4yJj7g+uYbnCsMWvug0s+ZUwqfqOEx2PGu
VrQY7LxNx+rAYUhvuqca/uY92I1k8HgjDsXsoUd7D0VTWalYgl29/lqJ74F0nbzT/Q6y+rhNRQww
VpR2Us3bYtvxafltUXWiCIsmFZbPQ79Hp/3mPN4ELavxuZlZDgEBIX7VQVIISoqe6PPwvG9TrxPG
kwAraihojX4RPK/2T90v3t/oQwl6B9314uOLfNhZJua4VKPamtzeae4R6C3kWNrRSBo0Pjal5JaN
sYVs2T54jb74wwADxdExfu4LYjOusHNLAZUHdz2skFdr1mG89gQZ1OLgD9HmZR4pCFnhdOKhGX2T
51xMfrQzji8BuvSP0prTa/8G0V3w4sVc7aTLSBmF+BHeEU4hXAGRw/170L+E5+pT+cDO4UgPwqf9
lk3d15Z4n8sQmva95+qrpQ4CUUCOW3EiOo6KqdgOQy/y6odiYlyFqbqgPCgornHdyiL4YBoIv9Oz
ZTQoF8sMmUL67bBR3Oc9uvzgOtWxjIozzMEukLcWiAD46eTB9rmSEcXjeb6Dc7q0BlZ4OusG33Gq
EHT+kkkJa+KjPwZGBf8FiW9qqMlPa3mlUoxIzxpC4PUzYUp1Ky82h7dDpur3M/zzd53IUXJ9c95K
R1VKOQPJyDsYR9tzk+OrN5VSf1hXzkp7LxfW6gxoirM6B6MdqhPjA3p64WL//mvhPVKfWPYJUVZY
uS22bG7Yr1PcXQcEuTat/uKltMVrjhmhmg+xks//7j5AWBxa1NFo6a4HBTa9fEKR3bxUq4q5I7Nd
/FL8Ginyj0ZJ1/EujuDKJI2yXS+NF7N1kQC8lyf/wuTK/0nLH6FRcJd7GFFY8EaQykNVz+9Gau9Y
rFxdkk8olTCLyVv8x4GXXU/9cjufaJ1FM3tJpmTeI9UuIv1Fu00rym0jT5bxOI/jvQyJqz2etIT7
HQHziD9VUKsKKw9midKNf2rKtcRSUPE0UIydRjMuMdBjP2mJFB1Qo9R5LTDiuldnolWIBVr6hQEc
LGAQHpfdgMaPlrlCR5RkTchbJ7XsO8cvbj87t3sATFwhC/nc5tNBwe5UDYDK0WqoMZFGnHL/Zr0o
PXDvup4ljP9cpExuOvk6xM0R/z+/B0GewB7vXzs61bgHSQiznlGLifYWzz1DYPsACnD3qE1A/tVx
Tq+227JFy1G0j0uC8OJd7tDH7urC49J8dy7M3AI0jdFIultkhVOIjyTpJt4FqgxPcc8Mpn1kFr3B
x94zGfA1FsWUpcafmaeu0ib/ZZpm0kYFBe1Wcj8tjLXglHi2fN0UyKQmT2tfllx21nFMve50cdbK
MqFTteBWTGv+3LPllUzCRKEHwvrwYXd7qgAlSwtpflEYUs7vB1IvQ1/tmsA8zzK5r+4VTi+fmVP3
Dpc40JlKRwllc/ZCAqnxV9kVmYOj6NGRC9Qy95FzkcelPO0hmWnSzl9nHcEQxdyZCdFvBmGnPV54
EToZvdZl0fZbv2DzpHRcbYIfxUAAz+9rcvGg57jmS6Q+y1+b+JnBtfo6AsUcysQRVxVwlvImcgRd
Qlj545vZ3n3QO65mSMnITfZceheUXRggOFNmFnRl6wcmahXmCvEEc16BuTbac1tCIJ59wEyj975+
S//4QkfYzI9TgzDn+BsQj/xjfQ4WT0IUy8HUQLhBC0ZNHG9C1qgFJy1qrm0fT2ObeLXP7sWx3y4r
9fGj7ayZXqqoYcEjiyhCeszAcJAiD4e7AZNCvbvNJ5TfACPRXZ5q6PEGBT7hCJxdwk6I9hJWn9hD
GpMCE/OEZkn08mrqhpei3jcHszVJ+DR1kJatLHTbzix3A8knUKaObkZvce6mjeKdQu5ngESvy8A/
QJKaOadhE0DlfMp4d5eng+XDDBoLgxt+dLuPHy8HVXvt940a696ZLp1g8XfcRqSQCnThc1x2IMMj
dXM6uVyJBLVmf5iEmqMYGgQnpXiERE7rXDsPlMJ+oAaW6Jki33ZwjeKiCsF0uhLE6CK7RPbJbqXb
sr0MygAIGUsl/nl2cP62mXrahfQng7hVFFf7j3xjSu/GayBHUO2dwX4FHBSI2G2gsYNWk0oYFE4G
DBzf2KizElvAdVcnYd2GHEisgwsMGXw+uvvLX+uCllQm04VZOtOTNAaTV5Ig1CEDnMS9GOp09Cky
lR9lk8X2Bku4iSTWJ5XABR6EPuhrc9xZk9hNRnwdgAsPVr99969TS9KAjAOCWcrzUm1qlvKEutOQ
Cbh5nsZp2fOKBMdY3DjYPxh46DPgBiSF4ruT8le/Oukl8MZELugptOsr4Z1szTJTno8xhSmZVbDU
fBe/9nC/FSHPtilSSOswKTprnWMcbG8LPDC5ESlXH3ufS8J8ps7nikQRzLWtwWEeWfiPGhZgyZQM
o2lOuf9qegP8yCBWFvNFupWstdEAszzZxYMi4miSxN55a1JdGZp7jsjuAT/ThiclXR0y+grz8H51
nb2CsXphFvfGnQx2okP2xfNKm7qkXC4SfW3nS/4AvXhcDNPXhYFsO5OWFS4+RD+Yp9fJmdN5ksUB
lupubB2M32ZRQ/ec/0OVAiTx9H1wO/6gSrxZGzuz9b2++Lpvt/4CzXLHx7Tz09cGuogHpWycS7c6
dXdELcD4/mW/qb85bIsCdyteGu9BVqcA3rmfDG5A05clZm5kQAekDNxF1XFK7EEkZnQY2hW94gB2
iqAs4qkS3p/B3H3MSFbYPO1X6SU/FT+IPz7yLDYFuXPP2B06kz5dh1kXVCwnQAKs0WMmrYW+pNOv
ScRpPwOU7+qAuBvfF+IsOanYs9sESK9MQRSpaW5+5cWC0lUcBdPKbBXVqiMsGW/w4NKTEDP82Gte
f55EsbsjDJBgF15aFw9xxva8qVojPua7mc5F+N05RARihFWOIZgGO4sYsdKiOMXqJ+MRfaB1zh6T
7CNsI0Y06V9TiV1dWi5FMngsKH9g0f2besiW0cQaeszJQfLg+NZ1DqdlFLe1mdhAZZ9b56ooTx1r
T7cunDXq2pjVPnP/mP67iKEhqvpAQ91KFZFb25w3DhquSBHXELEsposY4ELR6QACS5ZlAT5Dqx10
AhK8WavOhHDl9ewbTKOaRkMpGs8HtSG8M76kIk8ZKYAdnf9SeleP9eihE0nMMJV9u3y0bJReMpsn
W8RyP3YLabi64JxPJav8BWj9lnCNDY8VcgymQ2sEW6j2uyyw7miNJ2vr5+4l9d+rwmEGjQlCitdg
cU0kXkI1mVJaSsO4M13wiSDnowtxQZeaZP4cxYyv5q7Fsrfb+oGvOPCzuMiaNxIcSxfno5rf/SoC
piwKOJEdhG8hbpKixpdDT8VyJRdtXVxzQJRa4khtlf/kmpF2jOwore48+MHnFc2+tU+TyZ9S95Fa
a1U9WwaX+T7vuR+q1kYnBt6FIzE6EX7Jncsii43035NI0YzmsJ0UJKEFfgO0ZbDimRcDxjgSBp7X
RnSSy7M27Yx7UKydRBcP0bKdY7LsKg4EeQLqht7DNY+fO+uK9Gwqn2cjOb2Wes1QNJSrzCvDpFc+
xAnj50AtEY1kHv9VlJndK4e66UvKLjugXOeNbmYEheZPvd/gVrBt5dhG0b5t+R9HBmisLlYpFQNx
8Ycsh2s/ABqCBnyM4O+5E8bsck9Fv42PxpHt4a4r8m15aWyBvRysRvAxBJDlIe5wTg6Ubh+o5leu
LkPLCgU+5/fGNoRAG1/yna+D0LVS9Vr7IsLpb1jwy23BFhFv9qakJ4uD2Xz3lJBCXBDaabw387Yp
kDA993WRtwL5p5BCh4LOb1ducL6ul2SXlZogUulniyIv5X8QxDEY6mxMtFCeqQVltXQZIsHw3v5o
TtJ8c2P7j54wD2S0f5THkrVrYEu/yrUn6Kn3htHPa9bXCDMAUvJ4cWloRppAc6myyDY5A2fOdU7i
xbmPIdNYRsXwkXeoq/x2Re3n9TVqa0kAQKvBMauQUsIb77CGNSZLbQ4zNCANz3na8Yz6RBgP8Ah3
pfTbBNK4khh5uqrk2UBlqmoIs9xeEqQD2Wc1RFw1oq8oC/8cDLJfg/Tcrt3ehW9SLudnL+q+HaNG
2/uc5Q5QVkHjvnZN2v4UpyKbcqXTc0GonWexAl1S7DqvJQ0/KRVQyGitgSLt8BE1j3dqDjhUDta1
NmBW7XtogyWF1yF93dieGLL/rw/5xFruPcyW9IYNZq7qOx0a5KE0FCsMgIHB6cBjPV7CP/TBvqut
/eVW7PR0SZzIWDaAffRWaYTlXQriv07vRP93W63l6DXqgm/I1zkXwq9wwtQ4tuozop1q/OkEcGtQ
OJqfRDDaRqRzx2RbZbHIBQ+vBEayk7HRMLRLutU6fv7KpBkAYOiI10/JEBZDzqsmUWyiwzBBXgzK
rTkHCbFs2gjBI2ZjV6mP/FB7mm5DWFz2z1SsntuvlCy1AVnrx8tMtaIVUd4GNbfm/GBFprjwzkby
zEarCJE62zZedielHKRsV8cpfNP6s/ibdCiFwtDed/x0bmuaAQyndMNu4M/TYCqkVUstnt92L/JM
1m++GEUG1M+wnbrf5zMI0CjXgbd/RGxSQdiowG6Us7eGjP0B0Ky6yyfDe3ffZKRCDZuva5XVfeg/
7AfzGaYzviLSVHYX6ACIlMCTlyhKGPC0Y2qpW2UPtonuDtgWjW9RwxFo9tukKE2A4PQ328ZyjKHC
x8o3dFjLaW5Dq9IC5CRlLFyM+cjLPsP81cuogRtyWr/2DwzWlMKnqf80GRopU+lAOUy3m2ktm0Bu
UBP3Y4pE9gDFpD+WMCxcTVZA6ewAg0Ppf/BlOoIzCWxT5MxtkPtFTKd9amqDdJsmO44ldHMv59GO
UZn2wZomLQpAu001t3gWfXKNiznXDX8qu3HlkrzJYClb9QA51LgzlR8mENN1ECTM5Lxhnp4WvQau
GRyvI7xgyCtwi9XxC2qGzOw2p2InKPEcM3pmipao3jF42WXE18VQ8DPk1qF9SS38x5sKDd3RDrXq
3stRRs+UBAlaF6ppDp6CkDr1Ke5H3MKUtasm/0fcJnhLT1arcjH7eX4L3dLmNdeTGp3ekTF+g4nJ
kX+Q7wmIz+9u9J23qOLMUSWpnTkPNM7rp6cafu1JWLq8YYy0RZSfU/+cwCEeHaWNEMDVDOZ7Hiyu
xiSdGoSMs4YB3c4alBuSGO+MP+rLuissGam0IpVRtZJ5Lofit/DR7zTnt1xM2ont8YjHTWCxLGeP
dDmCOzxTW5IVfCbDiFZj6w/XeKKAOUKOef7kYzalTyn6v9wvk2omVIZkE9FW6s/VVmcjOBaXtSNy
hKUNHz0582jMtCVIAEosX/GIlgDuBPI3OwHcwTxCeZgnvy8+3n4nVhbGpLMSPyfGSp9i7jjAGBrc
4jNqBf8/4TvfhO67aG37bp6j0zNpiBYnJ7orkdk8K7toOle+Fg6r9zHZmQrp+fvZVY5Yt3RGZJRM
sbxomsVEbMqs+rlpdhi0oYH3x0n3wqjisxn5gL4gImDwbTLX4SI9SlGvD81tbK8bx9EMZFttC3ig
V3trWHp10FrFcuOc/+NIID8bDMtoRXaos1dZkLt5WcJ5Y5qPZZy5eQyJjwO76eA28yJtazrUQpSW
Xh9hbG/yu7TIWkdTjWNXWD+tP5U+qswIE6xCqZOG0haocTAivF/dtwcNgngNvmtju1WagGtAWKGa
tdG7fYEbbRfkHrraG+IPhl6+2+tUDlekHjLy0ls2Kr9c8a77nhv2S5J2V9RxACPT1q8XbWPtKeiu
w9QW+HLa+VO0qAcmpZYBQFVPHrf3Dbx+OQ2Ot2NtasUrwj2eGsOBiVJ5dYFQA0xUPccN4ycw73RQ
GlHnHgwTJWt2L61HoI2RRh4mowIlfyswsTqdlGV6qAdb1E34qF1AVixgCV8CbjvObrsJiMwtmLEi
jd55K1WNpt/LkuepukK+IO5yFZrYrTbZcanwO5sstSKt7Xr0xG3PXc3MRL8GGoBWFSgktLiEtKNp
P5hv/PMiwDApjLFZ/l/ZbqBPcNqubArEyrMdMAlAZbgjrdX/sNF3YGsWUNlN8VAXoT7tTxaUSVtu
rHY2aUTH7fpLAtdKzRVVQ1y0zsyIeSlTstUdsSuG9z7lvTjmqOwL+eQJNCtseRuhIM1/UJjNwc3/
FMUyfj4WrcyFuvFNjfuqpyNjcT1e2qHpk77XrE84YFhRcPSTGFO2fS1YQ9LoSorwiUf9hO+l5OZJ
D+Xb6jlDLT5fkH/0KxTMdhdo06jWVHMZqfVLrKIdxCawBpCvqR0XUXbhqxeK5uSOXRqcVnQqyxKx
GlCatLNZmH+OiJpGkw/paSCypEDGCLetFG3fOotK26r/sTn7lx/a6j9sFZ5pkvzN2WOOSl39dOys
HOrDq8Lkcqwoj5LL8bubTuFWQBKvzViha/GuE9cU0zL0/kLOeHKGGqLYKRsApMqeqx0F83JazjLy
o2NPk4sfc2YK9v5picmL4BY4yxt0xnz0aSMj04qnsfDxd3NMToU/hCmwX96uXvAHIC6NBHuT7zI8
BkSw1mJEzmbN8h+H30PgHevItlu+4KvLCRq6YpbOrzXFWBfOJP2db6sdvtlpGKchXKCueQc1F2dL
4nsJlFjkV+hjeaPMw4F3RpTcn5eqYfgKtLJddZ1zAbHlttr+SMGOceJ9mlt8eQdBywJnfckcCNgh
9U81msTUBDCyo3piS65BnhUNwr//geXf9lj/4Tu+eV7egnggPD11b1mZ0jex3FiIsZcIrRIcwbR3
R5MpvDG96GiaJxTS+UAq+d/WgRjp5cRVXh22cA7Sl1UD15BzhrY4+A4nTetqLRvagEOw+lrrGW26
OSF/81E5y9fWjAeHlpxKB8cwm/qbhKlGHPGWqKcCCyKWtEtKEmqFaEKioTkSAJH+kk3GfJyHr7OY
1BJ66fH6uq3SLQ3zTqx2SbbLyKEFrBDvA/Vs6MjZsMpuKuKbAW+PVsMlm71QsBLovvnF+H4nprbM
jWNDA2J5Se0h7OkuaXsMi6D/Vmq6iRJuaMHKm0g2C0FMcXBJEP7pir0i45HPlQf5mO3PnqeSXNaG
R4/DZZ/ggrM+fWr2OqlHF3cc6sfbzeCqCqurueaWp7dWzQpSTP7A65DSapNUiIrJ/DEkyUvYjHTv
T4Hmyv5BARXBu0Mfe/ivcm4Muq+5vA5O8sfGXIxiwIsugnQCoveKYFNvY8VUDg/BecmWHALbbm1t
PspBHrnK6yqdOVWAq3zkKZDA+qXbp104B7jcno0cq22oZbdhGY9jaG9kO/R6qzPgMTDre5TZnGpw
bSWLKASFuiEqVvcegAAnt5BdnNO0oB4lIY942WT4tvEkZfkA8UhpFMWHZ8uLSs1nW4//ysL73J39
DooqCKY5xeATc8n2AdlyaDzJ/VUV5mNMppyAcFLCHUmrl1LXkFu8EB8UibVtomd/JrKlvYTvp3qh
nlWNv49jkTCEWLl3blVxl2p5qrRQAiSHH90zRcntcjV7ovOhu4HxSpqK8n93dPPY2hYB0EzEc8GW
9C+O5ERO9MRUEoG02Tj4bfQfrn2jkyUuGyAa0MUdyXE++8fbNrVZanjdHkgFP9v+WfqcnSZY5Jha
TBnpHo//qKBNjcW90Vw90ZmxrRP3w5QEVtGgswBXd3UphUBV7b8MRlYT/R9eJzZTLwMYU3WVEPYA
0FSakxSCBb15R4LBdWITf7jrE+qVlr76TVOLE+vppSaRhOsNR+fdOQEDk+wf+BwjcQC5xkhb+zWQ
T/TKSMp2FmRF5G5DtJMeAVpvIPYphLZyd3uZ/Qz0ZObhwybUzUOa4a/zdVbRbF1TrWSC6aLPR++O
3fCy4iUrzuo/4YOqZxv7oL4BisfOd0+lRwH7WmNKdqMkZvqn4dGBANqJ8fVZgyw0EEuS+0dn1L+o
Txdk6gQFDNsdg/xTVnk+wHD4eK5K6XN2wlxNt8jWx+ZGrn51Sy4/9NCTztO46Aldf8kkfX/0Ch5n
ACkvdkUber+aGyGzBhG+reDsCL478PMtcvCr9Z5SJI8IoR0g7WvJ/ejzikNjNsYTCpQC5P+cWi3F
Ly8XClKGrUfeIXF1UL252zaysZBz0QVDrYAgqCBO2G6SDqTEA+Tig1iI2XzOTKJC+bfTakigQBZY
nFtWb0YyHYvNlcGuE0WYYLEvhX7tlH7Pssok75tN76yg8dhUyZpOKt2bSRTDzbSFY6V24zqLLHZo
f3lPv8bKfOeaSZ5yYROigneHZG+ndqjXUyN0xi2V0Hi6hT9BUubMTL8mUXsE/SYp6pOlCTVFmbTf
QAJtd6JnoOyuNPD9mBfDJaX9qqX7s9s+mfmOjgopFCF6SIO8qYc9ybepONFjEVsCp2biUO5MEbu5
VcoDIx5FlMKkQhoOJmJ6hxcus5F5iZRbpxh6P7Wkk/BkICYEUYtggm3WzzAs0gr0IIh7SxPoP8SC
HQEQdfOSFHxU01fhGzAE/pwiGHVSZ3kZfxJhXt0bAfkdz4Aag15fY0pbGqQr+6fF/XOB7y6t7MPB
fKGIgEq287zfF6wM+gsjMi8IuSgjpls9oOiHy9g8XHnoFhNrUykvNqv4oM6djGvex1PDIlLHoPMY
nu599E8+IhncU+zxMkG6p8JdV7qODz/qYhzlgr53i0Dcfk+W5CTymAHpRpm+KVfWo0glbdxwd6U2
eur/dmPQHXq1JK9TM8WFrWIffBYyHOfntjSrDH4EkgY7emUkZPs9v+AiZehJZ0Kps4vAnrm2A7Uj
9P5juVLkg/VJDyPFN4nKJ3129GQDjxbNfgAI43svjg3sVGH5nO+4Y/AGGLO9kT4N9ZQo+yc+2Jfn
4/P919XUGK7A8TG/NqxMi/oecEPupyRrIIwhQpH3XMCfo7GjmQbxlX+mMvAGcLEH5lBqmguw2IVT
9PVEIATc9NHQ0p0GRPBS65xTopOrX8ivTQ1hO+rOEjvsEMVRiJnR8krFhcZCPtqXUPlipmJK7x9r
S7iqxywtYkQRXQV4ZvzgAOClZNeDRefWCMoL9KDjMH0nxBV7GF6iYOZq3afro/hUA3TmGCIYpj93
PoWL5lDI5gYxYAk1H5QomYxQvU6ae4u8MJweiHp4r+UfOtCCDeVNWW6QhDU+Kl9eQna+PES50072
MUoP7ORHu5ccopiyQugxFhCenOK4STwbG3AQCL+xNpRP5F7Ev1xFRtJsMCLWY8Gt2cJvIyX0gwR1
F+pPDx7t3tzocRFcUwtGw65jHBGRWmvX1kcOuA7lTsHR6tI03G9k3ri+cT+Nv+7F+zOCfScxiMbr
0ZwEKzPhnHD4aJvF6QwBK9Ru7qp8h/b9NryIymLaZI44DlLY+marFVuAmYtSwvzsDv2cN5KO+2e8
73Xm/pCebcmTkEelKYXIfLLouVeaMCcZ+cub/UF/2BtbF+l0jc9ri26Fx697XvGePtGDNr4m0t3M
tOxCh/oVnfw2RmvfvCVVoqY3PJLxXrLWW27PtC2P6Zb54amI8j3ml9VhPYl8mLqnrEtp0/vgj8cM
vh8Od5qS96UWxNxsiNHV4yZSZI0X6Q5B0+yOR2yCC860cJyWVYO/IXI58Gdr0r8s+LaSJwoYNxVr
EspDQllIZcsl63Ci1ZyfTdILkqq2BaeR3v5Zgj6MDrfXn3TqdjGE9bsHFbnlwvSRiBJLjSKFSghK
wgSif34pAqwyaiBUIKys4GYzgeABzB402KDZcgD/Jt1Q12FziLxw43ZEA+mvdddkINMttPEgA1KK
mc1OAHFvWaOx73Nl0+GoVC0OhqebP7iHi2FZIo9duaQHOgg7pEo7BRQGOl1CFbVXVPGLiVSHugkv
LBhog8VPp2rka9/9bErjkkyKL9lXUz8Fcdf1+bbt5oa7235b558AB0liM3XTFjP+Qp9bi73thcic
oSFbRNdxh+jLs8LhtinG1EI0M/ilfePbJcyWRvI88bCLb6MC2UTM75rKdMUG2LpHI3V7tW15CX0t
dzYCAXmXMk/fTqecvgLVkgs0dahOBEADtn+kXqNizVme9J7l2Ro/kx4sfXVhiMHo/wXrzeAn1rKq
n4Pm55eEQx/wcaI/ekm58DZWDEfcBIh9fCupFRziJXsiC1Pubw5WvWU3DnTGhjb1AFgG/Q+BaYZo
XPkQq0sAAbkSFMzcRdzqzSJsGFvwJ6UG/P5kjgUD2uyleypzMMefg7qXQ2urvevhQg0U9IdTYMUp
1IccKHc3pysHdVBlhYbZEdqQYInNzQzd08wz8q7nYKiwITyHBDw8+Mrs5nmBSyfbd2qgvoc2HV5D
+ot5cB6FxZGDwMRyDSCNi4U/zgf44wM7GlqLlg3BUXUB7sYTjyM3BkMqSchMrhUARAuV0dNwyjcv
TcxfjbB/5w5OZG2xmw3VkRHzfj4K4Y/+2mFjnMWqEYJ3y4rG3Fdb3mNcS6eHu1M50cu7thLqZMq1
HbzWEVF566m5+t+pNNytvR9L6wFFS954uaSJF2XSzBLwlLzh9zrmyoyt3qcjVwuO8vEENeUo8CW8
nu4EfssEkKGA42aGwJuus5ffCBycKer/W3jH31kMSwiRDEH64QuqAtkNsylh//MJzxDNy4EfproN
Zsyrz2Tlm9BFX2hlSyqGnNQA5c2qRnmU8O9Cjx/xhNlgwcUreow9huCAiCXcXQpg2S4vvdobLVGM
hoaQLSN9ge7N66E3AicV9L9VCqyuaDagu/W55g/w/l0o2I+fWOnMXs3FGEjT0BarUuSiCPdL1RRc
b8yEvPsCUzAjyOmyGrlbO0m/D2RdIz2+sfbDdfY2vXgb/GY6f84+Q95YEn0b6EkSG7FmyXiI3YV/
eRIyqlpdhEPbNt5/sexjPqnHQWnLonFH+bEwQq1isW8Q8Cx9waW4A26MkNE+opFgqjvUN3RmKsnR
2Uv7S4KBpNjYppzSiqQXyS/RTERt4ylHiztcvqmxIXeasxxGYr3vWddrdaKgn7/AgwoED/CJMvOj
9jJj9CeO5dlyIJtrcK+wGJYcd6MroIRic/YIxzPNmfDdaBCuPOPdBtlCkk8b1a0okCIC0qlFxC0N
XiiU7qqpriDhj6nkTLpZV/TDk4bs18Dra7P1rgEbFUyE6ZuoAV8M7JpKztuTWFmUQWvNnBR6Ht+z
/nupKR5xen/QIhpo7145JsedUHB33xIG4D0ZCC3ZMzPcMkWeuX3jOcIBkYFDAcOAhnEOQ4PsNiQB
10VDGnW0CBgVQGr506xMiWWrzxN/Q1w9FX3pPsxUZc1tcM5LTtMesk4YzDFYoB+8oxxWGjVTsu+t
W0gZvgsjsHcnvDIBcTsY5aTeL5qnIct+NDta8MIfCQJW9FuezLZ2W5Z3FautBux4dGBevxEdPfQg
WmI6vQqW4XFUbQBMLwAaCPElHjk//MAMsukWsowMDgwXFVuxucYQ4cAHWf5AanhmKdZEz/LCHuun
/pEUt9iOS/7HGNItE646THgdUsHtra67RX9xrzt8hsDQIxkPRf8hHLhwnXNeC7AL0QWoFLL7kKqe
P0EmAaouAE3/arANycFzdtL2WaaocIVdKLSnFcesBekxDnlIXrERd1zWKkT4gF72eqfCXWudT6rG
mTuYEmtRzcz3WHXqbflyVvnCRAc85U7gIP18icGyTQ1vJ2EPkY5enmDtTN6wcg0z9KPpOpr1KVte
6KYDyqY8VMJ9DISOOlJsnkGPx9fkm2kX3bOjLVia6ik8xp009zRnLSSFCaovW95T2UxFGCZphQqg
6fIV1Hf1f1Kuu4W1HzHXr8GBCpRa1aG6MhjOLsgAFWipZXk8vtq6THmgg7rBAFcfNfcqMSz0NDkG
42tvSbisQeKvl1cBWKJrUZiZRDvzpBZgWbLqkMb884OlfMT28doXbKOncP3L1Ic9BL7hAzHvw0Ui
MH0jFZnH4vnlOirat/d2a1EFpOW1p1S3ltCQ0DlYyAj0VABNLVYgDpcFrk7cMq/sE6SrMX0lk8wD
kDIGE5kJyyHna0kAJ2YOjL+EnWmMSfZ/PvVXT8wb+j4gEglWCmz2ZWhoU9zEi0lNyNIJAsk/XHjA
yIiZy4/6ASGG0A5njaTr+j1TK1P7HC7zHZz02NoC8R650yxScFtRtvIRcBVY5tMtf3gabTnKWftP
MeGES5mdaQNCaoe6hVd65ts6WDd+fTFr15ptUu/mlA729VyJpIa1GgOH/m+A9VsL1vDn63AyuWOK
QaBCgaZpy50l95ti+QVMlzMyaPu8rZCjJIY9ifqYwgWuxanojA0S6VKszahwbkR7BNt//2b+Uyx0
zhtN67Q360gkZ8t6TeDjTA6oNSCv74gd+5K/WrT9nfC6ATI4NEsOjgl/QGEfrZvSzdX62OV5orPQ
LzESZFKJttabAJ7zAG1K2A50kLbndE4b9hIZZX8rUMNf+y+j8sGl8rGHkeWPhAQhKSgpYVRrrZFO
+qxwo2nnW32k5C+qgIzooiXcXxi1l1bMPOWrBEkSfru2rV4tOfSmQlbdFprpILwGqjC0ErUgV4aR
RU+TxMfTfI4a4Kl1Ipucmjjk0ge+BdAgnThtf97DHJ6l8ERp5AgrQeTREvTevv33w3X85O5tkZAl
1HljQfWEKqbnlXePkk25eSbbk3mLY8+my4SNQEDqJNdbhELJ6hvYnGGt03Mj2eP58YumqsgZt2Pe
/MFj/jy9yWIYHUjbPprebD+7ihM+HOtpyS+JECVyM8awITXXcZsX1XhUC+spL08bWl5XfpPuS8L4
3IGx3tcBa14XtgVutCIFfiZSsx//7YzwGw5Q3I7yBUulkFgF2xwMyEEQEzs6E8e4Bq9EypVvUT/m
8zTtpyXFQCKEObjbjsDVcg0dn4b9XOYHY6P5Jr7ME1wCe70j4/DHxDPLGdCXeLmAQkLkHa1iReLa
SAuTsN8jthXcv75ZPFmYYI4doDecNlRecbjlEHUM1fiZ1X8bNJ1NLvT4aFxXRrqvqDJtJFZ0KjZ4
c38AW9WKyaJVtgBex1gbluWKQ/X2iFiLrgHm8frw1aX9yD4RI//v88yLvOGxVGtNhLWjJhptVECL
ygA2e6dOXXBji7GaOqfY0vtnfGJvtsWG1gbWY2B/cCRNnuZIgmtQQ7HHCo8BAXQf0HRtdFNvhBvI
k2yShNEUrJloNyFKJOfpnslvj9RGfFolt/bRjfG96b8BQvNN4Kwu1r/QWVsM/DqRySvfaU32FP/G
PjLcafz5YY0rxYOMqIFkZeB7OqE4B10KPLnSXFKqR8bYo9ZsF8S+KsfLn0hwni8OpbjCiFZywlsK
Q/FZ5M01h12EgW21mWk1lsullxLRolu+eJMePtUl/MO8grOxEGY5Lh30jLg9C51lXQJKhnQOgueU
KhP3Tfzc7hEwMQhvd2wTvepXfkzlcvxM+mQcckdgHoa8psuVZjxHrk+C4KXuI0SdYspRSQfhuMHN
yd2m1IVC8vkVBnD7CLAkESIQkX6q+dIcz9SkiDAe53uWSmyKCbJeIMaMYh/1bZCfVjNXoP8y75PQ
2pniF4zFYjna/3UtXwCrkUoVeHfyDzR3fYHNpaQkLS+0AwGCyPIIo8v/a/46VMimWQEZelZ5kQOx
CigYKThVwYRpxK5oCHeAPcqGzvJ2XhO11hbNt7gCKmVDTgrToyMloHs7dnffWKXzGJW+7pnPlLMQ
XNiZNSC9IFAbo+D3xnBAk5WGv66XJ6qsY6mIYaQUlSG6zaJ+ZV4Ye9kOCCCVkR8pccwvl46wLh4k
HlBpfG90BnhXtvHdnN4bQM8lOjSpYCrh4PuAR3QMS8e7kxfB/pHmXHsiVda2NHLEJuatKfE7AgyN
3zKhhjhV9kPIF+1vt7USvCPwxJp6iMMw/Zs6eVECdnwgsRGfwKCTIuAuvyvMO950LSGHcVjIELj8
YQ2EEe+TQlaPhv8lUpyDF2j6yrFFvdiL2uE50ghf37Ftu3xzyjsA3DpuXZDXlk2SekPDEaLk/dbH
/TkTldk4Xzi9YTn3/ov7aStpO14mjYGItHNwJPPDxWGR9YBNic2lQWlQyMgqOdYCnaCRantop/1q
4YrDtz9CUy8Jhc0gyfXrJ8Mtk+IW5jrhCK/EBGPfb3zOP0KqAKkHCs4cCAERzoP3i3J9CNZay7B9
apg8OwEY2xhfl/r7n7bKCpjTb2woX2wknfEz+cvtTSHrCOgxgxJ4Qm2E7hMmv6bBSgAV2khCMY5k
jLoT9bHfnmAS7YxXSvTBkMgfmcK3If2Y7ZsbpP47642TRB79uSynSB1ToBWy6K5nY0pQTfuIVrM9
eyaAxLq0nEpTW4nqyjJRG1KD+ZfjkJT/W8XHBFQKcAegsJgh3gyvMKDdF7dGVpxjTVKHQcQV2qv0
8N7yG94lUDWrl8daEIOMd9k0G/jh+GObDeH5e0Sx0aQ9gR8w6Hut6rmM4zV0xM+vxS+4Y/ZPBBTB
owEEOQWTzPcc1PLMhWC717F8TfnirZG1ExE45GVDyNC2PuIml47H3dITm9NDoqoXnCX23ZtWF93Z
qB8thqDDfZVD04ZfofRBkMAtfdH/LsxTsnwdAEMz86L+tqshDAxLS2lgBQUWbmBICE56OCGUAv4A
bsadI4PAUt6GZnQAm0T1JFAtl6NqMaa02WtEsPqgPUqjAeZCTPykE81q7feOzvBTnAU1m45t1oms
dZkUVAF6vQqNJxKEJK3x2/6wyLwUTmPGExzreSd8Mwrd0+YhQgvGap1clDRxMPjeaybkj8Q3eS1f
E2mA8mVpgxJwTfKUE9tQ9PpYP6vBaFGla4et/QZy8emPzm8g6AmyNyTaP40CZAHgH7XhAk1UZkJa
L/l/ePTrp0kaRqzAcijlCmKj0qxbhclTXIeUzroPVjF0ojbsDVPWC11iBzJxTXEiDJ6akMLgytZx
7RHsAUaYfFEaBMEBn8Jy2nmXY0ZmO2IGRRfhXCxfJuWhNrJ10EbCBQRNW1xA56hxLrM6HiJZjuf1
DTv2jca3A0za/jsKwu8XvtyFtD+jsD0yaTiiMEt2Z0zdHWUdtc4843p+iBRWpyV5T41T5M7v0lSk
5hQyHd8QVKuGvhJaxH49bICQ2BoVimGeWEC9ZeYlsPc/6Cz5ztGuLHYI8VYcTUZuZGIlBLBCnTGu
1V7MA+TYrKsTBG/w3mJLHc38KcbRYXvXqflugoSxGUsgk6vY6+mFDzWOCfWgPh/zpmNkvxjhJgSv
6/kQYo88TRkZCsn86vNWhTMm0s9Kq6BxGr2JHfVgtjcrNUM26uJuSwlzRu4ofnmmia0JJmbgOgRO
dt1bgEF+EXPNdeyOw9OtJbB8uTnODvVSB4kmp5VBt61TSDvvNODuAZZWG95oJ6nhsVpW2ommQ2A6
gZzRaXmFZYoJ6bNonuqq90+5fVBH1gGUxd5O++JDMRaz/y54oNE8etjI5n8IO1dlr9QyOdtaWiQ0
uF1NabOHaRyFHH3WDfJGW5lrLyMcoE11VxYM17RUEt4TR7PnY2pKvyRp/Jnqc93r4BnO7lR6Ofpv
225MBGt2Yw4oxwnoHROty8q2wA8pFdC0IcyWE5x0OhY2WIi3JcXDXmrUfXllBmut4vOSqi5c429O
S5/m7tzDuy5mRoRM4iQjm5SVdt1BFlBn9s1bl6vRQg1HI2tyfKFuT/4czJnduTZX/zLi7GXv/cnr
XSglPerSHEi+y9LLLTuGm26ElSz6l4/WWHgerDXT22y6piTcHYRXjM80pfd61w/l/ZXfBoyC5BoZ
zKUu8K58KQOnZ/e8AsVKKNX+Q2CkbB5hp0uYq3URpTHnlYoCBKJs8CJMwv3suxQo5yEXQS6V0UYn
JLzTefmkXqRSPAseuBSHjoiDMl8mFu6jEnL4IGZkdKJHVF4za26/f3LwpsWqmtlfekht8eFphZel
zM22Qc35NKUMJY4QaaUsTKDQdCIiQtkXutDqSV+Ov9dsHfKcJRDmUPk0zzG6ktqIEbSxc2jPCkvg
yeIB8zkH2rxJbYyOMvD+EgF2km0rhLWs9MfY6H6ao4to69EbNGPrHUJEdDfSYlGYfwzc2XJ4RZhu
5JlIp9RjFK5EDYX/mIbdArkKayZ3LXySFNidIoH35v2qEzPW2C+HCRLfWlWORYVB+TS0SraeLiiK
DNE1sZmfLwOaHWKFtnuQrp9OQtAJhMsOQI8U1PXHvd2WEkZdTxw2bvhvTl5lZwrMIoaiS4wGzbVs
H4JTR3EEpm3W/8btnEfzaPF6rTBj8FHcDYsi1M6GtJDqUCZ1kk1dj8uBL69Tag400kQHovb1hnRT
G91OLzrlVpPqM8fHyU2dCFhyHW+h4STKZwvcdxwfmvqzbsyDc5WeJEK98lvcBs92tEVtHJSR3JVD
6dy/MxpZVuoZC6QxrUTHBcy91Et/ncEW18OVZzwl+fUiuzuHtdO62GjM45i/p4qQ7dWdgK8XXbw7
d3OiK/DFM5/KsevrtGqBV78yPBeN4MQ9+nkIMHDP+5qFqK5ClrUVnUUNe9a2gRLrbh/Ta92EBB9H
s3+RY6Zu1d29Z7+bAQa2B71+PQjaYlDwuwhX0qyNUTBku81pdO3BP/IZyM2raes8HB3HJ7bI39sn
mSAuJV6Xhatzgm7i1ZbrJE/Ny7D5t0nfQMRujVqT+l/Lr0BKCB2gwC/MWcSLqOhaDhZ+F7tHqyqR
pBzn7lMGHpLkO92rTGNCSrDQIFjWoNHZG1AHGa/h/0a1XY3RPtFRI497sKD2t+SUHTMh/m9DDdDd
n745vwq33UeA8HaAJB+1OHlbZ1iN4X3enOMQCoVdp4Y4gYFIOhMUP3Q2wBBHkzADIg0sJT00DBfi
J8HNZzbkK10fWn2RJRZUApEwjW9MvyCqzMBCI1AFtSRG2K6n4QVfbimHYQwtD6miBQtz9N8l822X
CuxhQ93ESQ6RsfM/vA4TG0YKemwDn6XuDjd3Mr7tsNFDjbEGdcflKNwUx6mL9LmBgl8SN6yLEm28
7Vyin2iBgREINVW2ZM6xL8aHf1PbLKTl1wQ+m3adAcjv3wS9b4jx6uj37zC8TMaWsJTF6JDRnyJb
gXfrOdSCO2CvgMX9o0vtYVVX9rGWt9weEQrEZgkGNWpYfDLZkJ9xlFaL64z5mODyEA5LmZ5Y66r6
O60Hiac1awncz4+YTE71VZ5hnBgmEksCVu5LU6aHH5M3v6KY5Ta0t+GgKW7dI/2LEnw/yqBg6z2b
UE+NPplPgiAcAKt4u97oxtnsoilLLan138fywanFyPiSTFKV9+cJ9BJfMUMk1xh/pnCwwd4vXK0x
Qyh7+wGr++VCtChapDaOcrn02zQjTUT2L6yRj/FtNygg6N1Tuxj7PmUsCuG0Cko0Ue5bHxba7pt9
CTpCz46B64jbAFWmylHb5Awo7//gCH9UpHIVkWeRA6MegnEClTu6GAWFfKwWBPXz/6Xt5hJZtSDx
fH37ZaRVsiSlvBdMSapUPyAPEGX0cEdLeL5EEiNGMOJdSTPKrk5rDitMCD0K4tT72/luaTy/WFXS
jUPgmouq5iLRcbt79u6b2vDgyfW92xPcDql8ncMHIZlt6s2fIOv6Hy5qxZ78dBYmxxcJ5Z6+r/t6
CjgVnrFYwCmG7EEaH6NYGxvRzOuGtisHQ26x5y8+3UoHnv37x9XuNXMlIQYr/ph4HKD6GzmuKodG
4n0H8yk2bCZu2M6kj/8EMRmhOHk1A8NsSpOWlbzFhx6+cn20a8pGPgouBWy5DdrAVbdm9WLKkh4o
YiXu2P5barj+kdqbrg56imUAucl1Q15WfEjQ8qKYGCOfEWS9d4Er+a9rQdO9WtAoa2uTJalCb/DR
7UOd+jX2vOjWUkBaS3u3b8srbCfA3vDtf4oX2JoBUimw9MLGeVm5naL3Y2QuhpXiUzryKwZuNx2+
yXAbWXmycMgTPLRo9n3qXwwHoIoG3dVLL7pKCYBd+Mp8u4qTQkdDZp/RSPpmZFPe7kidANxtYpQ8
j0O/5PgKnjTbQ9QnUb63A2HVgz53Q+hYpAm4c5znxJ39xjBeLWcCaiV4yspWfWi2M2ytMti8B1Hi
Z+C4cyI/+c0N9fBgmh0RLr3CRPEsfTJcqfkqC2XgFpyGBOxuPgTmE841/GeC919nNYp0MwvgFz+i
bSpuHzQtWHnR7RwgxLVEEUL98pCVgk2ITWxUbmKtQZ7oi42MvkH6Au+wLg16CKGDDvA63IRq6nYT
WSCgCdc697N3mQ7+AbQop7eP5df5OTQmZr1Ibo2T8NA0JLKYDLqykcNC+kCs0QgX2mPoANzEmyuY
ulDUmUiCgj98YUvVkQCw4JEwdpL3V3ST4udtK0ytG+ERyJypDtVhdvCiPv9we6AOhhgPPZNM8EmF
c9OSd1JeIa6T4ubAbqH3TiAiY6nz0Bz8NYbQZmqhkt8YzHloJ408QK2Yfpi5LCzNv36N8Cl/ooWQ
/syAbnUGyB8KQRkFFWynMC8FlyPxf26HYqvVwE9Toh2cp3GiEOY4iTkmg3lsSox6QculYfVmQbiI
aG9EEtCA+gK6EHO83nFLtIkBj5h4O1xi9p9SmLrqaFVGD9NEnB+d2GNSp17HG9L8RIdfTN8k/8ZL
rMC5jD2JAcGrK6JDDQWkgcbXASLDndAXHnkxtlNawr0lexfagc6OtULySwjBGOe4epzg4EPTQm6x
gYZFfz8ydDADVMpAKES0ISSaYd8YMyjz3xhpmegUjPg9KZhjcZHyRZE5HEvO4vhO/BTJG/rk1AGE
xeeit0A125AdeUHz9gdlkuG0j0zdjjqLnYMtYqMiAeYY/G2XzCDjuZzTy7cEbHZNpdy5/W9UW8LE
4fBfeUzihkFJTwycjUEC8f1WYm41Z4cIOBA0ySAtU62Rqf4IXtO0eHPzJvGP2YTO81k6cADE2d1w
EUHI4c4vdxOGHF5X+pRFhI3n8C34dneQ11eYalMetEcOrFk9hAGbB5ULjdnT0eFlY9yYlaLbLOdf
WwcnV5RI6AdzvPHHjyvY9N2aPhbykWenBHMenl8nZifkcjFq/42vpHSm7Im0+Md/xYZeMREEZvRR
ssegUpo+6c+OOh0HOTLiLjEIrFGNwuimn7IuZRZTC7uzGdCp7+iqb8yp+cwv3hIhnK1QGbMX5x5a
2TJMl78+ulWH9rB+E2Uq/svQIa3J2Y1y7tU6ypulviPfB03RmeAOeHZZMAPYqNT/Ac7zqfkTG2WN
61R0tk6+7+58fhLCvDjDvDgk1neS4jwRFefECR2v0f1qCuq0RrL9jtASFdtznn8jiOy1XFLttQTT
do5oREfdVphe+ZDuUDf/IWPmUaACFUk3uUr1/bpRplBxOdT6R+pagqsi2ScxdZg0loP1EZlp9IgG
2lEcP3wKouWabGQ6IAaQJRw9o6kbmjmKIYduJ3W0MC8qN6oItZ2yc7W8H2f9r3ZdViWtUcaUfiW4
G/bn9KKJtaJddMECWPQ9u/6662+uK8MPU6FRbzJAYf/UW34+kylr/jqqsI+pS/zGKA6Wgio9MPS1
MR4cr2anIfrSCZUAMnu3hbN9/unghnm/u9AeGalnfGEZNhnNNsJOxNvswoi99xNl1XjLMnRsIWk3
w8BzHG4inh5691W36juh+y9IECSEwK3KuomQKfJ44hm6vCZaWXmy6KyNvA/gki1NcLCm3B5WV8Y2
yXaEOuuVG8z3qzpcIiE8qqlCdLqfdLHy6VBFNMCw9rO9B9bSEwSBtn0qkimHa03ghgEgdvpk8NYW
g+t272w8W1Wagg9PbS5bHNu4xVb/nfONLXptdYuhk+8p+tf4CIrZ/uPu4EKNx3K6apquHMCAee80
y+iovg3FdSDRXgp/jAm+9AhQDsvyETEq4cJqkAPff2FdS3KGHwJgDsodEgHKZHupZPvYLrFvHZAZ
Z2dz6MOM2OnfSVqHxwMMJOxrmn6+L4+C48R1IUMmyeTlSIM05koU1HQtv0K9XScELKXFiXqMP0Qy
1jdloFt6pkYdt2tNnEzr0vLP+W0aWlAf6e5oNlMelZcUIYpHzVz7DGanwXUBW7NV9D10297AcMeT
T8PT7VR2McOVDTegeh/dCbFMQ+2uowKS1Y4gdlvNFbRqx7I+sagy31UwF6Kmhj4TQ1oLmz16bM1Y
hVJbQYJ1mdB3GX/KEROEm9chflF6j7R7zm0uE+LkJwpsNCkSM8r+rOeHmjQzMWUGGr1zwvxRZjcr
6LHTSt5GkP+rWauAy68DHoa+FRbM7c0VEqz/cNa2GerYJ2gKYCWF0znVr8xvDocmIFEXBVkfFKly
k/2a7X+xzvkjMqkIn1zIz7sw8NizdqdRm5qEizzpcEYrNumfkmhgryhuz/i14Pi12qzoSuVXCP0Y
E7kqY+7TXnGsYJg3Xcoy1zYhBWWThyYXEYtV8uVIR2g/V/ClM1LeX2LfrTlv+o71PexZ0ngY8wVf
XZgr2T+7+SMRVJaL6FZAybREmghusDFJMWaIrbE5g9PBQfrJCczMjGJox5PoQyUDwxHbyT1edhFE
a5bWLdf0fUSbDJk38vzP/0piXxg41MPoJSw1UJBP9CQweeTDVase6bdgqSpCdgFTTTWFYiU4UyGf
d6olG6Pr5y33p5EyXNVhBRlQzfCbjVrKU3csBRlYc/u2QPqAEMFX/f/UgFHUgenZaVeUNh5xAZPc
6uDRp1CgAw+T/8yL5VPyrhvV/1lTC/CBTlfoJANNu/urEZd5STED/YNIa+H+M9J9G2+tynUq79nG
q92PtxEPomHmQUdpyO09twVI9hbXdcYPyPbdGe8XftHaJi8dlQIXybeK30O512ZYFAHgTR/PQv4d
1dBFvlEqn3+Q1PAYfVc3xVVuueT7/aiWTB2OKkaiN1w+/jKuncIhT0jYbSUtDye05ib0amX6nHkb
qOz31e5mtR1m14M2zyfcQ/jNzjTeRWJ8lhiw5BEY3cXyjq8L4+7yzOrcnlxV/y+EgjCfYzPP2HjH
5RLhTPBqDwjDX3tIemBcImMP9PLlUaSV32+9KChyjT4z4WyZEEauXzLvx7pN508KVfBUOBOhkSbH
4V1MM/ZPtbdZJcCANjEGxzNItlZ2C1am0hI+i5i0FV6vsnaMtsbwWiqGutIsyrbuuMPfZgM0DL7z
1bDDUWcy1R2olS/bjtUkbTpWMu1QjHzVdMAszEivcgy1f/Q9XkxnjxV7RN7GpXBTwnIGfjzIyxE3
jQdsBv3xlwmIZ+0I81dyUSytPyZaNz7Z3NuwZ2fH1P8A0/43pemDt/qJLsdnCQCOy1XcZvvlAy7B
pveSCg27235GyJ88tcFEGkMUAhdLXuR4LxZxh2pHfU0VMF2c2oF1PMHx1/LulLFh4mXxpHembMl+
Oh5dMR675dRgZgx1jLweWRC092zUtiiFCni1Zw+gtk8wGSx0XQIDuMwzybm77HCR5i2lifYZvLEg
SLpVuRbBDpH+VBjEYJm9zjGUpmM3YdBCHEx7vH/kBLNrhJYIG9Sy26peKz4TVD3pdAh9Zj/22iFT
CXXoP6kqxhRC8aWBlSn2t3QYRr/7M4fLVGzvpte38qpUmb0t375s1qW2QnXH16m8WzAmaE2eJ4I3
4IpF9jaaOyGOx+3qfxtFceF/sIHL/lX6H1fjr/zmUm6Uz/ie2CMlDi2bpUgVo5RSTgcxSJtye9tN
+VOnpl/ptkZ6q87EpgBRLtbjIvPH5uepkUK46H8nWdl7gX7Xt8rKaynWCgpAMrQA+7WrQ2lo0/Fm
2rqjDMoXjiArySfr60am2owVhYbiGCpIDIBKrBQO09R2trvMRsvQOwi3xnYynNnBAjjeKWa+CvUQ
SPSg/z3y16eqCUi8RVcM+7a3cO2dbsMvN5t8tfj6XXg6SaUq6hE9xkREWDaah9ZnXO57PKarINAW
zuniGqPE3kMLRu4IUFJbkJxkVCpcbeTc7GTFH/o9DgJbYEcLmdCrk1gs0/RHSmjogJgozDGs/6gI
O7NCT3tLluMjUuoQ1nvKI4nwtRNSKWwH77e9ge7/ZI8JRZgVM33Do16uYLjWKFZULIaDVCYWc/nQ
nQNuz6I0u+6Cy3rV6b7Qc8ALOmQBbBrUcVHDVbzTuHvtDjSge2O4k9nNQf6PMYh/3D/BGq8dK3sc
JG9yxjKEAnoYS+2YpGLrKAvNkyAjeFaeNvPM2ITJvUZd9/uftzdPJvi0zjP2XlA2VscvAadagSf/
kPY3Asuq+9F3SyPYQBOrQoO8vPd3Ax4d452WDM4xPH0yIsSASyBG1E9k803MYXAWUWMTHF4S/wDz
/2ijFRPatf4TaKUaCeHHFnJG9U7NOQf9c4qxstug2peSHrjgsTOoefhGmR3f/wzlefOjNAFxXPuB
D3wt37kDKx/fFB6YgvSAMjPFlByAKHJIBekmQ4F/th0VJXob9kM1Wqn3vM0Ju9LitsWPNyq885CP
rYVtDVnhYijEPr6gkjXldOcVYtArozc9gDIyDhYGOhDcCGpStTI3sRq/pcp3zwogL6Lqq8XpoxWV
IrrExKARPDyfVutU0BjrUTt05TUluwg53bg4I8MF5b2kKJVXMPdDzDOLQDWgr19U3iZVax1yJcDq
TQy2MAuxhln3ubKKJKrBvZilSo8ZWMBflWtInJEpSHAIgEIUySO5M6u9hoG0zEuAortz51/u2kOd
9HmhXJboJPX4/pVyWr9ZUGNjtmEZ+fvE1cy9CQIrL+1YctZJelC07EI0Y7Oa6/2foXlcZ9FnR73k
inCcPMMSz+r/vKvZttMfBBxizBbOTt9v3m+xFv0gyPLsjZpj/nYYc9z0XoSlfJOVbTd/WiH2NKDl
jawSeJCOuXPp1zbR1oucIhoin0gN+4p1b8fC3L8hogOZXm3lUOyrP3YbePdQELrMeBHkkYnTc/x4
7z/dWEdywjD2NfsXHux1njo93B3nSraHXoV+Iw1OoXc+TK9ucpUfujSX+6M32eAebF5qNYQJ2di1
Ow3nbV780hjxWXx8HSSw2HDIDddb08/hZ+BUjRkZd1ghYHfUMR3L3nhPZAWzFhGoFgN3LuBMIKEh
o1rpLBhRT/oMti7P6/0nOFVxcct9dULGLblhsxhElpIJH6o26K5z5JIlefb0IhrBBJP5DlkNNtHz
bG7sZKgejD1kxedlW1Enufb4wcMEkFtT5WQwn7Ptz1gZCgr5rtgBmCE26w64gVcKFkWUlAIIUcWt
x39xpQPwOBc7dsNZOcBOI6wHpK0yzz5GmnNUb7QIsd4uJZlbkpnR1qTCOyFx2tO3AB/lOFY3wI8c
+/SAZyCC71v/f3hJq/K0ZtK3hZdJABnCtmDyaX/5xl/JjMd6BxIiHRdewRK4EzaNLh7wQb8230SB
T9TeEByC6YuToClBJC5BfgTPaLh0vE5/KacFbP2QeqZPFWjJmzdng0db/fIwVzMHMBCdUa4rrwkF
Uqp+3xKwV8PHpGG2+IvwzKskY3qZts3zqB+gcx/vOFw9QFB/hTlkZO2AYdB/PBvA6xwi43O2GObv
OZuGTRvysCK/nUKylgxRrTkXt85LY8X4EbbWmRgiJnwmLFvH4KP8HtWpnEiPXDpVTNYXo4970v84
y+PyFW4324W7YMRMNnC2FKMOznTWEzi1xPMD2x/stll/NJl3Vn4OpNJP5oUTJTjpSpi3sDGMG1Th
UmeRtA73hhFnCASPNBrrunEenfYtkHM1vYg361xSpIqaGr40CH0wqRDR1bI8SJXlYvAA6xoBtawj
ugrZMCRHHmmZAP7fPFE4JAwB2+3MlWXfiST6+lBpaz4mG3lPm7XIcOu/67SStnYmftZh1GoM42y8
7PLpd0W/ld6kLKUnZaocTKOxCJYq4jOz5o8FHoC61SjQtUEnb+BnNgWqZzL0k72LDGuJSjOa0a/w
M46DYr+9jFFlBVYRdE4rl5Mi5JmLif93C32t26cJJzX3bXEXXhWqIeJ+Dger2xDYoK4ivZpSo/HJ
8xUa2ATBHenrhBAQX8xHsMn92hj6WdTDtCzo9fbd9jA0DvbqU8TzmWSOIqqiksHqe1VfnNMBVAhL
urQAW12hM61PSIz1mcHSfuant5Q5VaaYXH1knx2zUsg6kmFppg11lf8jhWPpqkgvJeGHXaqKLa18
5YMRU5ticZceGuLplrl7pPgTaIwtZRtlybmpPp4rItb3vzLade5sVBy3YQLvvXyaRAACi5lX/JYo
WxJBPN9HOLi4woRJVSG/rFyShKjfl+dOqESDXBfO04rWy35CpSs++271sNBG09hE/GbC7hS8EvIH
Df8msQeDsimsvUiB6DhBHIxuFUmg4OaYPPx8GTnzANe4cknF76xHWMYmX2G2QK5kKXhv2U1u4BUu
cb2rG4+p2Ie5VqwDavGkbskHvKTFlQiPTFtq224abrxN3rGR1T3BVZ56XqQJpDYdxIRyVDERb39b
Vrvw+DBklQYmxzWa4Nbfy9cqFa+GBDjuXPC7b63B9I6iCZBogExXdnlck330HQW2+Bwr+RMBTduf
Q7mTmc31f5/k0YYt4ld2/rjsDqAqG79spOTlZtB4rucJ8ZCQmHUudHkDhjf5yOg1S3NAW3tMbzsp
Lwfe025A1j/ffPLMA8pBoPUfsA+USVm3SDeKzReL4KJzZhMANkvOw1M28yuGCZW9cYrD9GBd4ZRE
MbfUydIODgwndw3/wefsYEE+2F0leDxj7igb4TGI1Z+qVaqxZNBGgkGdFapxQHNMlH7fN26xziMq
IrNwfs1Fyt+R+lmaLc43XPZClHI9qjNce37KcCQEfmcwApCvn8oo1Nd0LhUs76qCz+75bpq5NzKE
UbXNOQtFanUuXoUHYm/NI8OLscIGe2tGO0A88bV1PYupdl9/OG5IZpscXn6QQYTF6bYt7gwcQUyr
zZGeO/onh1H4Jl1NwIVqPUd6iiPTnKnDHYmx4MXyK4YQLiNn/2KsqWJDdrx5qwS+2fUj1+Hlsudo
/o0GUarKdsI3TtAqvk9CwxtOwF2hawhG3rUY4ZX+lyO/T8nq+aqTGostE8kHxupjdQHavPld0+IT
LCLeVy5fDUHv1ND5iqG7xKGMvW9fMF3rAQRBy7/8NXVN50cOnkXuQhvZFFMuv9Ns7rcAOsILKRZV
CKLG+AV5aPBooNpsKDM2ucHWi3FjSLCVmC3aSmHFYDbr+BzkxD9JH4AxFhxrzkuBr5BVwLQtdy9U
xW5VdnGFFFfjfpgD6dzBKW5tvysmUGSZFciihztgqx+UJNOelCEqS9c7WaJ1+7DUvo5apyr5RSRC
GGTCMwMcJclqHfHeD0S0nseH9PgDWEtnuQ38tJab1zU/TZbQkmQZvo5DTHaMt7qxyIQ28CI6B8wJ
M/+C+l2LDveMhdOXyquSByB2NQUdkHI1HJ+FrIknkYm8ZpWT7NtrnYS4LaztJY5qvvCGITbrAJBH
Aa/kD+8+YlvY9Kag8KyxOEYYUQhyYGDsbkJpAN0SaewGKq7bDDMdFNjUUC9Js9FUzgHFKLrBpJNV
ImQwpefmN4uAu6m4Ulpq9fLW9lCwzjFh7pEOUt6KGpra8hDolV3A7scOB6i5RbM8U0+XsyD0f7hJ
38dwREo6qU6VdgFuXC9ExvXHYiA63Q11HAMdQTP6QRXAhliMNXgZgaT2MAspgnUhzKq5nQ+JRwa/
GV+lGr5j1dC1DJbxksQdxsboxvN4krXlnVsTCANc+JVE4t/TEViGM2IjMtvEBGRP75DQE0wHgJ6w
myYjbG4NZHEwRgvQCLcJwys90ELhgprsuJhw8lza5rnxVVBO15nsBSnT2sh3K2GvawsaLOKRZKp6
MEzshI3sB+TsGW/18xciefBtwo1zKEjkt0Rn3aoL3ZuG76tP1vR+u0BdoBHNzE9vdlj7i1Yd0MGX
ecYJBxzVpl8m42zKo7ai/cjCepGiE6KneDk1Ro6uKa6ktZeYE25fQRu6zdiyBNo1CWvTSONECCfU
bet/iXspZevasjzVmXHImezo89vxbFmcLoY1A1gTPUNYOv6Yuuen3sn0Ijsqs6d9GvVFIKYeePg9
ecDI8ZiaIZkRYdIo4gc1GC6cTc7o3OJ6EUNr/zoc2/FWme3I8swfCTyI5a9jEmeea4+wQY21xYI4
M4G+F1UEcnkzwQxaYGuQJ57m2K0+df2ch4X6jRVAnBpw/cWrgBnyrh8ycT3qrAIa0Ad0hoOAK06U
OD8RYd6N2lY+5luEAlbwgjV3YItLF/ZanhL6F8uKmMcrdoF5SKa03PKOMCkzmp0b14rHrtQjLYxy
hT50oMOM12slXpvbSl+BzQosonRy5v243WkF6Oc0qw9oJ9D0OjLKPmgj98KGfeZGJk+GpUTLYwx4
N6aGjfiOhLDeGqm9k1rN8BKJdFKRkRdAHGPAvJYWppiGwFMU65JruR8zH0YbzHiH2qYXoNIOJm59
rakGXhEFGiPfv06uieeHeIOeRBCyMR+cWysc84C8LNfQFw2KXqZ5LHi2z5/tWAycSg7epeqWNNeh
aMHJFI1E4XtssPGzH4Nv+YRSawH+hpmzcwq+LP/mQyjjfzYautEpdZrl5bAtffHSCqJkkvx/NMZv
ZVG1gZ1Uy5wlBM2Cjlmlj6a6PtPibeqLYMdNplyksClxNROf2f4uhZG/lLn66sFTmvTWArpnBahP
1rqzNfpsv92h7nvdGDN5osLViADfm/6EOu+bB+JJ6LShbZT5lVcXw0NLHqggpaWvmJEldsEmmStA
xk5+bf06ykc3y/3zMkAAUiFyf76lBdCgEhIJuD7tSUYJve6A5SAEjjXD7hjkAIt2cv6FRYQVaRxQ
FPqPujbPJGmFo/ViJr3En4vnT8+PEcaYelNaHhY/EAW3ydH+StsJaxCud9gFLfx47nEhmitAUrBm
5hg89ecLvgxS1eQkrUjISSSEaTOhzbNxsnNx3gl8IO2cnHQ6qhbumQYCmrVVWBDdIQovUNAdTwFK
m9cBKUcrUbbW4tzkrS/ci1aq+uEZQq3quCrvmqVhP6jAdgx29yg3GLzkM5py8BP1xA0lIlF/+wAX
LMypFlFYTGl4Cnr4pQmsUMwwayq119XULUd1OQ9YoBHpIJqv/308aK/Kw0ZQBy9FA8TNlYxD6Pz1
SrSiwD+XPK0CS0vVaUBadV/CMGENgcJggQ5s9q5LDyveQZTNsmYrIKJ1oe3eQSdKu/NvZmgDLQY8
80MDSQ/XLeYHLN1hkdQZAfwLK+EkI9WVCvubwbIns+kUeBIL2l2GTrkChI9xsIf3ikA1PfFg6Qnm
4OKHJXe3sLZwZ8Bylem3IPxq6fkfQ7xoY6TzsGTYn8pMn5a7S1Ew/YrTNoo4uhZDBm52Mf/4HlGD
OmSzxwfS9r19+AcebhE+22NYS9q9MA75xqNG0eoVYHrZ/t/YgBhcbTTscprP1DHFo9fTR2Qm9dY7
7OA6RJXcdrAmgGXkpJ3M6YnEN4SXnhfMUe5B4KJKETVFeLhgd/soasv+i4g5kBFrmqeb39uj34Kg
tPuW5rUf9N1ZBT1Su9Ps0hGDiwql0lM1rmY7grQ4wH9UaxadKagVdg2vy6DLRR8FK18cqp+dKKu2
iqAoiEXhiRJcfHYX3KmeD8LWAuMUeiixG5WGbMET7Xk4B3xC3a/MPYA1N/iaAq+eqywGSgGksVLg
Om+5rwN9iW6J5kqOyMoK3XUQ+ZbC3JDiN+ltpB9uvVo/zier+zjJc7EhJqu0QkYk/79iIED9ASKq
GkBIqkkSuEBP0sBwqTffeNRauZP4Vk+NXDuRi/srY/HcJ14RRnPhdSGeCyJ0GVmbxgi2USnH4BUJ
T8+DB7cELuuQnNZkk5SWnQY6G+2oKA5jrj9A6mdZzmaFzPoDpuwRs6uk2zGbaWk6Hr+NjtUnnAXy
gTPV7lfdmaIMIAfumABirBFaRY4gjWPa+5gBIHleh0vmH8w5BfDcdNwKZifGcMGY0U+a1mKTyqAA
JivHSBED4lk5crlrAqzvFF1ICe3wwvQfgJL0l5gk0jswN9WseVmf8OgqolzqcaiHikVrbJbiMEah
a/kWaSDqCvnyfTSFnmq8lHWTnTIbSF0F0RaDM4GnQiFBtCv4EzVe4Wu3yRSdE5/hAl9HkriMnFdA
eErhoAnedaRkCTJ0uh9raq84VCWcaa//8Pnpkpbr+TvSVrca7LkO82NHbow5cXmQEObr3+7vLb6P
fIh5gKWryNf0g8XZeD60ntF096v1ez3Yth7c51FZ953yox66tbSeGjON8eBBzVgz7eqCArDlVBQM
VCfkjs+R9F0FVBraaH49vFKNfl0Vx6izHbnfQ18YWdkg2t9hf3uFS5NaMxwIzOx+u+M/bCP5S28+
am2/uNtEdzxelvnsPVMzV+hDrYtlmP48PyHaEK1gEHjGu3n7t27JrU0ZkmVWgFSoV7jng+ofZUTU
OMoUoelYLPB0zi0wDz5FYtsV6LyTn60oUt4aLAVN/324CHfYikEQpSYH8cth1YbnDPDBam9YbpyF
u7QbP5Hcd8n32fYU03M7o9KXffnYoRYSxT9xdzklI/j/xLAr63Zo02/wFW5a+issNePEalqR0kgk
7E3WXkgdXjosSotxUgGEefW96M83/Kc6OYfIrRrtJG8lFvzfUFxYwH0hESKRkWIn5Uk2FY3uWSfq
t4A5pmXMs3mnsTOr5mz951quz+EbjnG4hMOtlwI+r36eYjQwMwrUtCOZWdIPe/wiZdvSTWG5C6lt
z92yHAH53Qvv26BJP6EGkPjrjUt+hRuBtbeuuTQ0uOEdEv07WWw5HvH8/rZM/eCM3CTAjL/azXz3
9t7bCyyxyFbme/EE8fh9JG6IAehJHILKCpZvlglhtaPDnwi+lsjSijC6ui4XLMXpJKKhVT+McULn
zn3vH3hAybJfcM02sPnxj4z2Isn9xPg7iW1UUfsX3KNIWsN16oemAOfFlwZ/14Sz9tg6OX0rKFpj
QQgk/tkHolpZGJN6DkYZFZqXfuKnklqecf4BAfbU9rqZv6DM4BajzM2F2IcJ8NaoU9Hj1Vr2lOIO
LZNMGaSjCtlUMZbTXIXiSz3kpLSWMSL4jQ5tTCsWiUJiGxE5iSQs/6aJ698byo8AL32PJpWoSSGR
c9RhmyZj8kLzQ822n/Lyz4X2/zpAhnyx03368IcoaJu2fzGb6U4GaQxBhLF9wjlCeUmpgOspdYoB
/u7iIxZEYBZhAozz+u0dgJUDtdlmzpqljwjMhgNPijBQ5es4wD+fXXFb5CfguEEYYeRqV2iv88rQ
ef1xzLgxfXjPlhGaNaVY8i4pga+YTjBJOao1ZIfntT2OB/Jva5G5ESUXQXjx/xHfleupWrEVGVFz
EEDztT7AuaAp5II0VzJU9isrFFxp+Tr+Qp5fUvI95kDZ/vGEXUp2jkcC03HH1IVwd9+5FPtzRNAv
7xQroOHOCzf9r5z6zD/kTyyVHFH75II4BWTqP78UXAz7vBbSkUlICB2PPW7LbDFvf3vKUKpVQU1C
9QtvdAjJa8cclZvoGGdz+vKCe+aTnym2b0WNGHElyHTzOy1kDn1ym6QjkZerg0VW3VusMAvK9/bO
ADMku2tkWfzoSwKN/ZhfpXlAS4C4Oqe4CKzVVUbwnNQ122S/hk03+Z8aTIfXHNYCIImdNumF+qpW
N2W1STnCvPJpBmF17KSmHEKJ274sGzvaNI6clrw+Et4zUfszML4FDu8viHKNGslTAZVuTMtMxrJG
jGKLm+CIESRWFP6Y4VQSlT4fWEPml3cEi4XPo3GJjdwyqrGjDcIEF+bnNDgE+jdWmZwUNQlfBEPC
No/H/xT1WN/TJsjAzv2phtZJ0D0X++bCmOBfQ7/7Ni0TZKfdhOHF9lT985BkjE4QuJ72Z7832S1P
NHJ1Wof+5clqaUawah8w7kJbN2AyrN8nRWOFZ37WeW3Xj/rXDeRGkU9byI80ubiqXtNHCtbi4qOQ
icuHvwyIMLt9K2gJmyom5i2VSyxl9OvOIMg6thkhXNRwiqi51qzvWxJ70w5pb0XjUzjiIbShyB/E
iTe0RBYQaBoOMnUSHqeT+vzWe2saYnmnsSsxxihHtjChYKMX/VAVk1K9H1bVWrbsWlFT957w9hoh
Ywu3VQ9CIw0gIbPVIQN8VDhac+eFO0DKviZ/35iUfA+OtdlI2puicxzGl3xOCLyES96USNus+J1G
DoIfcVSjWXh1kSDKP2CyaDWZ2wvi9w9axGAt+4GA6W3TBiJq3iTR+5AyPopYtqgw8H6tbvP1znpV
hchKUFivCGlx3GdOmXPySGAJ6jZkP7Qeey/30cU4KLjc7cqWQc+1LWOf7qI/eTHh8PWcXTGr48BA
L5EFKZIxpJMc7jvx3S8B5wn0ET/eVbYiwdam6yduTeTFbga6Myn8Wdyk11y0ynGsqA+biymXPqO1
VihvTu/MjE3uc+ws1oMKmLSJojvqy2pRGPWdpUZp2HG4Xn/3NpHkngIi/dldXmS1f8bvQUdNjwLX
KrCrmSpVGQ9neIj/SlD8vcb7v0RAfAU4e862oY5b0rSgeIRujC082dMPoS7ZmnHEdjLV0HJxvuGl
4SXABtr9atOr49DnLO6ERTuMySqWcSY6vYXK/snGIpw8tul0Ck4DkXgpa5wTnXjGhAw9HsSxT+RC
xXimJ71iKyjyKSG2XAFVFZw2RjKwVDny+NySF6h38fjPx2QxapOZeGxh4PvezNviZCR7Td5gMZgT
vWZ4lRmwBKkyLG+baEV3QdNqRd1FaHV/iEhYjpT9oi02rxf8/keVAfVNz7vFuoNekj8W2sQSkSVL
ClL0MLitcW+gnM/AAseGF4Vchu/rgD1rWZ8rCPclHUBd7cY07FcDDxEiSUHjg0IZblW5JA+cxR+j
37i5LBt536IhZs5cUm7vci+dhZ2m6od0gcRZFZb7S0bNp24aJOJnbIHqv1P4a3LPzDN9tuvnUadQ
9kJokh+hTgPU8wdGZJW6+COojvzKqH1R0y4gACBOD18/hQBi/o4sIGpT+nRcSUNDyX5D5hHiZvrl
Wl2GX1XtrrJwJ/fpoiNCw9oR1ClRJl75z/vu3MZPvjc0dyiqWORweUmjyoc+bckh/4bR+wVDoDIc
y5YZUE+UJReiGbXpgu8TauTEBQKzr87FKMCpBd8xxVSTsbpwH2p9Xt5M39ANfMw/fOMtIVFRe4l8
i7K+j/l3ywKULo2bPTv91yVzjVq54fLHzRdIdAxiK2MyZfu7zbl6MU5m1quoY/EQxHEqL0zPKhw2
qr9RsBribCvFSem1FmH3kKhrgm7OJ7rgQTUWTTzwJBxFMhzvVibuYW7DgTeD8wl/iMRQbb6klOea
pi8aRCSd50BSR1R3qOkOXfRhRVVqddnREunMbj3rcZ66LMAZg/NnIrZZIksONj1cVosxwTx8zNzt
wt2ik1QMj6S8HBDQYf6eKhdweO1WLGXHse6vm/bm1qHnpwyWPbmjzCuOKSJO1jOjHzuDfUXGoKzl
2ag6v3s1oQu0kLbY+XKnUicmFLJxePIwSxHI3jIVPk8zlyJsoHNO320k06hXIFkfpN/yJi7TsrNg
2SgWp/rFxxJWUE0zGfBQ8PF/uf1fczncvyCIwzPglAINgS3X86pepkvTMkALGiTluI7PI1nJHsTZ
x99tq/V3p5aV6UC/u/tuaVmSjpr3nYc59AjTNBtdrDMNrN1jX3fJTkbtgwa2vxRoHyiQteKzHm+v
zTRU5xbZHTGOHUkbaf5C0PgcC3LMydMBJKCIVQXfQZI/Ff7qWoCGtELWQAGAT4B5u7mxQD0WT3oq
buLgCtGTvL+uqOUh5NBbX8KvgdOzyLLqF8fr+Dqh+FTnbS35ufC1a8gGH/qTBAdLanyfeJpyhct/
oqbhUAB4oNhXBdAl1exeu4oxJnrqIPi5vYJv6FuNMqDm0s8M5XavjnOODaHqQDaQmOP5zzEZVn/g
vvmafZuwUasrt/d2cIWJEmtcnaF/lQbxd8LyFF7B1swfAYnuxEZayPBk/iBheh/YQM2XiqOs2xDd
clZqdqw1vp2AR00YU5895/PDhxTCYNsFA9+RRGCq2ZKvmMz4EyQT7uuO8xY5DdcZo514QSKqpNQt
IrI5naYZp3keXYoLLXN+8FsMeNdp2VIwWNS1prckgt1VGm9SjnJl7HVj+DTwsgrlAiZ4PXF8ViUP
VGkCDqMYwPggrB/x2u5Jn20UWE+pxsyWu/gNNarmbT4seZhfMfQglmOKbCkrOMuqeA5vH6PUUOTB
f3O0KVNQEGBhVRwcTH8G6mdcZlqnDHWjCdEN3MypTGV9KbcgKck/O8IS343xB1SpNC/jBDuKzSn0
2tWsu0ezGQmkQhu+Ku0XVnhJa5eIKGRlMK3wEByHCvRkFkxVRLmrQL1ppSFvEz3JBBZvpdAYNDT3
f16BI270liOCXa7z0W/Uj0m3NGdfUtzv24cSagZDY93livKz6/ZMCzgpj4+UE4+Jfj9TGmKj28jj
75fRQM6XEVASTRHutOZ+i4c0S2lsWohmquVYOjmswCXoF9O1/s7CRa2v1L7uFn5TMmg8YrSuMNfo
robdiGi2MWZ1TWN15aM8navabJdKjyz7qYSpfng8QENcKwsitr/swM6o9yC4wxygfpjTxhe09Z8O
2OZ8gFzupYG0qmyDbVwP5IhyNao6M6YOw+GMttQoXW7eZpsgkOcYXswf8oZaW1PgDjwzEtZUgEpr
eGkwbWqr7EyYBJbKwyZtldmh82J5jbTXh2yIvW6rt5vDln4R6SRm7rEL5Zy5O5MsD8AAKsriqza2
b436y/169M5LCXquALU5bUNMlQwd5dCI91UyXmZJneOVBEeZboNgp9NAYshkY3gmiFlk1KFmm1qE
1JQSTJHXidSHSznf4q7oBKMeScyf4QBlNp9eAp5eM1pZ3aXbOlvs0PHUs+dlci4lFzfQ69MchA5O
HUYPf1DPYFZJ//tYYrJVr98TDz+c17G5J7HSnWiGt6oZZ5lbuqE/i+Pft3aXDYQBU7QATey2r0xt
/W09ncxhkO5Dr8lZsXhVQpjYg5nU0ZgfCaQdQoPnGd88OZ88j+YsH77BOiEvFXPau25C98AWVDxc
bm3mpZ2aLPIxXJPrX9pfV/EM8j/EoWAPHv6ttPqS1okXaBWztzac4ruSl7BU+wDCkyMhI4ZdwNB2
hkVN2yUGQ8C7ivE9+TnC+gZ6dihkqh+srq08b1rnxwuS9GFLPJtRKxvZsT1+ZT8kGxX53IsJglNu
up7eAXKUGnmiIYMyiYcVZGjQrQTEk/tHJdjrvUevFD1vkIEkjcA8kflHNr0tFpBe4gsKhnJ1QYZE
IYDRzHpsHF9no7m37MUYQ5/Hp8a5DRy+yzMbi2tgZzICYtGxMm+l8/ZpsbZpvrEjoNRIJxQxHzH/
vnccAN2Z+HOzxo6fEKJbTy7xV4khSHrNwkqj5MuK8ely7cEJ4z5e05USPv94Yte7WzTlG1kzaMfD
q670wbud3cy3cTb9Z5bEcQ4uNh5s/5ygBQ75VWcSyBDygBlAXFOkOZEppnpaxNBLaCzrjPlgAdiY
/PvVRnO7TjWqfGaOVpGdA7jJ0wtXbSg4TYYg71l13xwb11KxS+OqkRCeqBNqIvQ2SSh304eTpAyj
sgItW1MXQfx3pMJYsEAppZPH1sZEVwwsMx13aYnnl6OQw7dtLVE8bL4g/xv7KU1rlbggXyd1Ur5c
UXGp7t4mHbAUQj+ELnfTPHCuPEKC4sjQeubjUCI42RR8BgGeAYTSp9l8PstYipUC2W9BSmK3MFLP
rLmMBJ34GAyUsvA/7DpnNl8M67ngYEaWFICyJLnLYp8JTy5LNpM2JoNCir620QLNxeas5Z7c5k5H
fMlDSCwqk1HpPesKK4KmEBKdrf5i6M4TdUPOOqzghEPeaPlyzrJfyjaEB01RKld94KHKGvLLXDGy
lf1gkRJvTktsu2YQxDMeErsBXQ74xQ9M2YhTbCgvNdqo8RzOScwh1iVgemTYjuZfACvHISoK/1CB
mNen2Ot1e8XFLV0881vicnBgCnPrJaWSNaKQsh3AAigUKfN/MtYTm/IF74XaAjFnJmS+CsjZ8DL5
DdyLG34UJt2aFhxrgfsy06oodf80FL1QEAB0A8zwSjciDSINNRMafe2ksgfScYt3gilC/ySwKQXw
80bU24AwlbQKNoJq3chQfbfFL+Pxn0fHm8dBXWF/9zS/R6/8jAj6UdkPQ+09pU10RAtn0NPLJz+5
jZ6xT819QQUVVVSykUN7r7/VI8SarFBZ3WUwmEDRkPLlWEO9ymVCMpm9PyU4ggUq5sxI3MVS9F9u
H7d0BukhJS+wizZ2rL7HR87JtjO+0GPEO1ziu+7nkaRwFwYDlGM5Ha2VOJMskie7Q9z1kcFjTCJm
Vos8jGey/HNtL0qHAl2qzgQytG17kGZ+9fZ+UN4AzEk6//ziFlejSz+WFWvAv9ZOFmr6550C5ZGr
5K3EY76xZCEG//E2+1ompBsAOkDhXHO2Ky592yRHKZ5MVd8b32WOFbsIXwu4EeBQzyqQUddS+Wv5
XVmWgwTdCOpuDoDiLf4ap4EaMEvVBQyFz9Y2NvgGLR1BboZM47FKajd//XYTH6ymDP7qfHgSGlQI
G7CtLBY2iA78cSurOqSl+cLcuhmmCpzEL0tW+fxORGJtzBSkdfACXBVbfQmaBBO+GUAsz1b3AsMz
8nh6SZtg3yHEVs5Yq65/RHLQ/vM+jN4lNbHlrQprgMlrzy3TsjD2ETbpTZKSvKR+ZAieWQQinniU
9ezkzrHr+9AQ9lLhkOJzubyLrKWUOIIn5Or6sfbycfqbkpNqPwn/5trSP+M6wob/GVuCyzXSrN5N
XHo2t1rum7II7HwDuecMBDx6QXEn44d9B6RhpzqHluQhQtcZjM4m08WdVUNS+iXHg4/7jZgOnPsZ
p0X+EuCCzlWHrVuVdPnzOaKxqzlsBdxk4hUwpa6L8DInqOLIwX4j1HoCEiRoe0WSsk4vVPRR9B2t
lHuIGvsgQJh9jvI4MMY9rgPdFayo9U0b+FNMk3pxn6lu6A9JeDGnbg49jRw+72Of+wKWokRhmasp
dZ0uFyrLHpY1ILC3BmkkPTTAP87GzEZO6Q52JA7/6e48aeEa/v+8+3exk48of9sCFgiXjZMkt+Wz
DY501gT+iU48HvRn7wzV3i/8yVVT6JKs4idtkK6EUk3BVFu4jZNmZwWeQUv3ISW1WzQ6Gqs0uhaD
IS73rjL7lqi6A1JmPXih12E81WTWbBjWHVQTULOJTUq061evGQPuiu5irPMV2J0jDqC60Jjpv3oG
lVF/1UDKaLPBI9fyHqmgseUeKtxT2i12gbEC6lCjuAAEbrt9vF9DWMsk8QV6FdZTRWqCkvK0avrF
nM4PfvyQ1mtCoqtMVlf6o4d+Kgu+PwRsmmpXPUTa3HK3pEQihZy/FqlduCTvBlf7R0YtkYRiihvU
NU49gFHpyRZ3FAKrvNPd3J1lPE62cXSsTZXlnQ9bAv6tnhASeyGLEYH5N1VB2mVtxv7rAh6fxkTs
wiw/spAv7m9gjehkcg3OgTU1nsAadxwthvU3c3AEETCXKc0AhkZuDtr7YD5kZ1B5N/NKHb5DNoCs
PUtaw2zdz627NRs0EWrRR9/b8+zotr2hWhzig2C4a21cjyJnKG+zuqoC6PGDcYqdpYQRAHT+gSCF
caNxPJwhn96eM7Lq9xxqg5gG5SheUCV1wZnP40uJnSeWNeST7ErZ/sekYLm15FvjoZWv6apxd5+m
uWjMEqcVFKk1d2MDkKNl7vfAVPjz2/TAXwKxxoToQeF9vb/ZKHleK8YKIoUGQgqMUko6IUB2OlEM
k3GpvLv419FBpXKbBxQxhPbkRlRUpswJpXRCBfvmU/1xyFyvxTvqBJjK+7sFTAdhnB5rHdyLVszy
+CXu7rCQHW5ZbRoHuujPZIbMemWsYQzrHPo5tLZZ+3Ke1FgR6XhcNxWDegcRIcBNoONJhdI6p++c
We5/miQjCSctNoAW76u9zSzjT4Dlw5/pSOl7ogjJQxt7erhVIJ8zO85zDGef2Qt1TLwNJmrnCdLv
YzoQiWhZ3EwDRn5ijpvSRYI6d6uSbNof86Ta7iE9KAabljEsRs08/dlWQ0QhcbZ4oJcacmQO5WTJ
WS3j4HNBvMZR4KV5rrBBqiBgxJy5YmPdbk0r26b8r6aLBOglh0FiF82iAusNtqQHQjsYVx+8yUOl
cqQ77cFTFQFyHYmtogXhrpbr+25FvOMcG6C//R5zcjeTihtJXAGt29oDVcTk+MYKSj9xWlye5xlV
Xmk6/DEts81xOmdrqqjHazLY9ucSQZ6dx1yXi9dMz5PTTGRqb1eGg1eYXY0W52pZenEq33So6KLl
VEIKCn5Ob4L6RJTJzMBNykdbkTHVDJdvz27jbRCoWfz3BQtjBrzwCNyxVDi+5sbu9oEQS4Qg7Deu
CZEoSY6gsIpCNJBAaZII9nul0J0yVfoe7Upjo6dj681yRRBaX6LKWI6OzdbwpRLsonnGav8G7QQF
Ut4da0eWrDfLPc92TnnXFv4eIguV60y3aPknz3y9FNuI0kyIuZRA0u6IXYheFsxmiAs6mEhhZ8wb
wGwDti9QAQI1OAyFu1Ya30891YbncsjuLmrBvSJ+WB4eaPFADwfiQmeTX+DVq6aeUtZTHDBymlot
hVWhqD4DgRK3KdN3xDMCpPdpCKlfnQ8WVv43UMBEJBFvlmW4A4FBxSDoDTGmEKfgi1vOMwqBKQ53
2X05Ie7Fawt5NT9/VVEL6zwqhnFQD5dvf+//DiOnG/hIqB7n81hKN9pGup+sKLu6ucVseR9jY+vc
UacbAcYJBpRxLaoSYASvrTfKlP1bEvsgmJVrNGqFthJmBigZ9CPHHN4ma1vDsHSdbspv5EkGwU3L
m25TpKac1w5ZvTvysMuS1f1nuMN/sSauZ9BeW/SfGJktpLgqNTYF30UEd2EaxU3WfpYqIR1jKm7c
As9V4apqt3i16kuEzawcrxWTtkGMUtCMFR2aDZ7Za6wu7wrrXHv2wcJ7T305E2thexwSHtaIy8hd
DDEQE9iIdX8Mb4N3a+RYYGmIcHramPvGPvIX5X1e/zXmcJ7YBbQy7d0Ry6LordzQdAY2kF3gpANt
TWa9bHXx2OyAiO2YXq0si8SRpQm+PsLNth2uEawbSAAJZNmwuUQ9mB8uuXFH5UnJwSreNAhT7e2o
E73nj5M7aUJGb9t0feO9TS0xUF+GdB391nRvf67kVty/EV630xY92jfB9wl91Hij+w4HdlKwa4Y6
8asQpHoBwbM5MUle4ALmiLAvG0iWQSfHaxijlG1jJCMV1U/wUXGWpB1O/yrcTunWA1oX9+YAJg1p
n1QKtti0Jjj6B7lb/bipsEFoOGOHGm5e/LQPekcA86wnFfzW4XJhQDMtq7/1OMBHKqNAYt4vj7VJ
5wBdzHPPU5tKMJDKPKsQ3s3pd3useXuMih1oiAN7+gdhSbcKvDeu26ySjUX8coNoBaRKqgaam3w6
9a0tbotnHqJrAk/zgddNck6Bsppx1eKETqNLcFs7gMXRaLZ2a/mZ3Q+nV7IQRmWS868k2kl2DEPe
YQ5X2sIp5AufK7Z5Gol0fZzH7VT2J/XWmqfWT3XvjKcYSW14B0/1GflynfqGKyc+xyf1rOS8DgkK
Ii73mmRYD8vi7XRIbsUN5nwsDkCICKjvycHxkd9Zub4tkIfPrLsscvKntNv2iqi8gDvWn0Ts6aCe
8yFRqHIYcEudoqH/B1X09HEbws3k9L4R6gzxVw+Dh8zafxGRxFL/whl71/pupoFi9F32AxwUFiBI
JZOkzdz8hGg4Tf4eBMNPFTcuvBJL60G58YK6ss9KUSr1wg0r+QGUrCzNTxAqmIAAUZSeXuSVNT45
5N5s0DHuDoV4GloXnSEaEdhoSu4qp+V3mTkbB21AC6uTUo/Sn5c2xti7FE8gUMWO5D4Zm5j+Wtxd
zr/KqM37qO/QhQ8LqK5EIxv/SBi0bYMG9CNcYpP4Ksh/8GD0Oeb43UOagoh/r3H0Zls1RSMmiUoX
40ezoplJjlkFDh0TDjuBVieLS5mtJFilTHUUojB32wLWw04HbbhHlgubWyf+l/2HlTrWS4Yjvo97
/d1A25+mrL5N0hh/ATp5Tk/hCEtuX/Mg+pyHhey2QfJbOctovsOuEIAifwGfDse6RNCPlE0jYy0j
Y3F0dn64tQNlh2f58xvT/wdTGi9NP2uot49eCxYFxCWyOACoUhcEOB6gzLPul508oy+M+gk/1XME
ddujjw6rZFz8S7G5H+nIV4VVmdMY0K3du4UqnecI3SKIctl6tJKlKPZJfvHnJgHsdcqOK5FsYsnt
sV8SFrEdhLVxVxqJho3/JOBKMbfrlowGWedzWVeRskzh6OwkpbNaptow/WKhAFLczorRUlAXRCML
RL7gh24dajFvaXaaovSeuY5l5vhuYiGLbflmGs0Zbb4sjSy67lDEwPWDJooyDzP8RhypEJdwx2n8
OxqJ+FpP9vTGJypptB4NNp6ZhVilR7jn9o5OLjDlpm7Dh6axTlZWLwdKKxpvzY2T7+UmUoTYcF1K
UYgDe5mpNzSMSxTrlcIbn7FAz839xUDTU+lBcWLWdiAElvel2fMYKdVEgdIh0V/4RkQ8+2PeohhP
4ECi5leTOJhVq6bpjtCXW8dVelZuwYHhwasfSXw5cauih8aerTlzLVYBL6up2BETcS2dTB9QncRh
WhYWxdp08CV9Vgu1/AfmTWsvhw9GgCJGDDY6LDXCFHYWjDA6W5s2cqXJDdi7wJBe1O3WC1tM+PA6
0sgZg7xG1DDQ06KRMixWsYM7V3vQUvvor16K5AA0AlAwUUdlbNIR5wLQivfWkRK5iR9FFiKdLHUs
uOYVRvNo62TFyq0YPg9rQcRYAAUOhE0hOwdfBUiwLcNmrxacHQRWjdruzHaKHmrIFAnq9++x/3ri
eYslv9rZ3LIdi50k9lS5gI058Fz6gYR8B9XxAlAC6bM9qgOlQM/VVyu5KEzY/J4UDZHza17KCoQv
YQ8GLhfVPUttvxSbvVp31H1pKKouD1uK96M9Y1be2zju4asefZVmlEPHj28g90YhKwcTnK72fHW/
RYdzWhZbaVig3HuRWHmJ2ECZsC9a3dUWouKYjy8AEc4h8cxnOxSC35ghh2mw+wk07aAtqsVgUwyf
RtBsml0qX1q+un7m5UBkH9xGXOtAwX93qxkt5OIclW88Re25VDoTJfRNJXKRxQLlukNuKii0e81k
UQLCzi2pHpijCXsznKftT53jhxiLuEVy4dDHNNPRhzM4PTCubd82mIxGy7qma0zCJOTxxonOoTz2
0JWG4cKk9xSuKrH69FGdpNQuflPTcR34kiwETYzOndrhPfoanv5QWEYbrnJLFYAWAPFQXru0QCUn
uNwIiRYgkMJyfLpiAL4VXltftHDlrkiOfr1MTF+554+twP/D5U/QaXnAxrQzh3uGLeOwKXP/6DSZ
7+0yJMHntUY9ecZdrGZ5fuiZA56LXrAVvd36UwdQ321GgnqtqZGagMbz4gKA1vv0MvQ655pr3drt
ABSdiGeU3uNRUcXZTGU6TRtiZkpf+Y2tIOw54HatBzTfDrMIaeO3cB+Lpx+utRV1OHje/8cN/G4A
m5V2vM2+dh7vl9JtVvFK8FtgpsDS9mtVoDVMzis0QpoUuzPmCyjrjFhxffgfDLrn36IRYC+2RkbJ
faM+hYH47wkguE99wkwgzsC8Ryzp99wDKM9BRHlhbPT7HfXUtrGU1lUo6ECpKnyERczMBJON0Fw/
fiLs/eCm1y9CKyAS+HFy0Yf+8aOhPfmNJB1RtK5PzdK372sg6r80+2rq7tPVkZWPLyrT/dYp244/
gXtz2PZjwCIe6wnKQGHniKzcub+4Fdxl0b48irfXo5rg85HOUDxHyOu8r9lwlS1fgbXCqhIM8ikh
KX43SCK6+G1hR0CNLL27ZDEop2fP50osIk2R1/qSrMEJnIqs1v0AXfrXFY6jaPNyPTiDninqTs8U
3Ud+PkkM4mPmww+RQ9hxZMDkCy5iP5VOZ99ppJIHUhpAGwZVZioyB0AX7hbFRBQ89e6Xgoyq25Sd
2PGvXsJ4gwLhd/a/CH4uK1UODiNm2eOYU7kbnwA925lNWRQBflIbFvcgTm6aaEh0i+XW1VKPnqzm
4/k0dI1edax8tq1eSTvf5Kld9OysXTKmnS/Z+v8l6F1RSZtrbDdWJzClQqyr2OzfGrOJlQ98h33O
FZACE9/RASeIU94CzZTY1N7yb3qjqx05+MSDq38hStBPiwLETY8+ItQP/PDUM9375G6fwD8VaD1s
Hg+29cewb4wrcTAr8iYMaYmrWARbwUqaSb9qfzqY39v8GpbeSmUksAsGcopks0DC6xaRCmDbBVch
wW41ZNdhPFwEzmWMV7IKC3CCe97ZP+94InMjU+616DKdxXXvhFJhagHbM/ZO3IEvaaQsPEUASLY2
dD/5r49KKimfySJzzf/kcNcLxi30DB4ik2AGYRynLYd7Yj29CxjxWbqMVKsHpSCv+Kyvl2MNbqhf
UbYRMpre+2VGCBCts/uiKFqome6qXtTMwkezsNYZn1oycx8JGt+vHpFk306HQvE/eyvgFv25zrHT
18P2vj5Y+X3BJfUqN2dSHtIZN5Zg6v9l7xP/9wgeH6QSb8ltaiO53ZRlGAzteDrWVmps+KptQ17U
u8OHLCTI/dsgBdsdfNATXnRcHhLU33igdD+PrEFJJlr0jLpPRKi8S2ur6X5HX1Fwft0LMaoUr8Dh
hBg/baBJUqULt7K5Z3eEpb/ntD7nnpF+unneUDUm7zFt8Ryx+FMekz1B+YV9NmKgKsUJzQD83DiP
V66SBrlXUN5lpWZTQElpdKFVNuK18lusuUzT2FyJySbstP0lNxLgS5aC2uUNZufInQTb8qEDYaMw
8G6AOVpI6ou0L18ZpLQVbbOediLeLqr9Wvc+ZKXL2n36Mf1w5sb7HSKwCu0VTN7z1maP+N2r237u
nOzqq/Xngoz+CblJQqtX1KAEIe8pSeyFEQGUZVqpma4Tk9gB9aM2/pLswDekaJ4iKhCAo7MZ/3+N
dFwFPI6OLhINDLjUnfFuRhNFVEo1Hvu/4yegHAp2OuWQFCNmWQY7aTAM7WoBLIi/LG5715qVwiGf
qkR4Ov5ZzvaPCk3hy5xplexLdiAZAys2Jt/Fs5S5bLK5Ul0UQAVDgVgfGgLfDbl204nVk6tdePkX
gAldfwhu5liIsFq0E0AlW5CYw5iEIyitFw/EeZERN34XdqVY1HYyXznMwiBh0DSfyuksxzAMlvma
fj3oQTYU1V34fp8d8rPU8QITJyKMDMUJNXWmOs7OwKLlcyBTHJvjy+tAjkuVyzRwzj1lmqIjyRqT
pYHqvEsS8rPrdwXgK6EHxA7C9PKMK0fFCW6RqpbXiK9+lGELmOXhomHSiUPO/IuZsFTeVj+7QVrj
GN9lDX0CxG8ZtIGQEahAjNbOrAMBCP/yvIDKI74aooeH1Sfmw99kNSNVVf+WshMKnsqUJ5wB+Hi5
5Fdxo3cGpHPEGKDZtpf6qQCorKYMJXhK+y/VPltUVsqz2Q0HuDjLbqEsTW/YlD1uAvcGNpAn9aN4
sMW48tDHOld7C7YoYR42TSInVachUYhBHNPWZI8AzPYUdkRSRKXEfZc7Y+MBA8TIbh6/yCE0+qel
8ml/ASYmeA1SBI+Az011RqzpYPoeXGyUlPFaznzT6Rv5XILTTlRFQmyBl3+MyCmBACEA0XtJXVxj
TIo/P3nqBo1PEq16p4o4Dd1UhMyOkfFY9gSg75OJtlzCbU59Pvsa2bbbNQtCGGs4HU2N+tpKP/oP
920SyrWESLiISpILJzEUWnG0WIs+6iwxB8PpsmwTRu+rjLBIXlcmAlen90tvNdBhPhRLIKrZGRhG
2KGUjRNrjfeC4ag4frbmkneVQ18m5WNnsq0jD9E2wmeDtNE4B+dwzcmIss5n4z0Lvt3qha8FT+uH
W6BC+VQO+Yo5oEICl3239ju77zIs62vbzty/prF0PgaKhWZH/DMutgZwKhHkShtd0rgQYqPohkBd
2prC2W4KYX+4KuID93ZftvmYHaQEG1uu5nyGYyZzh3GDgRN58ksU3N+YAAXSGMRKvmpBe/rJ4ADh
gD8UUi6BT3iZQiINODf0Ly54hfWOFYF56ELVGLgei6y1dMJxbIJMfg5VW4a6jxHLO2ZQ3e3e2nw9
H0mPwjb0SqV97lmwHNPFI2D93+bvUd0xqji7MHAywVeMYhJ1tFTgZqDlI4FGlr6WKZDnyG4hpQvC
QkZZ9tG/EfmOO9BezsiYADljMPhzTVo3PVhROPvpVl74HH8MOfWhTkivUf9/b9n8GTOduIpboAPf
RYEkEkLgf9RCplLWUUMyexm4zku03zB4S/JcQQU/wkT0l/XkCEi4zpXz7TQIdXYRRPpXfOBpGCyl
rGenPsB5EvYmKCnYht+ESba/0DlzhdwkRBIrI4/euNLznS373Sr31WUlAZiyIIRe2BYjARM9KJmJ
P124jxJtrAOhiFt53p8GPY3Pd7KQmqftbRS2lGkKOtaR1QXM+05Wmb+qnJn+ayXCVhj5azd5wYhU
HHWl6fPC7rNplJmM8qsbdDNbkYWplyisQI5gZNtc3K+JysC21MGe3OSXQZcWoNlU+7cPvpRvbwMR
Skj0+tfDDn80K+SMKZJsw0RMNFkl8yOrekxJ81NONxfwPViH5yG/WZdlbW+QlZ/QE7CknfJT1mfx
gxlFMog5hTPFNa8ZB/5Y3OIuEubbiXGif3Pq8dHC4yFClzWDIzIgochar8fXWofUxZrrTU0aYkZP
TH5OqbzqSdBsJE4zLl4WklkYuJ3BmM7n4BTbN3ckR0VNOwMahyqIWqIFFSzN/cNSKLr1gbBaEYWx
Xecjcb6e1Zk0Z0A2EB/48neip9XJY75+CrXQe9MnHJKC0yO/F4zKy3cUdqRkRLZnewwPo3L7Jm/O
5g0HIZ7jwRL+M7Jghhe04DN9wNG7VxyhdUjpOLcgif+0S4birY8EC249iasyYAINGTpGTZbx5lD9
do5Y9SBycQySqCU+iQfX3wY+rIh1tahEzMJcM9rCY34Fcnj3PTjQtoY4bzIQfG4/kuShshXnW1tr
pJI/4m0H6oZea2T8N9aarcWOPJh3NFLmFhx4h1LNuM52SGKx/EFliau/wfbAsWbbsXReTUSk71Wo
vQNhtKtGgwMSxpmOgPnbvOTKGwvvT2738R3Zd8nXXcKlTnIHtVP03d2eKGyaBoyiCMW5XhfoAzXP
JhHOq5RKTmAKheDVewrFvwPQ+B0GVoktQC9FsxbesznMm+RQ2V+OB46w7wL8bXXMxKQ5ZVuEvteG
RAFJQ2VGUxRP9jj3xdk8Il7w6F04Tl2x/32LvLKtNhiSw/+59/W1XYAZCfkPWwhG8T6ej8j1O1+B
gtQJhBTZx+/RN1e2RP7+7w8TTWvYPJdAy9pDA5KiJPO8tuLRyO48IZowjhIuDU7mUz8akdHOMKGs
+I/9dTJqN6LIOMYUCDetSQ94rK4JNIIbq12YcYn0yYHLLPDzbD54X1/SYacmwUZEInwuRJDS6e9E
+hN7cUguN9C/I+wlZ2JeRWn178qYpxhy3fbhOupBzTtEc5Sf9OVjnKxlJiMKWvTlUTkjSXiuvXfe
BHnn6ix1dO84pNBeDNlaT7h6NSKhKTjUieQ95V2D2Ya5ZwYI92/QFWDAl8pqgymhRzDT0XtMLl9f
dm5o3Im5sgU8zdnjq+021VEeGCcbNVSdnpKvyoncs52KC8atbhGAE6xDnKSDpCMZ+WzV3z9XjeB2
/M8zG5AGblG9ENDg2/d3jQs8+nu5rsVA/2jPfae+D30ZdFtC7kLotlGX//Fbpq5FajPLnLqp503e
5SERB9H7B4lu4juEGzuDgcYQ8aHe2tM6UQP/9jZx8+PNjs7uHQdVBYaECUgus/GeGA6B5GccFHu3
p2vhO9n7GabLrInwRvpqdQgNMw3qXQ76R/d3L3fSecl7YEqWVyjyD1ngc5xcF+1Cd/imMxqPp0un
IWDwR/V2+iQuaL15TqsTLbNfoz25oHFxHdFcpwibVacxayZQfE5U1NdiTwwmMMud/OCeKwYM+Mpx
Dh3ZysYhDi6Rp0YVL8sMi2YgOIyb17suCDhsfaBnSli0Lh9nxy002sX9HAWd4aXaUBKxcGulmE89
ibj5XQ2YpdDHrqIxgwuUryhZkUXy6GbxFlUhCirpUAuWoHwm0yxLtbjMqJ6ZodSCoQe7mVN84D9v
Xz7uc9/7/3Ht+YBt5V8VUdbxCom+1GvDc79P00WKxuaRVkJXAc+OKl4ewxCTHRD0RzThxX2gzpB3
Gf8yhHSmo6ea27/69TtpF/kEMP5rt2A9NtTjn5qdLx+syPMBE7SBEHFoibeCOcKZwcbsjgl0Sziy
0fEdVDegTe2ZKN2/nO0nN9oo5v/rpRMrMzznu9bcUwtl0zBW93WM3JFLL6H+dfiTTBFivpsNYSUZ
lg6ttNHQGIJc7hBdr3i1LGOcykIGDmGQKm6QuFWkSqA/GGq6WeHBbBNqQN5n9VazrMTH4fzBj6gi
83d724BCl2my3N2UuWC4kgR7UK4aMU26fBnNb8Pd5w2O6F4yTwOhyaonaY2pyoJW64BDwCRgAQQL
VBitK9OieHpDhX+kaIzPBFD6pkAYWsd8L9HXh1Pt2xzO5rzEjIeXydHogWh2BNsgwWWa/Tktk9cl
DgL1qA7A+K/CeSIzp5HL3lSMUIgswb/JU5IAqiDisUKgbn7y5Pxj8Sv2X3RsUNkNNh8vsyf0e1bH
dmezTwf9S+uiYO+z54emsMfRn2YOtn3fqj8mWfUlZdER0sDOBD35w4Okv7eHxBCVtydvc8j4nBVE
sAwWQdNTTruAlSSARfAFUMY1tQZJdmqxM2QKR7j37GErbh1kuCtGb9Hnq/qVCiwXuGK7jWFrRvYR
Pl/W9QMX9ck2aH96pzIIGj+dplkd2xbxNAgsKaWXFLrcUFSrLcOXjxaWSY/0UFk0uJ6uIuWvQF58
ItaNJ7rdA+3uPU/hTux7aLeGUaOLHiOPxAAGkhg40RwEN4ntjevKwLfR0lnebqEeRYxpRMvwSp73
CLcJUFhn+dTqyQfvn7L+UZDdMrgq7sW7qvFkO739kKcxy1uEi/AaMQp/FnztmKT3IMuwDHwhv6mE
ka2PdArZW9l5EJjvSpTPNEgNs6w9GCaG02oMG/iejfkI+MExJbkmGk28f360kVgneWtf0IbpHUm9
lPZZUMSeXs/Xs/RV5BCLzClf+sTX9JeSmbQjSWKR7OzdD4DpV5EI7kKb2Nnnw92PuekNdvAZFetG
oIynQfsnoKc40VcuooEhoRlmLArBGwbg81wyYyBrtcw2BlG5wN+N8o7HZdMRa0tGc2JgApWCRBh+
AyIpXusSTnirgoOVDMKgoKmeqj7gj2y3PnUfC6kqdXVSabsqnhBnegecRilsK3walxCFLj6O2v70
rBdUCuBULM41VxWpsft0tClrdtZZVJSOMoAL1JPnaN3tLPuxBIXbgUmPSmPqyqbrbCZI/5rFpmAc
TJXXGl63REWNOEkpGTzKGgOfD+96bzPV7R2FjS3Wra7G9zeipxx4cRFlICFNF2VPA+Duk3uHb5UU
oDPgXy38pDN+vLMx03MlD+r0Vx3wBVHfoTVzTFGOF1NnpxDm1ixOBd4zwqjR6OZWZand0++KcUp5
jwnl65eRDCXKYDmDCm4GxX0slKk1rw5RaTKz2O1o2Fa5ecGwqBHcktjQiu++Qo3++m079TGcNMkg
n3eeTLXRvJ0e1wuZvg+YJNvQYx36kfgCIzvHolBEg1G1oKf7lPR5K/STDYkFa91MTxB366vNpscL
Eng44jP3dsjhk5bUwzAtvlkmi3nT9XRz6CJDhGnRPdhqF/TbeLvV0mixn1QsKYHPBur/nRJfGr++
Pnw0+CSic42LfpvqKMDImeWTAWeOMGVFTzt36oMLwlKrikHpBAvK0lUicEaKir5DM/BJ8akv128x
ShBoLqY5R/1u/GAQEFdzdNed0lQQFp6HYQEVKGOM5BYUtENjpgZWOOjWCsiHbmnnbc9XaIqyuzMR
sWc+nnWa1WmKtXIa9BFwhtp84LI6m+kq/08JKo/fxVXOr/g1oG1eSbMP8vEYkvNUedMLBuV6otmB
5EwqhowdAlMFIAwdjcVImlfIBBGbGRt3AyhkAUqw9sWlrV+GMEGgCZMmbidnBsPfkXsKPTAZbEqT
GN7L6H4KT9J4dld/HF3PXeH3V/srSNy2a69NOrBFqv5dXNwbWBELT0k7LT8YayALl05UKyS6Cfx5
cAFg2rbbB3CDB2muUz+V3UoGYpuzeO7YhMsJoRGi9xlpJvwS8ASBJ718KNMg2aWe1RTP9Xy614gU
lFeD38fk3oAg1gDlOPykiBve7DgNeJf3ktuW5RBkoC7wY0f5zJmiRrT4IWJsCGNLeMoG9GZFHZTe
l31P6CLWQblF81gmOZT1WgwTQ1wiaR1akIgOKfCxftHAOUgzWCOBDea5hvHIk8cxniI2TS7nCtPb
x6N97I+NCflr17LuK7RdNCt8n4woeY1hNb385a72HuJRZVFX8lLt6RPQwLYrdWZ9ieShRW5RBJ7w
LKWY9DyyRSIylFsNzW0uRS9JJXwH2pfJPNQPPXLZR/+9t4MvIKHB7+dUJq/eOAfpddOlb0Q/vkJf
u0X6xVh+LJKUIR2tvUxo2hXMev7VgV8wy7iuzZj1t0KAr/4F4a47Nyga0gmOzI5aDjuJjXz69o7r
08qW5GF4WhWZ1fKSSeKsnvx8HcWzxBvFT8YV/OG7qaqFeDb4pcTDhBnCOQsE+LkVmHj86wNg3y/3
caoDzDQwF1ecVQHbeqg1ipfvap5DyO676k4BfWbChJu/nTlhrnc/E2GTwolePIeARlJfGI5RaEnp
nZhg7QB/sQriM5YeeBZsvlSXbTI7PhhWXmzUfrTYt292ScwUcAqci75z/AUU5Rb+dAQ/af6vEuO0
t/flInagHQ8yNSLbWUeYDI5d0ro7XfGrTjAQQkdmwbwy//yjHbwSWAFitUaB2qhT2Z7Ad4naFTVI
Lji+/Kv+rsqwIQ1V1zvUZNNToTXvUcuY7RbUmNNj031BIkJJADZ3s62YacyqPIdXIzYGDIGaeSTd
rd4QzHIAh8eJfGAnxfN1DYD6M9TWGVVMJBXcRQwHuOaR+ub1TFdKk7h3Dh0F7OaSjKAktn+csin4
H/yQDZm0MUc9lSrHzQmys/aXkDBWW4FJa/zJHmLjze/nkrGq00A4ed47giAIdXweWhVhUgj3Zlk0
BQhf3XBkBvxlFAAvTBbiEnZFlx5/BvN16/yB1OsAE6d5MDaHtsfh/JUMlGQCSPCHPgFbh+s32rdj
wki57W+188N00J+U/w/wD0pVyssOfA+z+cKI292pl3PyZuyzfjUlnbhYCb42PjhL1vO8cavKZLUj
ggOD7lhHPen2xD+gsklK3170OK9nHJLbAMPx0M5r0UhyGGAAStY6eNXbeqE1OOQKWhqsvZc8gJx+
b6UpiQ5Gg6FQTLOg2PDnAEW+iw8NMMsWHP/Vunt8cPXsNlXpO6twrIgleY7qzTOPEGeCxvYAzzhN
0cO9S9+DRS4iVwk/1pq9e7mWyF6WrPfWlO8uTKK1QoQxLCr+FN24F/o8F4K875dM0tFuN7szuJyA
1fgAdVBdxeuEOKJ6WM8JtAxbZh/qbTi2ODV61Z/IzsMb2FYXmeSPuREWH2onNNhURE05ObgSpeMW
4TdglY+OaRNBOqnjFEPFXV3O6nfe7pbSjsdSHjM+WiiwdG/rDjxixkofElsqeedKZoKvJGwz9SSJ
v0XG4Myvj2mvpfSyyzK5F0+TBESc4OwDOWDyVDmdAMKc74jAFPIyqaJBc0MNBHUmquKg+r2mjj69
xMoAWErxkwRlPBentPZk+CHeuvB/l0/A3RVDC9zRluCvGbHPksNRAxqUKdiWE2SiEpvBjeIXmIih
DGVy0eTiBKKZkOScMJfCUCUMDP2nP5O1jdgOMSi5Rs6k5tIbbvXN6FZlakuTGx05vguriVjWeejs
8+A13bJ9g465P9qtGPj/BJD21c8dxLMJa8xIXCASJFFfD/b4cpD8MvZQ3mMgVbKj79C+AO72gVIY
dvVcV5gwAe+Ko9E6p/NN6D/jbQwwq4x32HB2rQu374rzx7w8hjZxGovGWkouokRH0BS02nTkpO8Y
PQfysCoExbq8AfoRChxjdayBxR7sRsNv1dt/f+tuEtXI+5b8z2Ej+lSJsX/DYsTytXBrK8CW3Xq4
WmJslcd4oPB2OfvqDeEKka1Z0Jin34Tig9zMO1+D4gqBT2MODaBX4YeD6LhUxsdIZrZpU2A3BdDG
gVky4VOLNBE+Qe+7U+lWvXOP7wtPXRVsgo3BUVTqnco84yKKDhMH2z6t9sYTsoZ7W/pjOfgGmkXv
OhilJQDummarGnjNMvHNoRIZkT2zdZ7Koeu1wvDzY2EDyT5GUwL20M2R8TUoFvS91rukN+Bil5k9
BKvwmBymkCF3rafcI3FnZpEzRwBcXbpigGq0SUpfZWhaFz2CATXDkMM+5SJzLMYo9NsW/WT2t4oA
H31s2UhnbgtiMrH4wlty5IfSeFo6pAb3O176wtAfAE+M5Hh4I4L2ZnslhFrfeGPuQUXMuu9sNujo
Aa2cGR7b3QQCqbArEX0ijIlwPBZH1/n59hwNznrFu213htDMIXZTp2J888h8SaYXac0NlsZ2I9Fg
9e6DTX3EY8OQ5J5hUr2gQkEij7D4ntr9bRRbRsUocXKyMqpYqhkkYRnZH8JL2Gew1E0aIleIDQmr
A0/4+DxMuC4NPXTIo/Mgvqap4kRbYIdMU7VxcoFMg29YQXBzG/cgVSiJ39hNSLOUZp0XbPt2Whna
bJjuJ4W9H8JyyagNDNNURoWV7dRWNm7QjYUL1lUYZoLwI9ZRM0e8k6QIpuY1sIaWr+RXLaPq5l3S
bNZBChk6QyRaWLKAbpPXRHzm6iwiFRFjONIIi35A4HdGZX2zXVH81Fo/nkNONC0HMcyhtWJIVWOJ
DLNHHXKPm9jdjasw3IYolvSUQ6qhk/kwhilueauUvrdHnIKSD8EtW2jqP1PZP7sGEFEHX0wBf4RH
EwoiV+n4lpy1SpDq9CRd2ejmG2QsEkowu/XkEDa0lUVFNo/buylF3LIs3jF92wfwTjtnszOBAzes
se8OyB9Yt6uZ8Gs/ayTXh2rkEHp3W+Go91i7hxhsNdgR5RG/ZdrcPmnZ5uImYHYk5mM/O0IYhIye
aubbz4p8UpizmBQlpxoeHYsu7ZIKaNhgA+BALwlS9Q/kz03BSIphHLm01l7A/N3i8p0KVxoL7dZ+
5r6KizcJuXOJVtL/HbwQdsSHYYbyHlaugtobwjhSkwG/tkZ2vPWanvt1KF7AraFLGH7pMgG5F988
KZRmSvx+6zxPpCqfBIPqXijDVRsqHox1616fUqoQEhoXSuUW0EvkM69vKiY6ms0luzuHZ8yLyF21
IBZL8vj4KIav/4j2yiorgcproqoruQXWWFki62JoQdgYqygq6Zo0ds/qgRe3NPQzz6XfoKdilMWD
by8s+9cfVrQflsAjTvKSslUhZRpJHf0xKnfrK67u100EjwqvFKRM5o9PQ4MKKNTeKWiqunxNf0bb
8sKvPqGWjaE9Oip3SAfKmdb74B/29qAsClJ/Hnx5Uf34B7z31r9WLUJ32sMyt6RGq7B5CMTTM+Mt
/jhcs6b/JWca6ncGLsCRFbUto4or9wC5/kqUKJXlYQj4KkSEv4e+HJavc6avoy8rXUpLLU3+6cl2
SpJqZfujLAHkpf8ancbb3tnM7arLQSW2NPeAT8UrAn5iOCIo7RH8RmCrI09CWIJiJquqYZ3Jhop6
bmVoMmtnmAGYRGk/WyDzOaM0OdJaG1PKZWMocgkFfK7VSY1TxWPHj00SdjfGPC4xpDmorsT/zFC0
FlJukygz6DF3l678Olnm5A85NV+jXDhF5TMYJ4Akg639ORzAHSvowtDTHsdETHan2tTM6vAUepLt
Ek1Etz6jPvbD9vA1NyLEZoQvIxmtiJPEZjYKN+UCXI5knBSfAEuA9AX4gpXD4OVCwOV7N6VdPn4Z
+bT3ahy4pUspKDFZoCkZg8WvRIx8+vs7jGQmrIxhQfoaVluefTGD0bKTdni7caShPcjtJJkKIbfU
zZ1ysr8ovBHjhu9TVcS0tR8x8wBg8JS9sXgvnEerLYivV9+d3mXxDGWHONwZUCOUuXlpH3ECLK/I
17Nh+AUpYGaBf/U1cy+r5g7HxR64rBwlZn+1a/ibD5kaZRTyKSrupirEPaikGkevZfTGHLNARH9k
Tf9LZKWYzwvcHiOxYRTQZmYbVH67iwYqGC6VOocxclYVBVKdFza1UxQd2TA/i4x4DuC7Qk7rnVkG
ZqKZSH3ew1hi8KDnQGiGrtxA8NCj6yb/K+EBTl3T9F1mdtS1dStx9p8GdpP/2sTn6XTBK7NZ+h4m
miZhFBpck21a6jsEk/jurUooiGCANSyJ3uq3SaY82JELLB8yRVS2//U57YCBinrYVIQkVxAvVIJk
mni5HDUltL+pLwq6iFekBYYY6GOBtnHrZSJlktGoaHwSAB812ERI78yHTLf0mylVTHOXqsgf+BtH
hB78FBjISVM9ZuTImOG90+fpv11SzNEYOlS3zCAn76m/nDiAER8ZYwhnN69OGFuTDb0+xxCEvWPW
b3+i0vLZQt6WBrtp+uOIxa/cO0UieZM0EyW8Le2IblPYbQO/y14DzJHpsjZ2giwHPSBxkxq+1+Iz
9wEhbm3Heq0kKbkInwEVGDgwDbac7Qyc+DpuiKiEaYKZTsb3ll3r30EYzsZknGwP0Z7Io8u5OMz9
bc/tU6PD+ypk1ZcbFfO0ryilb1760tiP0DU8VN/RS8HqjS0NH+WF134gEg0vi6daNU9KUN90+Weu
XAMaln9r/oC9PnRQcH3jLxOa/Ngb7yXtEhzL9LaaI+RxBdISjW0phhZU4MbHvdXmxFTL5dGpWkXh
2a99F6F72MAgSll6zuKfAnxhSyzXhOVgYpKZvd3cDUPNwID3BCk4yDGupFVag5mOlx2oIcBepAd5
diS2SwnwwOWqy0qOIE+ZsUJW1Jorfjhz4Lf8Pm6yvfGVfyOv9VrCGsisNKR6eQla9ek63DYPw8Yt
Ckn86euWG7CnzRr+GycHOrqH47PolL3laBlsnrSHx5RdwemZ/ZFddOossPkDC0R+aQMuBqGZWYo7
os+QjYXXIrZVym7qJQsP9VQnSyqjHKoI4rsnTk9C0k2hH+ACveClHO9DCn/YWVMJpUYz5b4zi9RQ
SOw/fR5FN8Qne1Vbt/iy45aYAjW58PYBtBJWvL4g9Hqn/8YvKMqC6Kg+4Tr2LHrOn2W0uvB4xfXw
UcluMoU6j8bJ3r/dQUk9xZ1ZoXpu7rkQ/2UQk+OY740ZNZ+oLkx0/5Jqd918YFXI+F9+gLxMu34e
HZm96cSTchny0/MksHYPYwNo74GOw/9Cus0tOv59M+hapXru/+2KHDoKEBkduU/Tiy8S2c4YOWyZ
ZdjC5hIIr+qWNtkfVIqJ7WDF3DMYY1AXp84Lqu5+z8dyQSkjwefmHKDJ9maEf561cXGWm7QpuEP8
DdyLIJbFfaDFXGmxRL4vVl8hSw8k5w6DmZ1K7KUHhTrrhJCR6z8vSIYesg4gqom/OLKcjr4CoKz6
POKIP6e0OjJDQXeqykic+w76Bh49glZTmGGX2cJ27gS6GLi/Y3A5abOYqDLcNM6gf5Uq/DjNRjaE
YLOozJ7XwoFwilgGgO/+8dC5H3fA3LHkNRWsoCFOSD0CS9geMAxxolTLKD94253o76ZXaBr1Z2So
uzRxVI8toQfDO0ky/tLWQoxStOqrqokDEbqqC9r8YmpOfeONb/NnpgPn+xN9YIkdU4hanexl07zf
4RFEUfooXvLQX0Xz3Sy29DauNs7ZYxLUW5kYK+s0fuAOyF1A7SVzwU890Y5hxsPoRPqI1tTuClDB
qiYjmGGCZCQMcrE+ppCN55aNReizEW+04BlG8wUlQ/V2xTOtWpPeOC8/ovq2UGvNBnk1eZvBRMK4
j/chmMSrlFUm7mCp4WEvZIMRMmj4i4CB5zAuh8nsNa9WUBm3SyJN/4KCFJ/b42Lg7Lm8epPqroyE
4akpI6VemXMZerB7d1uA8N48Gn9JEQ4Zcl3hNSsB47xDEKOn8fe+386GSHd3jMjJEo+lbLgUHRdT
PSnvImaItnuvN1vxUEgf9c2YWYyygjlTjFSPGLjqaxUfc7GyrHsYCmfQPb/EYg+ygCXhfoM64M0I
Vn6tShvAErkF38IB3MA236+suQP/uv5avZgwGEqnvVeHS3Aesn12Zx2GDOU81E0rrrhXHpV+QSH/
WezP0eTJsSoQrtL68yuoRlJORlkgLmiSvm33bB4srC13TiP0YVB7L+/eblRwjaVHzQZeydfKssnH
4RLqUb6IdWsY5kQEzDhbAwrac/+DtrKSykhcezHzgZp9QFg4qLCbSZffl9XDgt1ssa3uXVDzXF+n
OPhj0sxyb7tL07sH83pimelZWvRyFCnJ6YJIIhjGR7OMnHAALzhq5bYRRg4JHDbNW9OOXnSrNGaQ
r/VV90zVMLoW7xYvR1swh6GxRST8rLsRyG/XdrGNLps/VwwzN20IvXxIjqGoNTEt+E7IOATCQdVX
gEcEgW+kIFw2v+UY/ccb/XnNhMa+K4wBGlP+6nA8Ct0T3sTXTkX9hhqDVLH7JaS0p3Sy1/lTbaaI
2AfwsDhf5GIh4eMJPMh1d6VOBJKQgGske+9g7Kl0HtGrg/mkrg639JoTPuZQ8DI7KizAn749nOnL
xfv1pJwWs3bHsPjoyuZpK+ctT7IrFBU8srIltDU5J8H754neHuIp6l4f3lMsbMDF91yhjOIu8w4O
zpAF1N6co+4VZqx99HrYfLoXg8yhRh4Bl6kILfvU65iuhgaBKxDa/f3HDOXOtW8j5mLRwtegaV6O
/e4KMkf2kdaimDJo8DW93okXL4QdNvxtKClTBa9wu7gIWRyJ6rSp02kWC9IEfZm+erBiNpTAXh49
80oQPbfK7viCDXovmR36k82VmHeXRoqvU7/8L7lPrDOrt9B4im7hzDj8FY9skt6RWQdSzzjvhOML
AfN7uWmrAJAL0poBA5yPD+XSwCg2QaTAK2qp4EBXCRqE6joQKQNNHTWoxS2JGUPIh4hN9xPiYrzA
GZYlF+QgD7s/pUGu8jDS4GdBXwyXwAQcpL2mXjphwovgC87zgwUTUfWHdoJpqBsFFwpesHGUIZXN
v95DuFTc+f1VXkmTuxalBcm6ahyRd4dFPa81H2wRuWP+R1WrIhmQ6C9dFk9n37P1gtKocg3F8kT+
MBaftBInzlTWB298EizO0UfGPqAcAFXd6RXzq/4H18MO9xHu/6/GoA8NjmsOEBtTMVRCDdQ7MRWz
Iko/R/UlRXTDCl7G68XohzWdi/Gwt7IO5tWXykIHiw5PnBebZdyXpOq7NoH+HJ1wiIOmhGi9+vTb
KRwzMRYCuNmnEOywjKECESrTmvDCCp3GjmQ6wen+F8hM0IwsmZ/yphDK18mUjdr/wNP7nZlBLZvR
UIP26/RvuxVbBbQ1MsMsBOsfSYi2AjYQuSElx+ihjkipGkgcnSt0uAK54tcLGHfqoTf7aRuV8XpX
9RxtdYz1msS5FQVzMvhOXUwaiT3xkblk2YQeosQ/qhwoi82Co8g9LXnOksJQXEYsV+RfrTSuv+5m
HbyuLlJAOHa1NKvd8wgR9p7HSnQ0yBAS2Mg4DvjeSzCmpVMYWXaIagTHBwO06BWliZ93vVSAlcql
1X5er4bZHhIQ8nz94TCrA3NWOOCWkJk0GiktVNM9EXX1TQfkwxmMurMOVq+2RzZBzQ0jOXICftXl
F9f0RKxF6c4GAjDtlV/FlzoVFi++w327H5Xaei0W9Bw+/kumrEKedwU4aZr7ZHZv641u2ofJyULh
eCK1QLwyGxIk6EvcYjoPPdTTDknY5yWbgF0SzaF68+RdImcethwAYCz7wV+lL2fj7VQFlBLLR0QD
D30QOrcTQ3lzu1GEh/VDhJbla1G39U0huyezANYhS1ebDSwG3Oa4GrM4o4gFwhyvX0mjV7Ix1k/6
JEuRV8pPAeb8QPXcfWTOyEbPMr6GGadPNk2jzMC+NRuJWkPD3qZuf6ULuGpItWlS3J1JL3XVPRtw
43uC0LXxtZbFd91Py19VTJtztk7gMc3ak86p1UFNjL34/ABChBVw4w62V8Xwu/+D/BuWDx4l5D8n
fKJKa418GzCPK9IBl02N37DK+4UGxpWzAhUintesTdAPaRtdj7C+Pcjs79P9hWCwD59qNi12SKgm
NhmyWQC/ri2nbdlXyPIR5zWOAC2rXoE0P1nVEHK05d5A5/YfUIJQ+DHBiJNPsZKcJAQfauLixCLL
Fu4OtetioTWs6UX7OxbdcUTI/2QLJpsUAvcdqML38s6UuiyQ8WO1HDOdu9nCWUi7UkqLGn3n22tC
qAqCqu5mTNiyeF/cTXlmcqgfKv5/NFOcehqpq+EnpOmxygBh15uzkHnD2Nb05k5JGjKMjrHgiGA6
3ZbvrUGJEdA7y/Q3no7pAHx9rlzeA18ZOkSSYCtSKHnFJWFKIAdbkQ+EBFr2Cjkw8i07cPNZUbC7
mnn4oGfoGHRwBvs4mpTntDi1/c0HYdYqI4l+tYBCGXlOherUB+yHQS92Ggr4NhdNBQM4Dg5MjvOm
XPq11n25eeg+4v8ldxISP4vpWWwAtjlxsLAeAhyQisgau9Y7c6QNI2lHcGWnK2qfcwtMQ/3fObci
uHU0MKUMrKu+PAbw2ri1DOA8Szq9+QG4dsqD3kttVfl0M3/f3++oWZ4A0R3MK/Ew1vHjsRgX5YoT
SAQqr5zCHCbWNLQxL9ZZo8sTbgch2t+gVftMRzAiJmVfAIcHTqKUYUUg1+sKcSNHRvhAbN/p0ipP
f50jWael+mRspuMyHFI7BRXvKMkGOgwq+aZEzrbimm/RbER5eUg5PaXxtwvEqZZ+lxQvC4M1/fCR
n3k1IJrd8CafxN5euajBXTwfdVwJvYSoLZrhiThTq3HI0nVl+U6AfcxDBlL+lHonZafijlMF9bAg
p/paCIuiTK1Zo2LLpGn0alWtlBCoGV2KXQV62QLxTYyFYY07Oja25iKw/oqBRMOa54l9iJWbR/ec
g+y5D0cL0dOaP5uh1ZILIVwdFCLsFHNeE2Tr+4uoK/qERqbmCFqeHZdQ9yg+p/VcRo2UZhb3P/eU
ZDp+yXlhcD/MoLlB7/GpX/zhOCEFiBhUbh/mqIFUPMcpEW3ei8Kb/l7B3ini6KAruAsx40CUv+Ua
N+SK8q1xLsIuvC5KZgHMsJzYF8WMnvI3q+D9odkMIUPtjsDmO+qdr3IxgtxbpGxUP/cKqxzpEVF1
0OmF1Kc7Lmmj4bVHK+H5f/5AEXv13XVBI1Yowg+6zytQc17WnX7OD0JxT7ydRLB45qhFjdOxejr5
Y3xzUoLn+//qvmpvPGuLIY7+EtUisa92LCfiMBO4l0Z/kFt3I3C/HOZReWfU7w4shplUeTXsZAPO
fc/fD4CWUTJ/q6ImKe1QkGQuZqfqqNL+axI2QyDg7SQ6uTfIMgcTbdf0YU+u0Py9rnEedM+1YUep
c+qjDVCfypLkcUQ27I0gdG/uE85qmLp65J8LNUrByaS/jgAjkFFcxjkxpmCS2cCBLxC6K6+tciGu
ipu/13f5u0UgINGyokMXttdzdllFHuK2383EEPGPbmF92E0dRxqQu6KTD/dPTlEK2FKW4f94E4Ef
kdB5BjE8hxMUv6QIyYwLtZj4FQ66aXkX7PmIsJ+z9D+zeR9xZ9UZ2mH1qAKzJbjrkAu9V5vtgmWK
caWbe/6h8PRgRgwTnsPfBRHbx7YipzwAVPqLGCz0oLDhyUEFBYsDzmzVGYJ+uDfaXHyUbDSrKtSP
HiNdrgx/67pT4deOdENebgRqOKRJX1s6gnbeY1Q5ntlOcC4bnyIDsHMYEhNyYbLEyh78N1NIuU1G
rh1nPV9+ipdT3+i2sAWy8MhTxxAEyNse2M2Dx8/Lu0eukKXb6vNc9emKs6NEV4uzFI55VS+a9Z1U
szYLXcZWszqOsCuldQup6djg+9l5u5p31EI81IsC5K2T6APK5amts0sCym/5mXHS+vlmXRArELqL
Ps8KzNrKYZsWhYiOE78ed4oWBcEEtxcSHoxceTf77UalEsLuGMAfSQL5GbS03pZk5eXGyegEx4OP
+bXndTJyz3o0C3/d6ke+jeH6za0voxoeF+Vkrfkao/GI4ZVngg7fVko4diKLpV76YtojL5uwka7p
jBsME93KQ9tz+XzamqXFEGKyzOMA6mxJIUvOMYdav6jXuRbMAH8ARosaao2msjDdjHFJoi5opNHg
LSxDDgKCPO4pZBaaJ9Zn+6zsjrMecQL8XgwRSy6gbJxhCX4M0Bc7DmEhQskHV49R9bXShbQCGB72
e7GB0uupz4p7XQERnKp5apGcScXvG1x5eCGG8rA/hKeWq4N25QxEOW2gg9By7ipCgQYWf0AJc9bs
X+BxU/PKLIAsVQusTCZqDe/uoN1huz+yvMtYJbEqlUrFgOrARorjmqOTHoJPIo6JMgLCSW8N1NRk
I7btLctd5ZdFuVYroufV+oAL/rMrrJWyr0PoKTpl3O5xyYYgYJqd7cxzWFtJw+yqw+AAJc1ELl6O
NM7IQn0bJCnzFpu2YQs9LIjIUxbFpqm0SZAkOHpvpx8VDxlRQ8Z/w8W6G9PgeHePdZo9RnA7EVzM
I19E62Jryw8A2LvMW62cNU3AQvDMLVTZdGB0jXMWSqTSqNTb5mVbDS9SYPQ6E14UhEIfsjdcXr/R
L/zf5ryLtbmThW2GNmCWrBnQrykjSQXhLVNneWdWziSEFv8gnowZwVJM+FOtSONNCQHFvBTqrFhw
ql42XIAAqDP0hQhSofRym6By0c/lXqquYEsUEnMNz1lF/URToCW3E5zK6xshbDqtvlxLVWuKO1hd
FF9M7xWWVG76cAFpoqlMhTZU3FmqxXZV5L/KbBr0lKKbC5tTP3CV1E2cEbIGdE2sWSHgTRBh7Brs
0ejkERSH4/93OCefmwSWf0Z4sVS7XvL0xJdylHcgsyFCmnQqU81v5Uv1HVRdg97Py1ZNYU0Nk5jA
gPe6tgBpHWMCRYzCA0G9uVNGv2Yc29lIRUr9zH0BUqzZ9SdGl4m7CQxnGLc0FzUZjG5C1hIg2R3j
rx8J+SSh1rAqNKIYrhA7/QUfS4nPpR4R9e93WlG0tcF2EO4tBbLTmxhcoTBCE+ylcm+78Uq/Af4r
C1oKho8qN5WBk05DNm0jk091R/y8OxUG+Fx8/GBVHcEdgmEJC1aO/5U2rflnJtLH6h+fyuMDKFz7
j0f/Ny/05R2GkLfDXD7HZnCf5nuKMkIP9PGpTQRcHWeb6hcfxelUNeS6qRbKUcR8gIF9/PwDJ7Zt
Y5u1DBzpBkTB1hUgDbOdFtk0uNG4oU7hH8VeO+5x7WcZ3KZ680bckAwMnyfuqJQWl2ayi/YaVpCr
XOn4HwO7qj0OWMXFo8SgF5aLNiIlv63RzPLBbZcg5WZggYkopxlR2qVka3O5sh/BeEVKOf1TA3GM
XB4p9kmHRnjkvJGDfg3aNNedEhO6ZchIOyIXCSbrzLqRfamEke579P46tpUAYppxWBMH6DyeU6FG
GDrNuwBSIrTRqtmtZ9Q1v1WgaI+JifRSQDpORSIB4VPbHeHWRKeIOO981IZgBMPU0PSeEB+Y6Ht0
N7JSFXa00CYGUJxLRGHpnysZFowQTQcIMIH3eApcKVGh4guwfPqCYm5IIEvsLhzV/E50ZG2MCAEI
DepOV4964wtz1XB1HJDENdaoY+xYGZyuRUIRUMeotYSdu0jGpuWBGY+mevusQjIKQBbdzt1A4kxj
CNOCxyVVtP2lmCg1tMxz6E93Edi/LpjgBzNnl0SgJ/58wv3E9ssoca8HPxN54nXCrXZNAyffazeM
i/jIZqLq/BFd9k3WeWA8zMej6NJBk0zUNGCJcJp9tzx6P38fa1yTBgsnwcDklxQ2p8PXB6CZ7DCI
F1UZbTwLde9Zv5EM/QC5DZO54YxuMm1T02kwvaAcB4+9rlwsj+yXt/5qwlbng8dDPdGrz4oGuvfH
Z0HtMO2eTEfclu7Jak/aWNNtHuwLt1fMDeRUDx7NarUgNg10N2Jcc8HBofvUi59/8PfGZ6hED1Iz
2bODTqONEDBq8mRP2F6Sos6oEdW1fjRwWlwL+/FgHqKIajhZJZvQjf5J+ImVue84eFwPSMPBr5F9
qDzcxFwl4P8vkfwOlo5l523cuFa0ZhWwgZcE925/MktfAQYvDhWGteh+4S9i4lcoZ0rIcK9mqhv3
txNFlmbcm6v+xpFoIkq2B11bCH3Ai48lBkJz2ZQtdv0rDRCKfA4klaP8FQ4wHd6OBMp6VvmlObLG
lkW6AsbIrypKpST8e3oBZyCare9r0DheEdwInWhs/fTq+4KurYZDXxxwbcT96TeOtz8LMBI9HzM3
D7kdxqQlyBivYx4UVv3CyF9R1cwploZdhu7Ku+rEJ+kXqH8y2HIJkHl2fCaOJpSIGd1ooTp2WA67
2ORP7o/tkT7ChroaH2vBfy1G4Leto65XtuUBCgSEo2vrP3PasXVzzIei+dK+5ygig2lT3Uh/KYtn
IvkwL7cQW2UnM39iojWkkYxAsVkXZZsk3TW58s2mgSDq87C/PK/q2hlruEM4YIQbwzooBSo/8eLH
hXFaexKOxTM1QgdNIDTOnD4iHHcVPL2zccoc4Iawz7MC+2uXMFjV/u8ow2BfzPlZtCMN07QzVgbf
wKzl5ABs1mxGOF0pDiceamQnCN/A+CRN6uv17Ns0U4A5Tefedpo1hz+mtYhGLynRPTq5SiUB6Zai
fSjuxzRJ6pU7790EMIC0tmj4m3AHOvv4WE9Fj33yxLhk6VE8UX1K75C+GR4ngUuyOQqzB0dJ+nIR
g7kv0sOSR1GPxUt4RcoSUdcacsfoM2GSg54TB7XAalk/Lt5Lds0Ee7l2o3UhgaUUHyYYiTMTVWiZ
5kCfKAlsK6j5aYQxQv6DRfcoEv24jJFf/CnOGYL0pu0LPxjMdn+V5l6yT7sPYVl6X5jZNKxGrKzT
XTwko7Yw3vWk7f9HxwB8K12IXYU4EY7bFx741x3qtlTCbaPajCWqu+LJnwAAx3xBaJE+29g2nvHE
GFml2Lr5PBo5LsB08LwzBSXnD4d9Ug2aqe3/4pleqxPrJ1pZ/kq1nyaY+Kxkqm1LejaZ70KLVeFr
gV7DrpVakvgyMzTxmo2gl/DaIk5V4mq14ziUbVULAWnwcMXkC+TAj0S8VkmW14MBJvJwploKq36W
bvgZmZGQA9ypIfR5UVuJQJbSTFwtJCHwJPKDcDRXeU9uunCSulotMXHEv/NldbEFXL0mbsgocy1z
W3W88jSQ4CbxS2TgonnDLSQcRG8Rx0WOVg3pCrdv0E2lHEqVwBqplHFHv8GPP3WomFzrABdYsk6B
rUOJoZrJ6hpaS4FmBks58bKABood+DcYhdC/CjvceYrunxb8HLsbrNi2s0KboqPzh7/FoJSmhW16
ZYTy8jVzSIciHEa4Ny9IkqtfU2+4SUWSFV8L2BKc253FZwhRG+SH2jqF9pzI4XfSEaPsfkK/L36g
pM2bEaZ86zEkASuP9QSbJH9MN1MOIrSIxnf86fk+5uJqPqwlqB/z+FxGBjKlL4/Fwx9aWFvMC1P+
kRwtVMCahTiUEwx8QSEiq0X3fAjNI3ak8ve3dBnAhGuAve6n2ciV+CGOW7gItJNO9gsIA6Sz8nwj
io+ZnA3shlBRvi3QX2ETb/YvrbDJIVB/Fg1A5popfnvobUkYNn6H5AudrtqnH4/PNBwYNXQtv5Ak
i4yA3BK57zlPXFuHTj2nvwCP7e3q25pvIMl4LBHBN4s+AB2rG4bTLMbvOQkdkdGM/Nr+dYeXATql
0xlO/2Al7Mik74AuDr3R+1f/0NAss2raoXUnAXqDa7Sif5DZp4cGkXpMy9fLtXZv0CmngYY0bCVr
21EsepCDC6vaw+G51fVMAYxmfPGJfdmJVA8AhU7p7h5m0vDzBLB+Tbx5khi5ck7NnCvFggJX/4D2
8OORr/un8LvmPyTzeLyuEi+oOCA9kRwPHEBG+avXPC0G7msm5KZqNVX4Vv5rfj/t2wIA5lDFKFCf
i0aBkwUNPuzAhBUAyJ52hsa1AkWQv67cedX2ll7C19WCgBsaopRg2Eo/frvM/PkYZpnfc/7o5Gl5
+uG3CzIr9W+X8fEhdL99NGzSJ8CAEPbEXtDgBBAE1n97hYKdVag2fVvolVJ2R6QYu0y8NztL8rKi
VQ4w7zLmfQqSlSuthoYZT014gdT0vCyKoaNoVoOwXNtwuZGCYsbJTBT+EmztZmtYdOi8mpID7FAY
Z3AL2AgrFtsY8oc5nFDpu/i+7ga/5AnaLYxf+9btAbptnM9ETYaxPPEXdftCM7A/7a7QHIse3LLQ
eFW7Nohjb+9nvCB5jllT8OvUvBkPhoEwc5ZLIGCgVYSM6gboTi356MM7J6FaarTZKzzHWQcpx1dL
sYOvHac8NoaIPZ0Y4d+bnFM1ce9QQ/Ho9Y/oZZGr8qW1xfP3pe3OmvgROrWZknuBu9xG+f0sXFKa
2hhgUDuLm2ceDMdLUymVfYGLxPvb5C+xTe4SaZ9+wrQFbZgsx41jK3skgaIqASxE2ahfc1fgxLT/
psNrvaHegECKL93aCRjAP88hFLHiNdkjWBQAuUQZImDjry1XRNw2SUVr1I3nG1vGNWRXBHmx4aUD
Q2lnH1yVjAoCesEe6QaUJBVlbb6yksAFKaXSu6irVTD0ZiQ91RBkMDMSg6v/186eXCwOOyWLmmiP
oLv5zO+boAbF+CTwiQ2BIflZfcsGM/QOaiK12v65w2aMoy3PZtJApsuckI7NnddUsL9yn/gHpRqx
BHECHJfhjp3xXgohzXKD2BeWTkoE3Mb2Ih69ayO4PNoZ+yV+xZdE/xw1RXMv3zXniJb/V0hhxWtl
mufU/xIZutk/tSfJPW/8Z2TlYPKkaeaqrmhXL8s3iSScsBopnXKQ9HbhfIVoq2xw3TnVMLhkkTam
LMlo2rDsGYpd7PJMLLi49/IPZRSBqnQt6tRUmAZGIlzuqeK/vo7UPKagTl35cTIQ5RQrduESbDE5
xJspfEGqcXBZU5GZGlPDtPtbVDGpb68OlStidoNPSjoPRgAtPLsEm9iZjedKAR1mmifITFvqWqRQ
a+ZVyIqR4BkuHVIs1iROlZgTFb0Ay25Vlb6ZC1bjiSctKzE+SyjfhFlhvJUosdd/17Pyg88JtyyK
LSz24n5a/qgcuYB0f9n9UOURBqHbmdUjev6tDCXLrHz2hEguXltMtdtrn/skUPAP8tETs8M/vEfM
hxhXSnFOtkjWy94p5qr+nScsUzwjwMqebDzFCcfzKjyVPX++W/V4de21Ux9buhz/FcdUD4zJ8jSE
8Znaannp1BBp+IZrRBlTUsSz08aIAgfNldJL+7u6tWDP+ywyonrsXm9r+MoMc0hfuGXRhPvGJI1n
q2UWNZkTCpD/5ayOpcDAIkrdlvrLt7SYif5f7lmYxfowMvvXOOBcOZedl0tfGivN8hirDrXheYF+
4dR8Pz+syyJ/xMxXmNnN2IEGJ4LJomYfgpZ7v/E/FgDAtp00jUzxwlecHBxnXDWY2NZqcWL2zj/8
4rlcQtTEdwv+6Qp4m8bBYIYhF2qcwvglptcZQ/mRNR0CsQhhpiR2Y/mtXnV5Kz8PmsNVoGVRRu/F
873GzLhC6AYjPxmzt5pSsow9Tz/iZNwnkUH5liGMZDmUlJyrcx4saUjG196DkhtZPfyzNkMJLAS1
Ck0V2wh6sAWVFDYJN30iBw4jo9glghyfFJboT+gSCV1yhT5hIMxxZD0Kkg+YOz4Xx5qGIGzlqcDN
+3b/mS1LpFXYrE68Kqco+NmCovqXqa1eutSIUlS6rwKeiZeMHSGcp5l8Nme7h+Bp6RxZ/NmnroFb
2cc8mMJZR+g4u/trslMwJBPfUayK1aweac9mPMTMxEkzRu7wt/LoFP404hb2Ig63OyMBvwL74KOM
E5nEJ5SHJOOoDChDzmOpHh57MTDzoAgaNbjOKa3CuqGZjbqsaXXGQe/SWBwtNs4Zs6FwsEJQt2WM
Ml60UE0HjTxRxj+g1aDyCUEbeRNTi/Wjts0D/buX1NnC0mzoyv9G5IWeOC/VnLe1v1Ne0BBnaidK
/c7yi6sTX/soT/IbTxnSAnfS3405FPHo5MuxGDG/DVERJqhKJyymUNcbOPVFwyzMnPX6bqqi4P4R
LSQc1iWKzR4ezQfTm8YqyK5KTaOAIJtTetukCq7j6m04yoThZfTyaKX0WW27k7DglaV7dzuWBMH6
jXRh0I2ba3sYx16yxdp4qn/1+iLND8Y4jRRrzJ81EIxZTWKsEyEbNcccDRQtoTGdRugMTTK6jztc
8paTfriebFAUKKvdslOkqrLWNbuBvMU2In4jB83rGuHPsH/t9HOPUeBGr+HYZ2XBF8NRqEJdjmCk
kdiH9ATbmLO9vJ3OcuqYe+Vyj9JJYitoosUlAiKLcqw88xCJ3Ff2Y4ugC5xrnTEASlYN+KgL0TqW
AMuCkbumooBaNGCmyTWRBIJ/ubiz07jZHhhYJxpFEJZPDQJ2SSV2no2Vtv4507GTZlJucafZbJ1o
dmvYhUECdKIdfZDDL88/lsiMEW4J0EV4tEX38MzYZr4n41S1fAld3kGg1BE6gDzAPvL+XzXkW/sI
Dh8DuUTntYy8tbANDb2/XjxwK8VsgLhR0Yl7kI7gHVr7HjllTKcZnfGgMXE3HvWcuEoxLCV90/a1
uhL4DRuA2qVWyD3cW03I6xgNMd9Pd7pcKtbsx7kKIBCRgW4rZ8iy+OkmP38su1BuMK9WIOVEX1e6
jHtRdekH4zC7qdC1nHxYPuf9KFBx/F4AQ37J2awqeLhi34YQppZjWjNGpO+T6jZb6MnDBFbdo9Fn
gdwp531mFa8vKqIOtOij3Qe5wRWfLSjKiVJHIGRPKv9RLKN7dbFQbQDr1MjC2S+sWyqOMTMNfv2i
2Js9i02RkYdQXgqcL3TnS/Ng3/FpgNixdF6lxh9sDuWGVdES1oFWsQHQnEhXEHqSktVeed5wcUyL
71rGQDuw7u4cHC7Z23D/dQQu/2RQ441q51oQUO2gFiNoiXlFV6Lizfztz5BTXWHn4XJNHD3aEu+7
r8BRQSgvADdqx+CaSSJ+0SDwjdSugm4pEyef8tjE85LCi190vPziAExC1qAFH7XjS1gOwLiau3LY
T5I08Be7xq2qZFpsA5tlAuo2tC714izgjVsKq9CFHsO9jTBqUdqzznGVaegbBZcD2ATSU8d75tFE
6hsbfzSwHjlWrUa3Y2CB1WCLJmPY0T88aoYEc0aazQQ7Rmczru+jYgnDcHAWFiDG07qvs/BG71wA
ZtyxrrC0zd/qmMEYoNgNyKhk1Xsbrg04EeVNkTaqlpf+zTXQ6QgjG+9RvXz2kgbzCnVDkAKiWrZG
Z1oQzN5allwaqWJdDNY4C/H5IVfhOgMK1IvKi1iJcDNwyZIqHs79/T5N1BGwkmY05G6bmb1LuIYN
WBwusYKvRGBbuLGybFHRNMxhn61ghq2PluLvYfo1sXbU7+IY4tkWG1lhFEuC5zjFwss8GIVamj83
xegmDfBbeLwQSfB9HDmRUe/CZYUj4rSOGWwfp8Tk4wPkNpBD/CZnY32/YIVxSE4PT6rb7oEg8Do/
1E5S+WkNOV8I3xmmlswTnjY+ts3NwQJO6wBhjFSEt760vsWm0+jYtmJhdC2nBk5gXuXpIgZb0uk7
fQpknK0vnWuF1WabIwG7iNaniQbW4j0u2fXrC1o3f9Y0IFwyxXvV9BtxnKXMqasSLKlldNZqvPPD
eackDaUCtbEJ5x3bNzY4oXIOi5KHCzVkSfNPoqq2YJYx/tHLHx/ahIeYVafyrDLX+bo+4rJVO2FW
gwPKC/cNE/WHNECr28bP63Zova4UkSnaM/g0kgvgD4vKn+iccJIjje8BtIyikQ1n+44W/FdF4gEO
QP3SBSbIHxGh8pweJm4CWCvZITz/qE7HOfUAaEq5I2iVucvAMUpA0vMgvO8x9RO/lquBig6UVSw4
mEoJD3JFKigxxZaJmL61fsRWWkfsGGHYN894yFxiJokbFHplW5CK94I5zwAODXj8ledbfjd3JNwP
ZA6aThqhsBK5DKUYbkjKSxzbno1ml3ZyLIBlZ/c3CRD0VrQtn7Z0C5acYcaxGGyK4oihv9/epiT6
BjCH3dGx8yi5jcCzPrJTQJYiODUjRaA5bkRjdB/LQssvS7OsvtLqXfwZLzUkHBzZMICbcIyHhuNe
shHGJjDMHisZaWRDRprKVAPGFPLdajKEoZcKIBv/EvcF8DJ6+ivATObJU3XxllYjBuwdJoS+D4zE
olW93aiYlhkzjAmDeLtLklM3QE4uR40dxhzkVlS6dWvkj1GFFsbVFQRrO5ahvkFbXT85x4VvVsLB
MrTz1UX6i4mMIF6EwvxZzgzz+fRROo5t51sO2gcLS1nA2JwieNQbkeU5r1xnFwZBor108OMeNAwT
8947jlAfBeyMaIkJqHMRMMA3/1V7wuDi6fZ0G07xbMKUPC3ZCkNg0GA9tP4W/2SfhNqJ9+pUNsuW
Jl7Yrp303P7CTQsES2LAsWdG10VevWWuQXV3UzM/oFLO3bd1K2ca46cNb5ni6CxanV9atY6RFhHQ
W+Ih+072QkrYI27gFhpvdLfmwH/JYR3XmTgj695HpnNsFMnL36ryo/oStqVNHQqcE4bvQ9t/Uoj6
jFu59ZSkXv7Cb5M6cHELypjBHcoICTnsz5ILeE4Zl2WXh7PfY+LVnNWzMQXBtRDiDzI0GNMVV/50
Edhk+DQA3ZX2vTVMfHbDzEon9ZBBj2j2a4HOwHiYQQz6EUFeNmz3sUVGRlN7YXdR//X6eztnGM/e
9wFoK4gx3try3Q5glUsiX98p1Dr/gy05kI7kiEoAgLJMtvVaCKLt8Ng/XB40tRmv9jIz7oKMVtpy
r7dVEHiSZyZ0JrZCrGsuMeQGuFDK4Lo/G2HJurNWGyy3XjW/YNBabOOwHPVkOsbMj7QwJ/w490fj
xVEG/ge8IMG9nJrN02ChbvViIhq/IUkwp7nwOA8QpG4RxpVOoQPKyF9hGvBKIf03d1jGpCoyccv2
GDucTw+KTm4m36nM3tctliZyG2yg6edN++cyTbhckICyh7ZjKfMSkc7NbfV4DfuzO/xIF7xQ76Dx
tWl1sFyNqIGMovaYk2Q4VINIExnQggbeaNmWlX4QrdYzGoEXdKriIzJRyZ1uVjrX8U+XvflbB5f8
AC1OrheXiAWw5ffA7ZrCQsd1xB5achuhwPvjk/CAz1lF2HrND8JZeGVqrGDxVuNXazX19KDNWhpC
R9o32Pv+ZoH3NZlQ3Oh/cIyoP/45tMO4Mhi5o2Xga2EW8StxMEaq5qF4i2qx8tMEBTQUNIIl9qy5
NhnTFq6cTGaFac/qCPB2Bc8xbitLXyVnS5Ovl+InZD5k6GxTlkx2gxek2rcV+++3QjlEdh7eCrIX
/NZqXj/zpa72nk7ymP94H8x32ZQ9dsKVExlqksVHy289s1kaq2p0HYPPAXDPAEjnU0u0LbfhZPUe
bBFNkfRYK+gm6PhI0T59DWKMGgbULk3uNQ0rPYViebjFneN8OItJ/X25zqwSXSeioHpoqRYarLtO
xWqXa/QQVRb3DQ9QKjlzR6KyKEwM74eSPUpJ0Gh2wh/tGH4B0Nng1sF2a2y5eIC/Q+UCSpI85Q1Y
yfbkYXyeRMLbkZACai/C8xNR+LvJsmn9bS2UudMjL+RyuhFiAJACq6PjsOLX99oN7MZ3LGwtCJd6
faAyfEN1cQRdM26AZWdV3LeaG4ai92XoY4QforcQumitF9AEx5D9dAXBgHvfSd48g7epyiUjLBiB
acaiYVMCqlmRKwJeXU19fHZZKoZoGhqflRmxc+OEufixsxblcQLx7Kk0ET53p5AuaQ/hZFJdYv5A
PuQeWrYbA0wCLp8yzSVlBKMjnK6jLLf4nXv+AJQm3SGghb1oDRfTR3b2GWi8tOvb5zXH9zK8wjuE
v7wxDUSUISMly7XvrcynDCcxzUKJSCQGVjZtMsM1ocDm3gxbsiXZ/yLbr9IEoZsfWHNRG3G/7QZK
RKFDmFWpzVoGzkB7EEubrk/ijT9erUQdF5iIkOjEwaNTmq/E+gPIQbsOZ6Epb1+BhuXy+a9ky816
CjfzvHOU4bKHvdJ7yxaDRl0hHxr4AZnBg7SQ3BkckTXU7QSWcWQd3oqATLCYIgwG5OaRL9ILbjkU
xu+2eCtf8QsO6/Atm68VBc7ZLdqy5BaDN+ttundOcsqoNYo/UHJMjKBCMiIJExI9DVls7fBPDXrD
SEy+tSh3WDt/qnX23PZZWt3C/UMoiH+YdwnT4yXx2tKwpfFHoR6QDyozFexj44uou5fojA0bZvdE
y0S2n1EkI4iRI3HmtcE89gpsL3Mdgvr6EH8R1rtg/JREquiQDfKQqA9niSXQCYMCU3zuYxRi9JG0
pOxylAgOQc+Rh8FnkM9uNcgPkr1qYe6xhgBVMddFSwtfdkAMN6/JVts2ngqeQZX9S1sMkp510Wq5
mhsmERmwn3Sf5rQ3hZ3++eaeXUl8ynGxV/x3h2B/UjQj38mXG8YMxboGJNc7AGNJsCGceXXFXvXE
0abPAe04IpJQ9glwLPWKdC2ifJMM847kBGEZZdT3kQSjkb6hbjG6xFRsbzl0Pb+0kY9yXz1eYcRG
mJVqiK4nO6pr9I0F3Wcrm+G012CRDhfrn2X6J6iYJU/4arnkmO1oUE8Bn/uu0ebksyfP0CM1CdJX
sewtRz0nUaJRFl/HxNzGuYwUy2fbSUnk/ov4i3OrkT4WGvGX0cfVM11aghRdFhDv/nKsWSQBmvpr
GSEzRNbDyi+uePPOMZtvzMt6qtQ7vTCPXoRHtK+I1bWYLDtfvpplsO2z+YeKm5phxj1uTbgqr1j+
S7sulKuCqfC6vNJV8UPyZWmxXXWiQykv8jj+JSqGhfNVsWxOpvEvsNq2hNlqQDmVPICiInahYDDz
+QinInEQs4z7AVklYuUROL7fprKx5tN8QjXyPJhpTZ5/JYn9XSpLT8+JYbDQDw+uXEBv5yMJi8ZQ
Govrw3SXURCsJ5oTWElfuw1T4HUL7Ki8220jd40M8gvIMRW9NQvgCzGwqjIlLkSQ/xwJ4eTRIk2j
rqIdWbuk+BMbgcJZWMHEnEN8Pjw9pbd22LQcPHhrICyF7FOtrTv9SVhfomYxdmioPzvMHbUoafxl
hED09hDszWsn2rMMUJlcZzRdDf4HNicq8GLvFZJIjMpr5ZG7xe2BLANb39yP6j6wdnJ/gCNlkhVc
VrDp5P3SpEbjdOwwXEfbH4JQcV/9cyi5jpI8FtiO5tveKc0KKo8TR4VgVZCyTBDljy/RTPNXPkbN
Uxl8T7B0HmE8lqefNLDA7EMW043xXnViA7enha3fZiYp5JMPF1ksWJGexxNf5JdjgKNs/Wb4eljj
+r8a97FHxnx67Cah1eq5+ufHppHrf7iv6vDngfUwBb2YohNsFm/2WSDWRHhX/iJ9s5kILaqCwzpH
4A1QWw7U3CPVzPQ5na0OKYlmNApBVulVCH7Cxih5IH46UYSutvaJ8HGo14v6c9o0pSjPpmkP2fO+
clug/0Zfwi8xD4n+rl3eoYjOFTts2E0LDPNSZQPbR2I0+QeuLkSN1ZRuO/97rZ3CIp9lxql4DJks
nbgfI+5P0RL0axam+2z+sN6hObSIyBhI+6wyUc7pCuVIKBcg3kY2aOJi6UkPnse+u52rkw3zNNSV
jMozZHHnuXR2r5TvZE0iqH6XuyauM71KNA9PTyMIAoP+E03sPq5NP0CCWF6rtkHMcNTEsXwsijdR
6pcSjjO6v24E/B9YffRw4GkWd940UhCFUw5/5ehT00R4L5hPRXZyU1cFa26mf/ajMeO0YsZSDxHc
ZMAdFgL/fcEqxX2TkEKEzsv9ZFfQ/iXipMnq/ZDW+OrWej0Z9+A0sj36hTJX7oQvgP8sm/TIUbbt
dd80HkqH1Qr9tz7Yh20g9NsYT8i3wBoTimlc0SOIS0siQqZAQBc8JJmCue4Zpoufj2IifFsD9wuY
mxbxvw7AJ6B19aXkV1CM9M4Xc6lHUuvfLaZ9Mg+jwYzQY0WCTW9AoHODngl55XDiDgizx9H88EaT
83fj9EhYg5zyVBunhpgum1wiH/k4YWlPCzNKX2NgUpvJ2jMnYiUb3XOjy89njxOpvQp/NuvkbzWT
ENZLJ80ycV0Rgx8sv6fskicd6NKwJ5fxW42eD3y1el3hgyY6Ph9u/LobVgS0V4SSOIM15xX8HtIE
/vP2Fv+RoNTnYTW5EK9qZxbu6uLJnP9RFSGn9bQbDHmhseEC/IdMEpv8XjJ/p5nL9iPKI6Rbnafq
YzBlRBcYvJO5g7Ff7d1miNpT/S9XDMhmf2ZyoLY2ChEa3UsH+6psZNPzwGWkJDoKbdN4j5qlLzzO
+WAUd8J641L3ukGuWhsXSAVS8uQtRzYDKuEF/d/YbH3dVva0BlT+a+jizuKhCXtX0Q3FhN3X0N6r
X+0+nul23UcUW7xpDkX7nUFl4atU5WQU7UaL6z1Ca1PjxjaXKygio6h9968RRB3HJJuaPcWL53GB
sJG1f6TcNaPMjeqr8AQu3Y2eit7b6b3Nfh+zuVDrCIhJ+6cs2JLKXVAIw1CW955rbRvlKj99ytiN
y1oWy8ARLuqbgXxjQP4Jpgel1G9jsJOTR/p2K0RJl9pFp0tO+Lp11w6J/mcp81mFt1JFX1/PTUIY
pT9NXG9z3n7JGZCkSG9NWxPmk554BLB7pOimwoZejsNd9LFPf/FEt3loedTY2sTteoL3/3gPIyMt
Nf9vBgKtpVlmfKofWQs0A8GslUKc9hErpqwjaQev3Qd+Dg4UYhfouB3xz20ED/RKSb4x516/sFs9
CDnm3qGYWuZTQ7YYBhFT04mlMuvJ9oKH9oZe3mDJ55ZTn2Q+OlN4l9lHd9K5pSYJwUKWsQtDwQPe
wo+edFD8i/YRIo2WllTvz3lvL/4wdihoS/43eUz3+ApyejvTjBMhGyWGVfYqhuzEzs705rXHUqZU
0BuiH5GxYBGaNKRUXii4ASaGPAEWyaXEI6o0cIZHw79pWuKcK7h+eNnsVb3K6pDknMNVoFg0/hQv
gDFu553c4puio9vHUYxG1iw+6lOscc3aoFXEwM0/z7Gxk5SMNX/jZq4EXX0HCiWJ2uVg27ICITD5
0kNiFPkPg3x1U7JHXFR4STg97iEVTryljAn1+CEDhtpvvF2WoiGZz7ZnRiM4J+5C+N81IuFqsEMb
Zrp9omvow3B7c2MN7jpvXFuHuQv66LXuImIOpUwMjFchv9xV0EAT8KSX+QfO1YHUWVk2kZ1yBdgR
QYiimztQgky4LaFmdMUaSPpFjVcElrzUwm4e5jbL3iNvajLUNdgpJMszvpIDUV9dG6raaDggnTHa
XDn7qlLIl4Yos9gzYmnilCu466AL1G06SCCZue3cBkwK5QOGv2TLlBPXNAcwGDnGPOoTXLq03j/x
ECEXTnkGp952+gjbTIlrNxzzXJcwABEKACm5i6zTRMkFS3WPUPdVLyWc3x7ciKjnv9B/lDRqFrYN
33pK+eYeZtnitjVsXnyggr0LfSQPgZWkkLxJa2ajQc9Kd0ZIMulRY8mD9jZn0ZAjPrb+ERgRNgWr
dyyQCFOTgvM0Yqz1pmzAdJfyIbIYP23BfF7ddTGs+6YVOKXULkyEtdoBftjZW3sZUWegheGnmjqK
dRBsQDEKFAcmjbFd51ZcoTVfXeaFMTuBrkBmjpD5aJ3a7OaijavX6KXhGFUv8ZEGnJL+9Rb8/hG9
m8IvI9SsJZD2t/T+Wo649mwUTkqOwNvmLHvsps5PetiP57FqmZB0JNChqZ4ETt3ItkbIQaHsOzz6
pYTkMWGl+MhAgcLH0DmbeuXHk0NaWCLMY2qB5ihZ1oFvgGHyqxoeJUH5cvvjMMzGfylAQdfkG0uN
DOhcV1vc4Dmx+vyyWw6g5jdRk1kdPUnNgzBcxETakDcaiLlunABneR7Z9D1EuTNGDTUlHYGAhb9D
jZGnv4Q5vYDbnKxSRH+IR7VJYK9gCvz2AYUdgrliGOpANW9WkPfi465hD3quEkbpmht+4sWlkRPq
6Z9jqCf/p6zjKqPCW0Zz7cWuWf4mw03PZdnG65Y4aXV1AonjCURgrwBK5KhY7F1IDbyHvaLBF9Fw
WkK0iDokeVubEds6CMRRp1+4oP3e5R2vEKwT3yVNvEx0QJrRIOlzsM8ZHXA5Ty9yR3zy73xjGSgT
z09lTs9pa8Cv8XWJlq5EPKMfpi3+so/6//54F26QSuTMdSSVzQGc6ymQpBJI5c0PKoUJHwxsNNtW
JtQXdDvCmDZSdA8OqzTacyXC2Xy1Xky1iVrbV5vQmcbo23BybsAn9KjJxsCQggr6xuNCJDtyHgxr
K7m74Qrq6KapYMaZAN+0XIrkKMktf0N3h5umDViRD9/2WrMqONcX9T4KPOSPUY6IiR+/zXJvf/9J
1pS3dodSQBu7lsKxyusCerdCMtDQq1gnoE3ZzmW1LjAGOys6kh6jEnKRQOtH4w+F1bn+ryXjY2o4
IXU1x8krLj+BV5Dtq+e0JK/BbKeFZvAuTLWFvUSTXAV2J2ZNhFBLaxbdirQNG2K9iNQXQt9A+qNW
xFcMGjOFiwgFIFE5DrSkyDhpqjqmJSNEpdcDM5GInD1PpF2QzvOkNusMcSs3jKaL7H58eqi1X+yx
jfFAQi/yiI0FTjHW+fBhCZDz3EMGNe7rGc4cEJjoTvKGSD9sTyCE130wtLCqHJc4XpGKD3a445fG
TIC+TO2aLtS+ijNgBb9Kc5x7drzH5OowQv9S8zKzyGqcKSfvEly4ypXDrwNNMNUzGFSwZk3V5rlN
RcwOw0Q9fm1DHTmhr6ROwiROA9RwMwrLbYZ+K9DuYZRP+tzdJ8C3jwoqSLE7na9x4qOYzCnSjCZ+
pfOruNqvfF8O9jrGBd1mBkMZiXtkAil0Yhw8qy45yZtAvC1kJiMKLEenCf0vC33YNVu2tE1R7yl/
156PTB30YHQrpNhVYMlhdQUqsTWxtOx2lOuhg2hlKgG7P0fqRAWcbD7SE14s6gCGilVSl6y3SU2e
kv3PJdCgdM1LXgzT7cH+OUF8kWO7D0bB7Dgt6iKCctQgl0CVm73s8cN+R7FneqmnzReUG9dc9trU
pZY87hnScF8kCIuLQqtd1ceThrxM6l8b066HPl2MSQwGLBeyld91JiFPqOe8+YuapYOuy+zSyOtZ
vFduAYKpjwTqkog8JXTBq0ed1OHQYXVmIdt8M23yVcPc/st2j2D3tP9JX/s9aaKnFuCwCDL/Jybi
Nd9/++N1H203PyFGJ6FGLIXb+sMohU+He7JVkNeUo3waXRzIekWL/8IqDf6+O5oVFN4NNazCVEhr
/3NMcA5FhBNqYhcGIxpwoVexrtP/wGMsM0ZH29i6jkj919G2+8YEL66JC9Z6j5afgiJkeXSJ78pZ
ffhW+wcRJ8phZVmOliqjLVWPSumTxwEPL2TeziN/eHMafSRDkzxY4cFmVhmpACa1FueyXMQAO4Hg
Msfe+ZzvKhZvvDZzFl+08FnaYDx6ftEa/DUKIAXlpZ2TOqs8o78L5eIzTL3sMr93IuIurhFcScAf
tNYszsTy0/CghqQVwj1kqNVvisuI9qqCK9SK8+1dp48SAbnkxgQ1Lp5jqD/rkggOmgJ6/nwqkRMz
0BFcDo778+xj8eLaOXUBrSy3Q7uqsAM+u3rvHNVaSUmYmIR6b49t0EMKysm1jhDapbhelVE4ZOvy
3rMjlKsEEu41r7Kle/xWI5lJ2lAYaQEI4K4/NUJsmnlElcHOsHgfZnSSS3JcGP8O4YS3SA7FgeLb
lXd122ooB5m7ge9uDwpsEXxdo294Lv9U3E0s6gP5NlOO29pZWq7JlenE0vh4LpwQMQ9KcE2jWQ3W
K9u7z3agu1C9T4jHffdjgIC1T3rtoiKqijU3/UslKPDlMaUngzBxdpRPHI3Fr3acOD7F/6eBTxkO
pKqLImSJIrNnhMvDZhPCwN4DaOVaW1d333Pq9mCS76rjlTmouGsbmA+7FGwWxzpmrZrAWcQvFUDE
Lhg0oAw+e9hepSh9YEmkVKUtQoPVxDrw0YQe7URMqsePQRkg+IfJmjpZyliJGTzOdjou9rytRSwE
rv+GATOMvwKRYFyTDivDXHgsjI93FNiasahPQLkCdK85Y3+4Od57hISpY5enMghAEP0N0qcvrsOk
1G/VIeaiIx1TZKJhTzpCTXpK6ADqb7AV5zbX5E9WKOsR2Np/d1vH9fNB9okbOJiMa9lB9yrevLFt
TwmPeDzmgeq9sm573ryiFk+QauekeSf7zZCpmK0zxRP8KI72buTOkwVXXaVdGYmxG75rRH2yRhNG
i+rgxL7XzLCepvMeTYtMBwVIyi9ezH2NX1MAzDvL695+mcrSxc5YTF6iEzHreStcb+GT8oasGL+s
LKY47vyhjAbL7Y2y88MfXf4ynT/dO5vx6Q2vttFYDbaiZTI5u/0OyjQcUPLzNusgehzio52mX3Wp
qUz1fI953dC9dVvtx0dMgLgE2YM1dQfK8tavXHXLIV5+K7ML5ZfUPKAke6sNoIDj8Q6JTU6YO3YG
kOutPpILBuj8Gh5O+ljl+UO8m7H5J71ypYy6W5o6fGfihPwjctz0Hw9OcBEiyFKeY9omForf0j0Y
btiVCgIne1SXyGkG3dlew+/Z4ptPBqfUD0gLnG0mGlDIyu0rLlXcziqV9VqEq9Etu3xibQRHhGUg
VGYZm8IlRo9/by8mFBwO8j59z4hloRtCY6adrgoTGhg1u6eCno6dDC+djK2P9GCURBb6VWhRj0lY
z9ugx/WH6HxbUynT9CVVmx9/WAE5FaCtsNj3rvfZ9JmWxRVkHjU90aPqhfpakxg/9HRruPjrYi9T
PVwEjSKMCQUcbpr+YDCioRD3rSwoH94wgXoLJi7jcjAkutqQ2mLX0JNxWl9+E8Loq1m+W5YFbRl6
es7/9eTTfYZ9pZBSa1EKOj6Nxk3L0W/2TkLNQ3/eAyOZfIkmW1mRxAkbINUSSD7G6Wm+/MVmWjfV
qaaT56vw3EhW9buNueExkObiM086jrEzYVnCUeg7tl22KSMlidPX36wd3OcVQEQV0fPTB/9Eu+Ti
ntbNado5dW0nW9OaQkh3SYerkLJTt+0cWoLtWunNks9l0Ls9cL9Vo8HiW20aD+KnR7po1ihRu0N9
J0SX6QKzzoX65ZDKPH2Y9owKj5wk1xx5029uyB2bjdU5kHgGix0XREAkyIChcIUlXXnNwvzySr/J
hxM2ml6HfVg6pxePfAukf0nvjg9Ik280qy2GwM9Zhw3j0/cqNq3IAStfKIvnp8f65pg9jb7VY9KO
UEXLHU7kvrAHubEtSwFzTyccF1ETcBr1zAqOANxLYFy9A0dWWjzN2PnUD+3fXMrzWQUGH3NJdsr5
CbSdkdqAvChakxMoH5M8ibHPZrPYnnkbFzvwsXPWNU9LuI6gbMyjnMsK5iNSqEWacun8kLiSIe9d
1viqN4PCXGI8MQgTcDAAKWN0VbLi9+rHgvS17vIGToim5zchBi4zWKOExbTkIqaHmAweTgM2hS/S
ZbEg082fPK5BddEn/xIhuB78FOgtiFyApb180kB9o7aIV2vjYD8ZBbvxr2hzBOZm29Z/XictHzP2
nXUQ4/kmf1yi2PDMPcTrCrwvGD0zs0m+6cPdgNibmN5N/un6upBYiqGanPoyvfHicFXZ8s+KUwVc
hT5Nt6roIIXs30a1xvEvvkJR0hwsMTD0ISsv7Wn69n0Xb8KIrcpSMD6gDtRH5Qp/NuvCpwyFYZsi
spnOTwUTkq80CF2IAjK5xG0p7iL5OyNvoeIshk1YQ+iJ4B03wptRzwPgveiZen3IrnWHUOS3UEEb
UN4ZfG2In6P/cM/UiEFRRVMAs/zsHcP760uYkS+v80QVNblmuQ73FMgbNq0Na5LyxUVhvMIkjYEt
pKwWwckA+sOtNU2M8L6YFHbHVR9iCFkaco0TGWGyAMkoEC1SOdfuL8+bY7Cj5PTfdWzeZQBwla9B
vQ27jezGYRPlDknLRq+SjFPC5dGrVlXzf2/fmMSUJ1z7wUoXojBllobWgP/0nATBUXWqtFOPGUTT
l4C7otrvfwvcEnktTDf5rK5X5dANanlrdJO3qru3bZ6JGXoI/zVQBivOSXItz3oErnVcA4U2b+z2
9o2Gvnt7t6VfkqJptuDbnI+IAva8Tsh96Y09OVcWLa0mQxd3poN6UI5Uivi+28/8IYvlmDCVtRaO
0AwG8eU1TK0yWGqa7VGhrsTL3t1BjFbcTMbNCFw2tLlVzT9OVoPGlOU/psrOb6q1Q9Sy2MUiecoM
VA7ibutHKbh+P4CHMtNF+MiaXiNvDXZ2HukiBpeiBQc0AxNLy9oNpFyBS8bacXHreBA+lWrriUXk
irTatqIIlYqZWjtrnolhGN+ttDBmtOk4fSRIQtmRimqnqtyWefKQYZEEjJHc9P/B3j4xgxKHDj4y
kcXaSSUb8k0MqlkEhitF8xXQb2TOq1zgWHn0OgjVEAVWyMnPAfw6oycXgUMjk7kPAaIikxdUztpy
VypFYBQSqlN2RVg79AS35VRrjhJQxNLaQX+/+g1hPgS9MwV8p1ufwiBjK442Nx7tVmXXH3iCmdXC
ejAwjdjIZcPw2nqmhAPpbcTTHlIZPMROKMv+inJezPpekqTX17j9AXuFncy0kkOVuU5MFWnN8vhq
Zdh/Tt9XXgP8DXOFnCI5hpvXM5KtBMsgN841gKK8IDx5ajH+jyNHDNlLqDnqNl7fJ/oLl97zKgMw
qCy9ZhNkDpHXzybn5BJY6uUyGlbnfxYlAjYQbu4YzsxkARN+2Ec2tVvN6EnXr5GL++tPJgDZt/eC
li5Bu72a4HUBYwOELquVGXq4PQMFao2V8g412xMK8wuFMxeQ0wvECQetXMvuQs82kqeDzOcmUq9+
pw2uit57eWoErQtA5MRcHaVW2RKPkcnnTmbSfT+gl34gg7ffIz4xFhEQmqCuEDvN+6e2kDvAHZOo
Ajgc78wTeTOTVsIcIUJEldeXlhWBM22sfsMTjDzPByc0EwNd6oOMykZVOy9dJ3M+97SXfu5t/iro
K3B7grnoLsl0NgM2hDK6wKaXd5zwm/S+Zg4ZCOCho/6dRH6+IDMGFhy2R34ogb+IbaJT33sBk3ey
e2pA6D6EW8rZyglWl5Ydo+OLMsSwXYObrW2VA658ie4UzSKYtjmVqMq201pDMELWtseZXf7v184r
lqfcHytI9mtxumr0i5MhEzNqGxaVauhtkYvddeBS0PQd0Asdw61cRF8JANHdNlycU8haNOrPwQ81
vl1iws/BP6S7yyYmQpj+omkIYPsdXtT8JuyJmVozXewGYBkeb+Y25fiD41+D1FdcP0T9bi/uu2Vp
CqLCzcdORIqQllgGzeVp0eYRebpX2spNhRTBsCl5UFLKIarI3cjelnct2/3uaeOIkfm6kdeRMJQ7
1imCI1CDWBtIPVwU/hEVTNcH4DaKYqKtvCr8xiQB+2GxdQJveQmSv2IJJs+Y7c2XbkUsj4tW2Obf
HD2G1E3vfC85xClu/f7K3XSqKkX6gNHvKiOYdgmIZHKi/GJF353De7eJRRL6aDq/EvuZ2TOYGbVo
2jTTQGDiPLJO9RIS9aMKz5fqWwRBgYwScq2M60Bww9AymrGd/uL2yMmJP+gaie5zxZPqFa4QPMXZ
pNwv4ioup0nMhWDXdylzMQ3p/WlkrJ9PjfvmT+kn2UPzylJBvPY85T4tFgKsltnNC19M19ORY31H
VI3+FTlT+B7RRduAuoV0D4n1vMsnpNfR1j9TICFfYgTylYc8Mq0L6ejpJKXyWGdHU+ysCOzc+xo0
Gl6yAWwrBKX81aW/zjfQI4c0Lu8K6aZqu8YCLkOgYJ29BiBZ4eswWQclvUX+JGmSFF/GDOmO3ELn
y0OHOd+hp44nY22rl0rWJ5xDuJguENIvv7xiftT7I6dUo/4zkHK5LK60oEsq8lL+2azNWUZbdLIG
0nZV3ZBcCJGxHmSrgwUXoY7A3JL0S2adKYAB1YEhLNsLCOzjv0fqcQbOhxAgqgny+BBmDlmrnXOH
upTExT/88UgMltP9rLnUl+bdQpaV8Pv7v3qj2MiMuIVb3r+BZBJBkaGL1K/kb7Eto+w7ZfQclk2e
EsYAcJBCrxHoKE/oOE1nKdwj4rXbnUX5fPb4GkzkAN9J7Age9FKddTLb0b67KykVoGNIyZM2vkp5
E3C/gEJnHt+y2p938HdY49JPVxp52OiSS02g9TrvfG67H/nMwE3TSljx/q+K/VCiw6b+p5S36cri
hAungAiw1gkzeXeuVqCljzjPmG80Vl4w40x/pyoKByhRBzbUZQui9V2cBcnRZKKUcm1jFm0gR+OO
eHq4+ZrYRpw7QgEXaUJOSEP4jKX1ptd/wvSf8Bz9hC3YvL6TL5xZSPEwtJlBoLOBk3WsqDP95V0I
DzKYz8R5tH4IgiigpvW9WyzD1WZZFSglCKSfU8Zr88csWcjC0HJlxzKZYJv0xEPugiHu1xTBtEz7
mg5hcQFyRNSDHW739VryVW6JcPoEx9orHDvTzePRB1SnhiY6v5FTykXrUWYDHAoFKyMCgrN+w6xm
5yeDmfGKH0kUogMe8wX0/ryeKmx6hE78gqQDbF9a5m95Sf1xt9lb9dwnikU/KBa4yoyZ3KGxYQjh
wxhtSqOM3lZi78jT0b/aO5Nz37HlX7ios9R9CZRUFswIrNRdb7WG0L4cMA0lZjxqJa15oEQeQLCj
Hjs/VIgWoXHisiBYqgXXtj/66AS9p1hGIxgfCF42UY7043ZdQjjZ1wC86F7cL1/UK1mm75kUlrjq
NKgWowtwnKDpEzZiaNMlu99w3FIhk4mq/IF8e/jCy3vIwF1q+uen9zAbA6y5/W4F1kaEe1Zt6+/G
+qD6wBD0nKLqX6RQ9x08Bxh7JdEHbXCA+xBg+m2HHOj3NNoZ5EZzZYcn8pra+dKPcA/h/EqF7jfu
luq7v4MIzMD1kPtNbcIXrLsoxzLI3vkMuIUjN0F8s+RVSRJTqrQgvV2umHUfR5mQGPRENqv6qnsd
xiIgQY8jd4Q+4zLwZICS3epylSYoHVCQ3LcANnuH+7eajfwdldig34ewHhmZT77xGHTRQ0CXs/cP
aEKN6PYJm124vDDadzS9+byBnbxcdhi0mHnbS+JAk8mmNnvrXOTPoNcoLoQ3/tt9Axc987HVEd3Z
b4y4cKgtlQRz5ELO/T+rV+LBgCVH0/+dhWbURWSBmn/mZ7pLEkBZ3zxI+Ncu/UvfLMwa68i026nK
7gG6wSvrZH00TU9vz2L6qqjQuc3UnYwhXzimCktR0Y9HiMcO+tgm92DYO3jYjtKd2HvfhETNdxq8
eteirbn3UOMtlW965s9tT6noMdLJwk7opaZmG5LfqFpNfzIxljr5RVU4c1VSmRNh+zccfQ7ac6X1
rfvF2MB4OkUNZT2zwPG3x8kMM9ry45w7sDiKpQ+3ZdZVEsJV9qTCYxOCiScWSbPc3xZeHsjZaA/M
nYodSM0SZOYybeOtRqIDYnxTZ45KuSEtygKxQiq+DOmRe91IimKeSiUitMlfecblvkDkFHRbeY6j
apOhK5Ggj7Wdo3rsTerUHVd+Kiwwt2CAWVd7F9fximK3t+F+QsGaLBNYatobirzG9dSy704MESkC
TYh2hhUtpIXhSACPzPreRpSaMufQ3hbamoFiOcO2xNJYslVwUJCbDWpvGpN4AMn3bHwTFePAFOX6
jzbrqkSL9VwevlF+Y5cvmgeL5vGMbRIMehHVn6R2k5yOjio8iMPb5DXrPaKnCpgHzZqUNtQJJF+t
vYAvmvFFT8rc7OaO3SXxOZJ3DJmhmjYBa4XNBcGyAHsnig060oy8bb+JGp6pnj19GZG1ceANC5mC
1JggH/SbZyS0k/HnaYX01VW1bti4jKuPxMnAwmK7hbCKzgb9fGUwwWzVhWm83OXwGKf+zZZ4DhvT
WuvUbuOVcG62la1L0E9cIAbjbjWfYNV83l5KkBB+WoBaDYlBaDM6C6AWCduJyjvUCCAfeboQhK0F
n2EJ+sbfyLRauKiNY2a60Pl3II79ggiEmKkzjUhRJYxgVvyI6eDma9Ux8JysS4tiXbTE0LUeZL2L
AzmvSOtw6YRApkuOGXMeoZtD5u+18xAUO7Z3/3qysHJ61A3SEEXQ32JITEJhB2kHPgBjcz+S1Hde
6+yzIg7HNCEGLOSH1RDjEYBBt7HEne7UxYgN2IZkQic2ooZaRCf+HvFdMiFDZNhmrREzNm58ypJT
+zyPXurIRlQQkzoY6dDermv4Xp7rbGkWl1cBJm2d8IpN2MsdvgAfwNzZ/7N63KPQOLgYqw2TCMoE
Ke4IbzqvAOrgQwuZt7L+GS+qD2aJB6oZj3kTtDzWn6IpCeSyjkW+1dMWMPsHfeXUFbfY6bf4+9on
GTkWnKHaqWI7lE4ZXfEGCyR92xjfvkTZlhXYHLK9wT8raBfAPRL2Sdo/RndiqFaxAF/gkNm5NcgV
Yhz22dDCySDfjnNoiMuFVMqq9mlhebrpu/zMFwecD35BkZzi+36AV+jUfb1FOvS3IRuvPF2Udb7M
ZLKg8+5XVNcf9hnxk/2sRjyeBkM/fmq5QOoKyiLdAkrfOepokJ/gR87Z3RNN9gDstHeq4pprbpqi
mSVJRsQ3LydsUUR4oNAa5LgjkNT7o/mamdDozM1KGJKtQvkrYa7bYP5U5193HKWq+ZAaOjo4aE53
JOgxFMGEyhdj3AgUte4CPu8c24Rqgivzl8LvzIG7O+xDVTrQuo67TK8BRfizi+6iZbazZOkjE1A7
dQPr4VjeM5lHuRpM31a63nV3a6dn/QOcFhxFukYxD5XitIa8tNJkpJz7Ghh1gLe1EO5hfo0zsfMD
74KnT0+NDWY+N9ammxIUieeay1U5BhG2dIRyNsIjwlKXNSTtI7t2zySuRTjn8GWInhikp3jdImQm
7EYUxI1WqxR3xfiAUzAd3Q+tQjZTRB0hUKozkTALxntoR0YLItawbMbdEtbU6viTsUMomHN0IzYW
MgpzRNLyYDrVOrFXOlQQRaAi3mHCxw3NeG7lz9jHxh00iKKKypRXx7lSrs8PvZH2H/USBsrC8XZs
CUTx/LzNBHsWMdL/KIP4MMT4pRPMEQfw1VU9+JEHDmYNvwTLx2mWqocrZa78DjjF6GVvF5qoGEya
Yv+ZfS+evl7lu2XkyOlWeFG5i76+Ql8g6foL23vQrJqpxTmoLTn2ca+9sBDZUsFddrUJrrCqKWFf
q9mFAoZsHCYZ6evwONEqXyzwnkGlpwXaIZUpkyK8Vs3UeH7prIRbuXpri4sC54Ws8e2vdb+YFWwu
STqFL+dRUooHKbgUo2buwt4dQh63INtXgZ+Qe+YDHnq1PnsUnNitT5BpF76Lw/VFsEz8R3SmXzUN
1/p+TmHIbm21d84Ru9TANpxLZdPHr+LuDbavL2E04e1Vx1XFUlrqW08kLfHIQr58GiqWJf6mYIeQ
Z/iqKw+el8vDk0WM/w/s8i0N86zcGCxR5NnsqXUKlnE92F9Zuac6rnXYs7QQXjoGvrvGvYBajiXo
nw856it2CqyZ29gOcFbzVJngH1fJU8bdSPeCP+KNkDud5pTecsrIdoQH73VEXBmPfuHY9+PmjnqW
S+X5dPyUyibv3MNplXFJ1vGRB0/ipx8d+EpdUbQptvOQSi1Z0XfG4KFL7pbWbYZqKdwd8UjPQCJe
QVfZiUCbXeasuKwy9rNCGU8ECXYgDCDEvsOuqRSZCffx1a9DnHYnk6aAaMFjTeCPvXwdXkDmAR+6
JCUZ4EOj/RV61eLePzpQ1Q4vVY5IlUbBxLxmglMOPa9KZmyQ1eUoodVa/hLeDOufuf5dXJ9sYKH1
ilxNXM44xTKrMnJUWhFoAqCEJMO21jUGnOAcJu1h75O0wGZOqjsGPUtWQxVgM0ra9K1nBZU8kmH1
bPqCZgP0mjh/UY8QBMX8gW+S69M46SU8lCLNJjA3baa4z6XdR4xQ4SUUGI6Hnhmqm5a0zqtrWmAB
8AdR+1efp0kEhn1gDkwVphmNFF2Rb2/q6DM+xFnu7CTVGXwFoKKxZ6KOgDTIqBLnAGeiS4sEpU6p
ZizOP9KrikrLTQagELmH95F3+u0tHSow7UIZXLfx2Qv/qTkSIwiLmG/8tIkt2SonQAhqtvh+9Qwo
Ym9nWGy68qS3OCIwgcPsdYUjaHBrhjBOHHPLBEqpLXvr205GprJUAyiqwB217q06QJEJFQxBQiKa
41FOe4DtKejwsvU+vh9TRZ2tCtj9ZUXEqAqlNclCRuDBY3i1TXDgVYR55JE3NsxcQDmM+Fv/Dvz6
IOCRi5UrTZVgGCjx+taZNUQH8EjKKXUW6EZxwN4ExmMvBBsok6t7ULLUGRfxtdPm4O1/T5jEHcUg
BrRr7xd35l3/xR9kegWt6ShecV7JPtGTEuuGurf0aWIO44Ou8daVLjTaSgENTDBqu1A0MpZfF96/
oCMg+n0+cDpOJG/vQno6ZLluJSo1WfaaIgwZdOf1DCeGa2YqkLykVAmBzeYjI4fNgZR2pONihEOE
jgLAqjresnYqxiRyDmUrW56ePO0FcGzhgSMRP1RqpU+bTOVjUCzxYXBaAkadnQNIvNwGfKdqCI15
hDek2khzff3KHn2F3sUvdrK6kB9hnajrr7quFJxoylWmz+HR1NDk3B0zJhCv0CF+OBacDsq1PuZl
0N8tdy+4gfLkSO7qjiH/rqR1P60zHwJqflHTCI87Bys1f5Qa0Nv3T74kacz/gPitQ2caCutV2zXL
dbxeRD5KqeM0Ql8r3wYBc9s2vsbs6kX2jVybKMut6wjR+xSYXuOxEslq3I/TdzlqaADO6kf1GmQ+
sPPtLao382u6Fpwm4XRhN4jBQY+/M/i0Mp9e+YCOQzG/MpJiWYUtxnddQpmG2Du4jB/rNDrL9dLM
WSW+8pxyRsSZwm+HU9ydsz6jL3W70AYx9ywvhUrMqGmGZDXSH+qNDVz4scgX0yT+0b06G13+Q595
jy5ONu0jlISML37yL6YwaQIx1048G9b84cp4Fo5dZkAG7WhMHyqCO5DosVXbYNBqBI6e07tWrsp0
jhLspgRCgrH5eBErVXeFDyfOh/Mypd4dVIL+ESkCKnQS64TEipqfI6ekbSqOviFhCuLvvGW1Ecet
XGGVjM/Cz9aMZ4TMci/jCb0l+tKK8AeUdki5LFoxDtDzc2wxW5MdFprDCUIYI4Ac4JwdyyIspqk3
Iiv0kcKfZ+oUwdS/T6s3uCcBLPPzNrzdFTahnLZFnCvfPFTLL6qXfTfRLAsfUyIBCfE/WhzThmWj
t0alAyfc3uI+WEjGrRPZVbfD1rBGxCGZ68U/aUsx3lh8d8Q7mvKRlD9owWqzOASgUso2gzwqPSnN
g2avVLPsJt/+2piEksz0EWLv6JY1iuzGJBWaNy+0na1e1ybNw4PC5u7DIZUxnscCd3ZSy9qJwYOM
C/GMIDAy7a8jCBxIZR8ZxmR701+WOaLVkHAU3hdqGZs5o+m5vWP2ePMirtWu0KBdw/NAYhaaU1BC
daDoigFoe2EJazN4ICh0BD+tmxyYJv1/TXsKf5UhwjhLed70Tke/zwdQVL4hKYfHduR6NoK9RUgi
4YMQSxDc10DezRdrdHuGt2z6Oxi0y+tud4yxX0TpwwgvzZfRSU8nDFD5CY9KLgYYpELun3btDl2r
NvuPSIR8SHx1AZ80k4SzxUoDduy96rB00WEC3y0baXAwddrrRlYBGjvCZEtJdU9OJwVjdeldHOTR
PdyNF4iQnHgMw6SOPjVtuR+GfzG4oh8gE4q4vD4GyPLXpFY8EmSqpOkhWVqVDt89c0/EGHNrAjWQ
hzQmbapx81vFPNTR+K+s7HIFGfN+46RjU0+axiRdVUtj90TL/tSwv5aig4eqtzSAOclt2JDqx3iJ
y2iVVAcXTkRjUziGX+69WAxIvC1jt0PmsmF99YI8PyGJSD4D02+UnqlCtvSgFo9WqI78iQWX0raz
aDnoac7WSV27N3tbg0virstxpD7Dj+i6juLzcP891msf6BFrUFM/du1yPh6TBYtJoAr7hIkjahEX
lqKZyA6CA2K6hk2YNRRP53Nb+uy8B3800vaG2GlE3K9KXIw5lF8fkYPj2KeFwg77npAJSpmwXqQY
7tI7wUwLxJkqjd0yG/mOhUWNzzl/NOoroPS6OZYmjZvwE8yQVMPBDUJwb1J+4mqLJSuwklYRLdX0
znrVLsWdUj/IrqL2PCkAhW1bQIegHGQDG8MlEKJtImMGtwzhudXKSHW4k4AbO7q1wvASKjQ6Ta45
u5Xf4fQs5i/9IihtuHTx6ocNP0oSIOevGdw0fgHP7YxN4+pUh3DQyaHC1jMDTRSUAUmM02jS148v
SIT3qrJtQQ6kBBkJHtiU7NtpAoUr7Cz/YCr/J26K+SGgjpIAyGQtfk4QH7f4bEOQnnFCVKdO5yWp
vW2oRZ45Mjpp6hYEplpDxytcdgTMiFsqFdemTDSg08IYhTzzgjkob2BNkRNobQHF3rrV4NHvhX3Y
JZR1Nq8A9eVoBof7M/PsVXxDncUKOn6UlInrHe9GuuD5/uubB0G9+fe9jQXAGURgN8KE/zyS8Sln
E97/c6NQHFcGH8oS9abS/colzHUDMdO+MwsiVdN1AmShwldO4Oc1qRkr9PrpoK3JeLeFju9BOh6b
JdBFgZSINNanROZ8evsaDW8TajHf665jrgnG6DNy5ysI1asA8F9ZmKLSkW9Ix8m+tXTYZTRYpAc3
RX7M2MH8lVomM1z7f0k7dbHo/Ma1Sis6uRBMMd2XZl6oZe0UHG5b5+28DAP6653gwzPoKA7jIx0v
Wl8ZVdVU7Fn5T97Jv8gQiTKYH3LLP+BxGqOjLkWwRim0VN8jJPz9O0nmwSgW7Pq3CUd++regGHgn
3uY1SofAn6baD9rSFa5WjjplnDJpMTHR4VXtE1OvQa+3qIhp8ehK2E84Fn+/JerXMzA8POHXp7Jm
BVxWMe/0/F9If32r2JFgvkHwUAqZYPoFxqLjJxpfXXjYJNQ02HaZp97SkZQN/2w3fWGT9nyO8u0O
7nI2zx+sXSStUeIurRikWU9umwgKL6GAf9Fzo9AgK5dYb+DjSGcoQsiJdYzvEDMEgpD6fNj3O/Iu
09WAVmI04aja+0TjQN590AjB4rokoPCzOctn5TIuOKhk1FFEsoL1d50tNcCNuSwzSO0aMuKI+TE3
m8M9ldgMzCskl0mRpMlo1JC/cIz5nocQJMLldGZoQ8t4n3JSs5t3zqjWy6UGyywaOa7Vpfzwt2F7
O7oBKDdSLG1V0SRoxpsKRSJyJVTsGteBPnbDGhkWySEduqGgS9xjFJUvHUVAr81xgGIqNAFSVW/B
mG9/pz1eYen/R6W/7Qrbmgt6RcyREgpF8wWHuf8KGOKYmjsbGcUjXMj8GyavAqbll8VS8CuYqsjh
7cwxIK+JXBlorYuyLsSB8GhCcGFp9kuZrSqhzNwuoYNE2bKEb0Jynm5HN78nweflQOUSPzU8OxVB
qncXIhZ4Kcz1CxZR6GenaPzcOnEP7UcOOp9oMLaGhEwkFmQtaOG7+Gl9iUmHgAdWgANSDFiWENcm
yUnggDNnC2VF/0m8p3xmFjravFvANfURUNOINtJx8Z1KNkPEGIF+G7z00fLyxpVulaPfGmOnMfZK
1wBJfx693fEjJziUBZySMeXwK3lDkVC8KsP6QiLBuc8OGL7BBOs7DmEJaUVDx4qqxuwW0NvS033L
X8Hz6S3ntHOg/h8W5QY3xVQyaS7lG2E91gc3jIS7qgEy0v/c+jBpdVgQAXZF0T80h2Q16gXSbXE9
JE7xfQjV30V8V0bg2OFt6hTieIbG+nkceCdwnZ4be85rW6+9ElVTpVWvRgwFaUuFvEhjLLtUvUzA
fL+iZw072P2fDxlu7t78VqxundifzGe5ZPlAsV0Vo39MH13baeiS81GlI04FYdYBj/kzPqRVJPRF
VNWcur8MyFmjGuk8FNGw5gaviUS+tu/ctfb3mgiNPmP1I93haLj4CvcC8a1uCcahMSnJET/xLAa9
HEATwxXjNQI2lGXCxanOnjGwesbrsGP+PajwAzr7ImPR3pp2ndliYlKqSyGqVHNVjKrPAeALNxWX
HAPXO0rRjAJLs8sT6cbrnJcjXJXTyTI8SzmKdgTLexstq4a8fdVE4f3fhra0gR97wGZFR62QnrWQ
7+M/H3S2B7dCoH6nuI3+5yZeaFkfM9CRJMdIlyQG3RAQ8pwKQdoBqtknNlb6k6CSHtewNtoytpre
gPvNiB/ag9oiFjuAra/aNqie33bKikp5/6lNpbY0oEt0F2SGMCTIrQvV0JqNjUCeE6NbT2B4Z+0F
9RIUxrCHVD69Sptdr7aq5K+bsRInanb7BhNK/IxyrJX8ZVbX1wm3MXeAQwlw5qweb0DHUwfMpMi9
mXiJ8tkHb23pG8ajKOt97fILIz3e2a+vBcr/uuMp+2pJyj6V2cSiEKk2YRVWFQ2+shH2baAmdwlZ
qffhFAbTHx95GHanMzI/j/JlLeO6T4vkq3ehIuRphhLfK5ek4RCzT0ufKnazWZ8unmMCD97halW1
vxZiSdxBjBvZbhx5zZXJxT1m5Aim3T0xVovVapnQR4sF3/e6r8IL/9IiwbP9Mi2NFqwVHi6ctISx
c83pyXv7M+w+sB1RFmfvEZVLmoMIlR5ttt9LgPuL3bOCbhSoLDTI73EKRwQOGnkyWAT/myfDGDOu
vftRDkMfqQy2YHMmFTNli6mEGjMGOYuzb+EP+TQPdvW7ra72IkRsILVczHaGaS2ZCPezqhQMEikC
QbxUB87aZYsd3Jc13gD85djML1XWyo7/U7RsYauc+Bk1adqBTjxWiUC+NOkU2vVmwONJFwvMZNhW
WacaZBfSeaaFSWnxX+uYzmmHA7BZNAULoICt52gNFnFj141WJvF+XaMCNzK+nWgOW0lkGAZddXBi
oHQ7MSbDNqE+nMFIH6EXb5Ntw18SvV0yiT1DSS8Sub7Fu5ZKhy6Jyg20x0kU5q2lOtRTs5P0BX8g
psy+lHTDnav6SJHc/rHPrB1OK5qZx+wneiNKpfLY2u1Oqlt/5pd6tgTFbzbiZZGVTSpt4tRHktAL
i34dvyO0Ri4DBGqVqgkCJPOp5yGaeKL/7hBHkfQ5fkxranqJ+SyJUYT9xJVUe7CehoevbktjN10r
nmyO5y0Am+UhAImmTKdjuQDybemWlIy3ouYrS/OerXjCFOIVjUzzG+73UI2M326Xf8V9JkNaurdc
3Q62SfSK7RiA7wCksWM5/G+8SlH6gHom/GlvO8X4jMRrh0DpeoBkycW1lHCjWxxrBvHD1i9Z/MRA
YSG1KLRkFSZP8slgvGcE0Y9/2C9MzPBgT0YzY437824/UWKJrMZGR7vQNGXMK/PKlfj8I27EiX+2
kwRqKVbKyTssLUbgclJNRTCs2Dz0fRv64SbZTbpFi8oDlwhzkKQ7AS6Bg63IBi9162xbj+xWJcfk
OA9RbyKFbZzCK4S0poR4ZNUZkDlhhAcVREMzv92gANIFy94seJbOPqWpfFSgnjdmw2eGq7CDmSio
0OCtJYYVq08+PpTgWWeM1pOMiKuata+9OhCsNss30lzVM/BWnGpmcTb77xtA7zmbSMH+9hjliVvb
gEavEirerXoh5caCLL6j+Er0lzDW9JZNk60Xluyibo6ccud+HQ8y9Pp2H937fi+jNTpBJxse0OkG
Gi8hxB+Tpx607Yq4H1kq9gKL92K3o+8zVzuZW2eciRN7k8okj+Zk40wgc9qeuZSelUfM2ymgamNN
yyNrWtV1x3ybGxp6FGuvdXSgEOylamzkuZYKeKSkgWQcK37AM8AStsyMG5frEYgVWxx2rE71loOY
0HhA57hbfKWLud99zr8kUPvTpMVXzB1wHu7UHQDJ8tGalt2MHpJGfyrWbARlNb6x4qNOkaYuV5rN
N613q3DT134+4xc5Bg0efzusfww6yTmbqiXhIHMfKdktlaQpiyRQAIx1EAtM6cLf5D4CWkomNHgh
RqQLOUzOEWSOM+I3Ghkv9JlUPcmKzUpcDVH3G9vrzLB5H4xmRgpfAipV36xH5rNzAy2V4eCflTse
wtgq6kNauZRJo5dTP6LkMcBmgZOnyT0LiXoqruhbr7Rz9Mb96o1VPLeKjPFOG4syEP2ZNYS/Fsrf
MVS/5bFlxQRUpZ8qPEG1fvji5SknhXHliauD+AbUQ9TiogFUwEgBDgyjEbOW2rMreEi77wbZdtZ6
Suub7m3HCSxiRCwj1p2X8r2qAfG89cGDkFziZZgb3eQhnA9S+YQG9N0lUHiweTlhOAPrAG8cbLcj
f6foITMADfybBL7oUbMj5GCLjfYm0HyVdZ201KBghqmvAB4c8tegQYB/7+5anjrupWhOLMrEsvf0
fSpJxqEYWeh4dYRTt1gRYH+jd8AEwg8c/eMl5TG2GqK/fc/9a+SycgPwO8QaSTlDxgoyHPvm9EC3
fmrt0wAtM8Zd0L83Ea8jtGZt8WcY5XxqYvFE+I6zsQ5Dtd/Nd6ANFL7zwlJNr7POKKftxKWpokv2
YyvbffUXCVRX9nZkTVvJsLHlgquycon5IAj00nP57j4y8pIoT4ia1KXp82C/h6f1g7tbkD+AqnHa
Ykq6cny9vKAjOLb+cZbexqKQNk63v3wT8YVsQotGsG9ke1eObvKui33G0PD0qMHF93K9ujF9h5yL
u+vimJGlAmbKxNavELz2cZ9jKuZbK01khaCLxxCD3JCKhUjvZ/F/XJM9o6t+87kNLQ6h2NgNxNeN
UbUQa6OqW35KyqkPyDEumjli2IIfV0G5bltpuSIPFM6GOAPgOEqQ7axWilfabkW8P3jkh+BY+iDK
sPI0i7dsdgJf9M4khZRvhdqkAEqYpqsX0jAm+2sW5hCxY5AWAUoH0Mejp5QbetG8tCTrvXDJGDD0
N84mv6d7M0BIWRKkAnE+DWl6a9bWhJ+9vckVn6jJP2rZXT2RlP1pq1CWuARwmCqsx59XJxf9ZZJS
F8M+sD5nJF32BHD8l/blswn5N1Q4XGTdWWRcmX3slV2S0DLltcv+UtyRLZOoLpCgmYB6RHYe3hPF
7dlEsAb/Pdp27nhy6QeViiAM2z5gzKl0ZwDBZoai+eu81+WEySfGRRTf+NBH67dXVG9NSNWoQ1FD
Jef9a4WbfChHQFu+lqyuKbGjakUr4+5FaB33LMtjIXvSmEVBcaUDS/m2JuwK5tFOXhxLGBdo7piN
2P9k4XLoCnFe4VzDZqu7din22LYTpXgDDc7iQbR1nIZLppW+KHDOg4vbv19QRJqasGAT6gNOJO12
CtgV5dAWThRnRqeF7/e2LrflnpMMKdm7D8kq+h35jNj1hkgZzVtaEfSKoqMK56kJIrbncKabJg5z
qFJs3vOJHM3bnTzzXFCEfcyPyE1fhR42UId0ryGzPsQAVwt3+L95dYi2BKfxjNTDHKREhl3LQl7/
OALFTqJTUY6cwuiO8A6X+c9taE1OMH/67wXqf2YexZvxfd9atwpshtnIOKu7MGPBFZxX8dkTt2E9
hE1dKvmhoVAulhx7J28XSUBZ0aIy9c2cjd3iw9yQ6Wq/OWbMp12wH35k9zEQkAJuBYLcpRo0ETSY
k/OlPd4BHv7eE8P2/BJEdEyuRo5+Dpvha2qmCVuoUHKeFcMXasbbvdfOKPVCWCA/hQNJQU7y26KK
QdlWtG7hN42ba2s4MLiFsfTzjr2uAou3Bj9yKkH05gxeVVZAFqX7gqf3u737WIuCDrzXiO8Dg6Y5
cFHvHs/YtvLzPq59BHI6OStXam91KLbFjwcAm80MdlaiSlm/OqfeSF3igaIcffvzbtBdTf6tamVp
xpsHvSYdlrD/4XSKZ6GM9f3VNYiEKCA7HyZxN6Bj+78vWu0n4MjlSwwwJsL20/mMS7gjPuG8XG6x
t+VdovvHyDw2Csy7olh6Z9MZ5HEBYN2YB+9KSgxl0jRm/TCJ9bZFoJcCozQDQ40a1xqteut9+gZE
25Gur+fXbHroQEQ1CYDw/rjAalhsXAEfjQrBcjPhftXKOJq5ctqx/JrDsh6vdcioFyRpBKK0TXDd
zPoaIUbaw6CNr4BYPdkawhPk6HulvUIFbim+yaEyxuz1dJSDrc2ng9wZezacLi6tTpO5bRka+GZ0
sk8HVh+w0JmQC/kJhPYaftEUgDDLIwwlr5tvRcjNHHgROsRjohKNEeehfgJSaShugJeyYE0hM/PL
E3vmzjMQNi18sh1EB4Eweo7Ua619Qm7AJJ4P9/Xxm0+jJLnmNXFcQCluBVmOsZ5LjyvxOiT3vorh
zF5qAwpifOVDgm2TpzZn0P3LzSlkFFPHu7QtxDAJ4tgdH4eclA9Jez+Fd6MX4kf1bUJatUnPRUgm
uN75NdumTMXOzwvQkocL7mjwjONS0sDm8u776+ESuTNAvl5dgoLgRHkSaNtvidMqnTK/fZMX1T6g
Rfj5lASf3fgdGYF2WC0fia9hyWz1yau715COyjvl/1BRRruaMhl1r3Ekewhi4wbYlzTM0FuHCs+K
XGovaO4853rxDQrpNDrv7netMpGAjwFkKW1LgdO6EXw6/H6HxGrfeskxDYSt0D7eDQMoCPbIfrwX
ToaJg8WP2JlWhDISZ8iec2o6DIfm4y731lojF+YYyFhqKdSXSr1RvYajsegeVyMh62Y77iYZKodP
Z279pjmEpEUXdgpshuVpJ4F4/Mmg1c3/kt4+OiBlTv9pyjHpksyaC9C2++2Cocli64+xmds7spe6
P6UIu5bdCB/iPvg6huqGMv6S3qUYfzmlB7rfjCn8Gx8yCqcRmkX9JdS7EneCbd9L047sU41iLKiR
d7bY5tGHIrdBoQ/N56/Z3t5UdPtsaAB94g9kyL0ye486KMGEpiD2WgLq0i1Hy42wkJj5w+/ursHK
rgeWwRXktuxZPNVABpqsE2PpoF7x6yZGN1c2AKza/71aqU5cIqDX+QSMTn9jy15W/AQ3hUnwPJ0Q
DIuFyttReseZdVwZ7pdxc/8qZCwSc2kM83nLy4jM4Way3LFOdjArjZzM5/ZfaC6fxrSdC3LXoQ91
7vsqU3fIDK5Y6R6l4F1WH97NEUbfH0xURLFW6yDowT64XPTwzmjE9aXzSHXR/iDYjY4uKn1HKYvx
ShuoBIWPYTD66+dDOJ8XltiLJBNzMD7wyzlMSBP/UroszXHDzc5V7qM/oUTH49TjF0vMy1OeR6Is
1T9kXFikhIJNS6TR4ik/+e5DUObZWqMBm3CXnIFggAMKa75FoSfSKZG7e/RO39KrDzTs42sLjFoE
aVnpxhljEcfoePL2nEKLEZGDjXBruMBjUwYgi5p5Mjpk951vtIlgVEnxXaqPBsqrrwsdNXSMBzrE
wDjpykQEUdssjZQatOmOUOy9s2HWYu+o+QtgEe7GVSJvqpK/ibaV8D/YWNVIiXi4nUk8CydmgqHZ
AOy4PFZ/vJcEHviQIq3iTkkcKVf18FWXn3w0uIpLDZ8TavidDBuiZ4YTcwe8I53acvTjQYyb2J/t
z3avI2EWDA0+4S2ccTPOtxl5DRBj4b5yeXdN75E5bui9BeTSoEneuv/w9JmafvJUOP+EInXTSjy3
0lsynNR4L78N6x7xf5uOAQONSa6TznXqWPf1yRT7C9BaX1yhJP6qZ3ob/t7pyZjCDW/50hZ3kJi+
GYdfgLBaB596EBwCGsojr3+I5uPM6uyUNnTt21KhwIW3HSNsTrUtJM6ukvGsWvi8KUxy/tiGw2Bj
oKcdtbFbcSi3eMqrfB51ivLXoPzw9YdIv+AGAY4TcZwFES1nnhoAJUPrYsv0llDKYXsTnFeoU2Tu
sRmb1O+BLA9vJaQYxsA+CsbXRZOTqMcnB9xyTgjth2GzewcACT4Me5A30Yc7a4WVCECn/gfdxYBj
t+eKtR1BDvrm7ikPM9zWopVppLVS+4iXE/7xILtGxrI9AUKhHoZBzB/D5zxZxYvojNeXCRGWvtkO
6c7IcynWk87FeggeKj0BGaxIIL9M5mPJdJmY1F1GjgOODgzyxQCkh3icPbnZUPwJfRbrWTRdtU0/
8KkWLci0yS3rtB4kuJR2cKBnZp9keJbkBx1kVGR8ZmX2XhHUzqO5HOd5qlpCnY3LdfMdUwavLvm1
gAwN6h2dDLJWV89qrpacx0Row70QJMfouEzFQ+jeNuB6Jko/fUxg7++yK1qypvB62GcsFwzRf1RO
dJ1cqf1fo3krW3aDsK9ARjcj6ZGwe5s12+7JjL5QP/n2zV7QtCtp64SsQw85MibNrEFJsse5QNwe
vS1K8biw5GwjTMJ9ffIgQin7xQ83M/hUvQk4MO74FypnD79/1wNMTfdRQuYUGPopOyRKRYaXLhqG
/Le2l9/0whlQl65wFM3f3mfA11C6wsNlAFfuE95aONhZr6hOvhjJEHj3cOkgyc6HChHS2xxSOJK7
EiPOYy4rPiBcqsavGOoJKjV1ya1hEHvb+bo59c/23rYxNxEluGsfAtSHUDy4X6bcwY4u1nHUkq4o
BT5jAr4PGhKgQLATt+Hl+4yvASiI0PKmbdoHxYrWpPqhLfPpO8gHW/mSiAKhvmRp0uVwzJYrn0tV
WOyvNhsIKN0rvHBk3ZTzbaLC6MY7MQrkr6EDVjMb0X1H+ImGXCUj5pc0SZv5VbUcCf7rQp92DP1e
6g+Sa5xWuyLh+VfayiIyGBtzYcaIYiSm509Qu64yKtaNGS3/0WnIAzowTzq3pq6YQsmfiGU48JMQ
7qmdC/2M54dam+puEjyLJ/x7q87P5mifhLn6f1T04O9KMffIDQ6hBqwj4CLDUY9ANBrQm/vpnW4e
ENntHrAS/FcoYMRAJInblCSVNr3vNRVCC8AWDJE45kRUnmDZetTMucHG1DC8t0jgX5G6CWM2gNwJ
EdMpbfUCyBWLLTsqHtADM8rgm0kzZXesg9VBdVYCGuNPJAKifMoy9RNQSTkWvn1mVawAQosjXvxq
L7Av0xG1kjuu4F6T7+4UNnHlTDWMjoKbPqsgNqG6Hn7Kq5SCCGxPCgyD4NQraEOaG7FGc1uaDMtl
IkHmOJOrvItTB77F3KjSbJhmWmgGWpMkYCHYbbGbjNznpmr9Bj4xKtTnAm3NyMZJ2eK6w5ZYKxhx
fIUsjVnGT/DqWpb/tI8xmiwaZhyr0f8DMvf5tLHbWnAChw3z5pUrHPx+Sb3pfbfNVlwC8hiKx7Jh
9jeTNHXm9arn/8n3QRos5R/yoUS3fiskhQeY60ipnUbGjTccGuqw7/PYu0oA9m+zmwO+kE9EfTcR
PPmzyNnXdjLED+aiDcClFcFQR98FLSf6JT8eenf9FjTZA8Nl1qyvlhfYosbSQmuzF/ikFOrvwPB3
hLDryW8fvbsdTGIZwyFTeTyteyp0W46TxB6DAuc1wU4VcRkifhJCYxbyZDxWDxXS47v8VOHhtwvG
HAuKT5AiOWV19nti3Pfpm3iJrRZDxoTnYEd+EAE7xVvVNNQ5PtskbEIDUf9tL3Ih6jr3nPc7syab
FN0C0bMVFtMRdX8uVq7ydg5jhoSUpZGu83qfWck0KtLrKoG3WaLPZRSgeLyE0FMKLZyROy2azX6R
WcxZU7+HS3Wsme1KbwB6Pm9BJv1qEEovL02rJkQedWpQNNVQLDFKivOTm/LSrhvLhm3vqn25ZOg/
43pKPLg5HO9kMa4YnaVI+PTIuggXLEe/h4WlEwG+kXb8djRGXcBzskOyXoQFv+9fcg1ajNbZ9CTP
APHxZgV5rpo/IfgVqew5+/SYg5D3LL9Z25bxo82z/B7exAOFdeL59VKxi8Bqr2fgYTdP4TZJz1fW
tLa2X337SXQDUKPwMGeTEaRq6tARwg/ciShtOl1psDFVdlHWVVpCijR9HVKx1fJ6C5QiHcsKjHVT
4jONArqzsv/S5uXgx0l8M8tIRONy+yE0Gdz67/eiCdPoNkY1VN2G4XyICnWU31zABq9rhlG2Dq1T
ui50ja/d5ASJbw+MsVo9e9NcfRYRJKTorVnqUIOBTD+XCs2ghV0wdI2vIUnFItOiVzrbmplv3VWO
EJ+8avBHDG5UyfbxY8fcj99VxTRrVqkftyqSMEmwQtWkCS+5o2m9TnHPitmvVnDPW/lrkRjodjLb
kj7q/xzDzUrdr+7/+79w/upLN9oyJ9hU7OtDR7v+xi+eO2LP7cMGgxpVmMs1fxt1/lCrdqnFl9wO
Bq+A3sQxZS99Hb6l6DjU5kGt0uO+QUz5/IWNVnLcH9ZKNmGi1/icROg+130DjfEr6zY68TaRLq9Y
iByLYGGZsw0wEyHESV6V/bvG8aTzwmpdPOJIR950JKIfqPpWiCLbJlZ7j3MZ/dcvd+3A3P+XAF9+
Hs9jp44w6T3oPJqpGsI+zIY9jFpY7rK2pY9GQlbr2c+iBYU6VDO5Y6DSygTa3QMv9JuirfuocNlo
9q/PXgV6hthofDkbbRlGKGqZPU1EFNaTmlBM/YcxuHsA09NCE3P3Gn2zc7Jr/EcYmiWcEovQwygY
UsWQrN0yh9hJqzR9IAeVj9hsDjVLTWWSAoWPHnybE3vsGhH0rbtfwzbzLPLuNOHJiP3DHXVduO6u
bayiP+j7TWp84FpwmnwbywTyw09rnmfUS89b4mQeUbzCTXtyOMrlCZUtxXKuXF5ND1RkDyXwZsls
gIx394/cn3wHqP2EN+A5O8AXurkXXfDOY3pIrFvKcjzjrPZ0CqUgDcmIwnfCAauAWzxLV4GhwuVE
Lgl/Ag7cwWeutwJ97gf5Q7f8doIxVnGJZpzA7bQqbX/woifDOPikE6pNtgR5f0xxhnI6ekXPvlRm
d6TGvXcKOdUWhTooi37v2uPO1owsWsPURhslZuYk42Fa3WqwEurdQyHHYX3HwzNIy0lbZQaz4720
t4wOQAQCPfzzjsO4jzORXnBRBtma63cO5a4p8p2nVV1Darfp7P++dbO2QsgCRyO0cci/U60YAhBk
5NaY7V90rTz6IaIVjLUDrfCBjTo0Vp8o/6a/HGUoIf5L6sMXKNYOdclL74KFCnXkKUz7XhvhmWfb
VukO2c6f6J/9tNNrIjYNfPVcTdAIx+9vCDd61yaaSQ+GO0DVpqTT+ptpS3FnP3OjAK0ZwPyocJKH
ntYqv0YBO+A6kFrCcKdgv55X9/8Va2JS+kI0wQ6137GXx5GyiAyFhdVj9aQR5XTJYWlGrhydzIcf
0x02xtrkWEYvkTo9UzC+iCniaI/inIPAB1pLcwJGzrKR1DMCetkG3TONHiPRQGGeVVgRzrXtCYqS
Ncj1AmVhgaBwXkBj/tpzuLSOL0WTHoV115wAcywTRScNjw05YO156hgsXq02r+I+KO28+w6Gav1v
P+SOSJUvIrDEsFhpM3pTpuYVd3C/goS72521sbBNvomKVsGyHPC4fM/X9NjWXktHQC2LL2ygGBeg
fa5kVptrQbEtdGG2wHVvcA9GrVqH4Ym0mopNff/T+mFPmH+97nxVrqoof0ljLtXKCL6fUaD9OqHq
F3mp4eNuKg6lAOHuYv3Oy0aLHFyCS4Do055KVgDQYgB93OwLKmgtkqFt0x9HQuRmzQ7T5LTA4Rap
ZkXEYOvsuAOnR0skBq9D4qdbDbtIFpxrPxyr2XvaNG9WYcbcMSm9ZY23csKmX+ewCbbgOp9U2xCv
wNAOvTNuLhxCtvKsG+kzVQRpOH0veDDsjPI3u8FsfQjIPM1v6jgmA6FYua9YpZvx0YC0CKMaDU3e
65eNVi6+8CbEiHeG3NsIP4SuPr/lcfCo+2QihLL6XLnVbvE1lzRS2YIK6NOOTT8Spe6NYCZCs0wY
+Rqdxd6xM7k16xkoQbnXTwhobULJzJbBiHDydSrRV7qSHH2MYIBS1gB4ghSxj6fNKMQOjh03PEOj
ubFSqn72N70391KfYHNwkJyghiPOmBDAcGtkoqbhoRB5HiJUh+DlSji8ayk3ZTM5oaFY4580aZab
jSKlrXNpblibcOBAuiPIuhhsBW5lZr8q5Sgback3El4Fm2H3bwOG+F08KnE3qSG5xiChii9QQaIr
Xx5HDQ0qfgBx/1E13coc/JYFWOb62rvawMEDdVkjk6OVra3vY6QWjRB4BuDqefvtIGoKDfj4tGPO
PC8SqJOhImAKmrMmhqzM6sQj8kJWCp16eislgopjnjISO1bjjy13x03AMXBX4hm7YIpnLiOBV/GS
JJ8N/bs+YzVgXA0vIr9XWYfJxbzt6jm6jcQqqEaVRSfmHm1vsonYX8ZCPY6AyPy5NGQId1H+jPHy
78FRehOUMDlFGbRLZ0bByeC3Bsh0TWbJn5rSBYnW5nvBHKtQUdyRVJ/9uPNtkWjlpDtL84YFpiK3
WhexH6wOc5Vk5Us1ycvUgQs2VUyeAEkQCapDEqJiHiXavoNE7xlaJiHJiOhGI9zWHl/pAxszOHUr
azy+ZzJXtYalGIYjeOUjHw8YUjMw489oqMXWNDt5wh9fwsOe5+33fBLKvvbncnWbQK5C7mAIeMqy
M9hGInaUdikFcs3ggQqPk88OXmUg1qPlScBrSMmf08Zvb4Ce1cXo2HaeuJAD/uLCV7jYfIaQUO8G
KKC5XFnSEw+rsk4XAmKvsfgwmdGSi+mvv+wZaTSYu3nNlRnFRPvgeJGVu9dXsI2Rbgsal7yYXmr4
imBqAyRL2euI6zA0UTcTYaldRQIvS07X+9rhxQrPDxsj/1uRIxfiMn1npm0w/7Jc0vAIQWGX/6Ht
LdvYfIxogBrl4h+swPNuDU78W0j/8tOD3VVSnjxHENco+Ji5uOueTtk7cB6p0/qhbO8tq/A+jAPy
RWhWwLjDvHxTWGBm0YOk2/WWxgqR6WTGH/P5wyHzAwXClUSwUgWEFbE2NhY6h+nu7+T3oCUmqAMi
tHQkiuBBX0KEWKwKps2oQUOrs7FKfB07BXSmrmtQbKFCtSaazlNnTFL187+Oac8qVcm5dRcP9npr
4YbWdB7I8/RU5yAvol7efuVnQ/0n0VQ3RzmicK/mM/4geSjxcJReDWnh7ruYe8zabBoCBv6hfp91
Dmn/XkatayxAWKu457jmSG+awbK/mt9CdUNRbVwW3cxAyXxEmD5f94c3vGg4lGPzP9Ko3GVxAW0v
t79EzLMnNUTx3RQNTgNJgeFiBppe7ntqhdNZNRXP0ZGSB9FgqcKdrux+nf3gUSRtDE7gt+W0lOhR
MOdVxKVAVwJ1ATMxxvdbopaZYQK+f6eYiVcTYkjoi1fnAIX+/nbjzOCuR7K1Kk6YrYXvBYguagKZ
GXJdY3E/2+aNEvR0djpVKoJDm1tFWYHRCl9zh/KWgtpkAZV9WpON7/i7huiwh2zR2Gk43UYtH57A
pbxfOPgciqm+adR+uillOA7bBCWtn0stuZYJ4P7lvfVAY5a+VgHIF4Kh3wXFkCPYxxhN+37C+PF1
J3NerlBsYGrvbWBAK0v+BFiQuaJUCKE8+fHDPQ7mSiT+t70Q7MjDPoS08QKVuSjGb2LXxij80mmv
wCGqO7Jv01b5e3MKle+LFq2efUw036ZQ3MR5P8cS47cvUSM8og3sKa2OlJqBLzdeFftixEVjx/tb
AEyLlTY6xCiNspykEiDyZUpY9obTvBInE3Owhz84vKFTi3CD2XA3ZDUd57mLStrfdFCRE123cuvJ
tcCA4EElZSWSdrxiuEmICjyHBAuPqd6s6232XJmMIxOqZj0jcZK1YowQJ4FSy/9XHMoaI3RyYjx8
r45M2uJozCEN6u3DvEUoJCAbAEj5ylcRSIuOqRYKSkwYjVWXT3/29c78J+UckOKwnZlT/2qxY4BD
gtztb79RpqmoMwzb9JPIRw+6MtgU4DrO2x+006bf5xYZAFiTnAwHlDKEfbCnCRsSE1riAt2Ty56m
zUkj0Oo1agES/Mv+3jqAegxjA9V2YHcW6c3xrKUYMLfIaCKt5JJ8XS9/YMX26T0FyoRFJNU7xoQR
ghcG5PGuTEaeFEqC84DTc46VWPV9MHoYlGe/Et29q3OBFfTsPVNrNKOK03vS1Rst8SBXJ638Q/4W
mv5K+sYw+OHHmN9HFfavGfokdLYwzu1JOjs0WDmiL7PBl8Xouyu1plhn+/4gGSH0MNGTj/SNzsfh
VRdo/g/gwC7MCQ/LLcwswvswbI7MeM7XZTgRTouXsEYcaA+1sBoQt5xc2VWrRN1QtBnceMTX4nMe
oBUNccqsxuVpZJTSgDjKBMV/Kh5nk1/dXjzHfgAddip1GpYjg+XQAqqWb3Ltm6ECO2CJg2LjJmY/
W4DeAbo/d37H06qMyREvVguOgb3bVCgIl2qqQPsNLc9lnHyQK6BlfsrBztjvKtOGyCtRnhfF7QXJ
Kcx1DL6uUKgzbZ35Oog7yJvlLatqPWCmu+vbRmbkEEmZJex46tRdQQQPblfwak9MrpIM47aqXU41
4k0pToZsm4ECZbaDFen7Yr7/UNnWqbYWj1U19bLKVRBhzpcAsIQHIVFXWZR4scercq7uUP5MOZMQ
5xl1MViDNPXtkH5l+OTOywqMzSsaL70kImJ4jTp3NcwOOnqZJiS5yJKknpRdRn/4L2oRqE906fBm
Uvy2DalIxioPX94E2AezsR4NeA93Odpo612Vld/pJdyHBTmBB6Omp2x2MQfMBlAbtMfv2en9NJfP
oxhk2SGaCaM0f/AfBsG3/bcwYTolpg+M0QMzHj162/+Zr3uRKCEYJqcXGrGYfX0Lpbz835a/GL8E
+pYNZMnLyv9XVHwu8uWl9eMyNrMdiGUH6voDwdw9hDkW2yR5m034vNDMNedL3EKC9DToZ8FhtVO0
fgKoJtgpkffXl4N566+7aPIukC2EmMbKuQkwfDTn/VRRVaclXrA2YqR0eS8ttuCGRCPHkca44xWU
gr8VF71STHinj2gnLTEnbBc3lCnxEOcElAiGsGAlzicEEPyoIC7spYkoPIfD5nIdoGxYeWE9/R1W
BvoX8QjXiIXKd/OlWGEZ/OpnqtX+jmKyAB9lMWa7AkvOnqj91WabhABHVQj/KceCWa/tKvfgdSNv
bkb4Yc09C7BflbJTpQqoseXgnR5Stb79QT2OCIYXy6VlL9KYGzk4MyWx3BGByORIvWLnVs3uuF28
esofu6PlxAgX1JRMTPg5dfoxji9SuhdU+kDiwgSf0aWYmnEeeWd5w1Z1DNn9erCD7M22cbCIOrMI
odniQIHkdA7uRSZMCUIQjjEFhGgO9ibRQaH50rgHNAzjSJ4DqM7SS1jr09ag28mI4tLz+S/8Z63y
L8Lls9ge+mS6lQTI/D//DX61mdVTdSc/xBSFgwBCLQna+b+NOm6EijSTKmmtomPiuL8ONp5a0Wxr
g1r09iPi3s0rO+0ALO2USEDzAo56D4JIK5s5owbBUIDqusSxPpIEoFqHcoSjFkJtl8nZy0RDz1KI
kC0ISwbM3wOpwQwT5zKSQ/a9Nv/6fADP/brlrWZU0UWJAuWVFYVeq+rWAXOyWaTN7nB6mdUxcSqT
i+lM34fktRIgpJ+LYBVhlgFDIVXb50Ok5RV1Rz4JY4Spad3U8qG27RHyKC15XTXzEK1KsASaF84/
N54LD1lzAqq+UI4sPJexAwXuhzOp2lX5XnDcvdIXDZhvcsxSDlLJzYvQ0he3jkZske79XsSLhxLl
T//LOetBm7rpVuBqlZE/7SnFYMgLRbyW2cbisfka4B3GupUM0s8TUb/VN5Z2dsCHzRfhrkl7tfiU
cVzNwl3Hn60YJKJjCRyMaGog9ixfG4wEx6K6Ov9eMi4cf8cpFaVD9nlKNijdhaNRxUv0EsaEuxmy
t/Vaouc2uff4UZf6pns818gajwhGkce2GtE04qmsd+6z8kdJ0ftOSjYykLea5T55BN3cMbG1emiv
FO2uBQk0ORG63V1cTDI/n3TWlSYkcjz8fTNMYfLUOn0Ul+oZO84lR48aOveH4C7ZN6aYLT5ayyI1
brZhSJeeN+e0t5txVZJa8c6YGQVZtJ4MPAAI4sJnDLHlukXHzk6FUy+VjById7PFaViMQy4ZE0WQ
1JU9p11R7jJ7mUmha9gi2ZLBfkXz48F8AUsxzBLQ+UH1626NikAOCgvARNY7S0B2GtMetb5cZ907
QsS/NAfhqMHWmH68dEkcVHSkFnMCDtlEmfgv/Z6Brz8mYjji5rnq3LPOnF3j56IBp1ZMkuNmBAC0
DpxTbKglQc6ev+VAAZWqB6W4TCrSQmUn4PBtStAdgkSRZnyRR+35bIn+IOA4vAHGPxSkXwkF6sDK
r+h0tOXCZNAXFNROZua8GBlQbP1n9ELwbopwjSV2xMTnaBEj2tA7nVzw74BHOKsfonZEqdxm4N6a
crx2NWH3oHi02Z4yefzE0pgtIvhVIgiZ8TT5FHMZThZa2qhwSJ5f4Mfeqo0Fw0GM92nInW7NMz7Y
fjpNu5ytc7LLEZp39eQebGLufrJvAyqeP2J9WxNbyN1YjgpurZNQhEzALhBrgus6Qg577TOBP6Lf
cGEeYkogyTgZTFoXqG5E7IgouC3ANtKcXpigE3DbDXvC2Jv1s+rCa4x+0n2EpQXOSEiNebyxm4b6
2+VXMAcjot3JXbEk+A4X63b0woZL8jv5xqDigKEwDnz7dDPfjuZsrr9Cjzp+eLhPHhVnyI/EbzWy
egxkZje0awJkq6axFwL+3g1jWl1oblCVWL3f/aIiaCtGRhtRNFY2n0Je4+d0o6OWvBsyXKUnlFXg
KwddOD58PzKVo91BDKW9rPfLPetNSFBaEew5K6LSoppGoJ6UaMPbLqsXwsgBplusMRH9JadDW75n
cCYFySVUvBWZm3W8WMrgkMWuqUnlfG4rVleppAxeKFb+zYozS0VtNzlMqkVCHB++fZjZ1xrWn2sF
xbbj+X3tUUpxzzHd7iQY5YOXFTrk56LvE+AMSzZLhQyyG+qSmAbWzXN/BlohX9f8SoQADyjIC2NR
WAMKjavTETlxBcr086KUXHwi4mHhSvN+l4cBQqvLN1NvUTu9q7PU+/CthSIeDvM5T+amzOv6iztz
gQDA87VdSDbH6bxiBmqW+ymNitDRArsIh3NGauiFLrTi4T9T7yP8lsR3ovsOf8yY6v2avYFt4NVV
R6rAjZEqif6aJtMtK0xNTz8S2u05LGLcVTx/08lG5C0hpsmoI9d4ukSY5aVaiDDd9zITUYgzJCI/
4K7zeSsdKukAS18dg70yVza+O2uR5pdw4Jl+UgimZYabBGXEo5BrGcRA4147GIrgmwqkylpB1S1M
atKWtrFKaZCRLce5PdNhP0krpmYZBrcDsMcsWnt2oN8gFUCGmJbkchYtFBijdF7EzQaV5YA2Xfn/
WhPoDWvuwcL9+eSJhwixCY7oLbd50uTCFBASTKChJRXbvcl8K/drk37v7mBLpDgBHNN2o0CzdKE5
ELEy02Xc77hQYStHa7awXJf9pb0FV/NZloGrN2lMGH+Cw9MvwHI33XzFWK5gBlkT9w3z0duviDTK
IhqKnrY+KDFE3Q/qNByWzJ9VjPbAB9N3gxAIbE1MBs3HGQRk63G/WrB0iTMmEYl1U98auOX/60Hc
Tp9HqZ2P6nRnlFnYPHZvjfiS9jv6xRTGG4pdjLgSRKzj6XGn5D75oGQNs4hGzZy13d4cI8QMAeDj
PlODAHFr+OoVMhJr3ARvoZaI4Z0De4vdkxp8R7SQlUW3Y/IIi4HC0vK4IQJWvsItucEasQ/rbOhl
5kcg5tMfeqE1p+FpXs+CQL2xjvEdPxgGkMyyfjBTlGB/6T/tvd5JemDOMoCi3C/3x2w0yiE524Qz
bDMnvCEGTmKqAtjc8WTVTKTqIqUbr2wGpTnQPw5e8v75nkxeXHvtZl2OwUVbq5EoeDbYJHY/tPHH
xxS694J4GHswb8crZe3QkB8TQp63IRZR5ORv7TqJmUp9uzmOTUk1sjnTHhcjunYFited6xHZ3aKg
jehqeTluZoQZV8szRAFCKJamQtJ5ybPW2pmUjMYZ7wDHJgrpuG/2EjptUMM6JIqIOb0hrWSQBDg3
oGAMC40bqHVadGTNURJjlrizKrTjpk2gMd2a3eM9MhDaklKIdMDLbiNjIhd2ttjgz/a2bfJLCfry
+uycZERJw29c3SrC0lFhf3EnwRksL7hogTBpoAMsUgU0AOBWndWNFLtRhqTFvFgw1II2DnzYcQHl
CyV/VRvSp8G8yLEdpkST8L6TTSwPFhCTvwl4YXSm14atz6eUOAjxswwiuqlJitYUvEoOHx1T3KjH
rmlA9h0/P8hoX1/QYMo9imCtCiOau7op7z1Fxo94U2gSp7Gx6Rt76kFE3NZFb2nTV39rExUbfqzW
3PmoFB4RtwW45bZ8Lx3mSr/TzZF92npGiSozpjt44Zqbc0xJss/CEPBeEMk4AqXZn/k2WZuUgvEA
rJTJ5PzraRlW+mDdBRyxiIDt6fvHrM/Dl0anvEZ3B/3wGfn0COxhVy56o7u15AhARQSk8QhFsVR/
DDaSVcDIFN5+oT7jn6pwEURsov1aRyMzKS8j1R5Qm2jgbIVIv842eiSiu1sYjVgtKFZZNz0nw8K2
OY0pByvJk7t+CkH8G/QVzdsRxWNA4cwRPKyXNEFeFo6MBz7CCn/vqAZC6RbmqPJcbn4vwzRkE7NA
UvJIWopvKHa3UvTuzYuwT4/czLz3bZrxo4qTn3RsYCI0Zak5QCj+8EZT5Rfh+Bj/nDXBrL6XYMSf
gDAgv/UYbAzX31RSIHmMYljKFCdq2sm6+DLkUcAMdDpqBG8M6Hsd/hn9KHFpsPwEWv3/dNIm8Ft5
D8UQ0zU3kcKoGVm1nSLKqUOBl+Kl9pv5WfxCff9hTNQrjUPqDQovpfJWUQtAOADvyIfSP+k3VIyW
pVRm4Uyxi5JkCX/EpojWskQlV+kxMUb0uoDQCp6B8ISysq2eA9qhhE3lJmTk4bKclmX1sylFAReg
CjFUa4CEhVohSWJW/DOAoXOeGwolMPIyFOtIw3Sdn4jjA05COUl7zXbSHNOpxIb3cLKCXrh56H+o
uJjKJPuz7k1/eZTvaKLMP2Y9cpyn2/Vn8cYvX2X8twq3bdsFFwlj45D7ELRkkOEtCY/MeHoZ5JxN
Rn30WLCwa3dTXo3QY+v93ua1lYsmcyfdk/NJQXj53g/uRqBK7xu590mGfhnyAAFluooYHJ3cymQU
nkYsPQyMCnVrbp+V+VJybO51NJb4yxCo6X7PZXWu+wbNIfuPvXvHs5VA8cDHSNSUs2LN939IGiV3
lkCyeoFLgkG7gZHOEQtaOPILourozefRYn5UBdcyAphj6Nf9NHtQm8WBAEQC4P74Gk+vXYtEUHAG
YJAO/MtaCkf/3G5xbGdp2Rv+1LvUfwKFn05DioY9iYCzTOErGoOvTrw8GJ0jE8enb+kA11OFMMO6
0croAidN59Ke4JAyr3IU+jSPPGsV7YX3XleMlfRvFQR1sPmfna4p7sN9KiRP9VOvRNjeOfjDQkAa
jt3OZbZkZH5eoG4aAXouCTTkrxJnvP4pOGGQt/pMTNPrMpAUBEHUVuykKMJdz+zu2p+TybBrk2Vd
/ON08stwOlaz//hVra3NUtZ+qlVgDMdjgi/Mg2Dj//ONd4Ovl/tLiXzq8cfupyrdVome57jLsunn
89us31AKTLvA/mwCGNgQoBbXlzmQJNXqvPeDYPJs6/cKDR8OsaonSQ6r1GwGzkxU3le2WFpTvVOT
YwYOcSbs7PdXr15uvbyECcPHafwNpmQF50TdK7pcDFuzisiQCGLIrbadHVLHE3Cx/OKE2lZeOPE+
sNl23skgP/X45X03jAIxVFhKFpcNP2SELeUQmq/vgIV1lsUHdQEXTlKrxjsg7JqN6M9uvYQMDhoR
i8EAbJ6cN3lk450ABlCiy1WwiOMws927XVX4B/f9i8OPrIcry5agCN+cI+fKyhAlqzT97gSJGMmt
epsQ0Us9Xqk2fDf6WZcqxYzIWWFdl6wSfclRRwylu84/VvaifdMm1DtOlrXaBzYkp0APqwGSuTBQ
G31c5PGILrJhpPJrlkrb7mRv57ctb2OON170Tz4JWq2vYqmdeEMM4WZ354BUlbKwBpLtTzNKJr6K
ghXm66zjyDt/2kUpKKtX4AbkNscn/q0vz14Sjcr9kjCn4L48B2D907FJyN5E/NwWuL58LxsjvWns
OlJrlqWX3OnxMW6f00sEMtBZuZuVO6HtC7HX0oa36BMELYjvubMGc0yQvwQYY4R/Gu4angxwRew4
bBDX6rO4uoxAcXrnbmEjgoQi10FsQC5jirNFeQzWI6wDhD2kDt/8UGH4kXWY1HTLXosiMcVkHNfu
r7YfJZPeFNyr/+z/5S0NFpNH52SfF0bVoYgBhl8mtjR2nF6bafeMA2Dv2Wu09ygzYBIRG5UxgLe6
dir5PWTTwzZZhLJoSdDqyRoVbQ8pH0PO+EL+rLZJEB6xwnsEO7ejWdgbKrQM+cp1eV4/p+up6SMz
49kUaS4cxxq51cPXBwxJU+gAgfH2w//kBJ2zlq0YtqzItc47+Wh28r1GYyXNY7lJqlafUDbVbxsL
uzo/XHMu5pn/WhiBnxdGN2HI/nLz8e+jGw/bLqiFUgdtHeIcQ84t79pztKiL4imXM4OhvaA2ELWw
HSgIaN+gcoxgyDD4QvTwpYzqaseDqo1c8WnCHwRnbteLzmvsGkAYNw2KhSrnyt+JQaArLD+ZJA1Z
DnJyLUQTODPKGNpW5fRJO+wjw1oUwLsX4G+5ULN9jJvJXxnXHtDJVjMOXzdFkfxUGxyxfxQ93v55
IQtULMLtiBJymcCXef2A6eyWtf/Hy7R3gRQQlKGg3rJpgv21Q7OIAJyXR5Z56PWnHITPXDNTpwXO
/sqD/hqgXHX/Srnn8Dv4h/bJF081eLMcBZO9F95AEgAEXiZA9Eib1i9C3R5GaqRI4Ah5qKQzKSdF
7oJIj7mvMdHML8jwHnrNhsucCzlrkD4xvUlb51l8MLlgOIDxgJdfA/SNKjZUPEI5RIbE02FCUR2u
wju1ef/jBMcrdPthTKOnjg7ERK+vT/K604bA1IZD03BysN6IQU3dwJ4e1dmJBthZoBclIpNd38Lw
WgA2VsBsi9Hdijl8Bm1eSKoK26gajMJJBoo+cpMP+aSoAsYUf25/jX3JEDMh7pEar8EtFX2r5I6W
WnebxxQ9iIVPp6MPYLpgMG4AhxETvR7t0MRdc0b8fgyUWgT+q+t9x64v9qHuGVIA3qgqRsL9FUGB
9rPCot9UHzP3112CS9btwwA0jA2c6vWyhVdJ5lnf0ctpPryf53vmEAF9HsyQ4+XWLGsDm+dBaKGf
VX698ehvdwk76iyOCBqBlhAriEvjSgjIkxRi/eTYeiYYGEvh3uVdtFqmOC5e3wu4LmZOpFrsCHw/
2WGWVIHBen0cNF08xCy2pE11DR9Dyb00tyt3dTvUADE648ALPgvBiPH7S1nNpYJX+NJw31qHWdyf
TXSO7RRcDdmngcRf4qadVvvcpfszUbonWJDpVl8CLbgmHnf/1iGOcBKnKa0Jjt1kgQMQOZhzmuvP
/O9D2Dc3+7bZbv4SUJ5799SVvbH6YLaqm6wEkyTpL1Xe8tDABG26nDVTWD6zrfiovU2I3Rt41oax
++d3Z7K9KTnqrw2evaFRfJRriIpkf25EZQY8WBueBWKSOc79gnYQEeIlDr9w4B+eLn0Nl4SqZfFq
khKRwM3mW/vXHuFV4+4M9B5QC9XxS9N9wq0Bg3GdD5yXMYyTV8AKZxUXU6Im6528ImQOs0t6uAwd
JgfCC6CG+HePvRw5IWQs+FJ08qdsl54sZN07CDhcA8sGxD9LB7YU4H4Qmdgm49odJqmofGKmQqZH
OWI8Fqk2LukYY+tib5F0yopzKNPia1fDR1pt1KgFSk/dL5exZ4wtJT2Jjc+wzWNVhaemANr+t637
XKvWumObZyd7kIrdFcZuNrtaSHzQK0qYOGP8Bpbr37bgaan1JdY21NaSviWmWs2hsOS8GGu9FSlP
kqTjOD9Fpztn0BSQzzuoM3DSvfgU5lRr5tdoxWKhZdubpLQrErB35llJAe0zkkMJZkkFvd/wzoVx
nsfFUTzBYBVbv/YNFMscTL4z71vfMqFJLFJ64uZPlW7QhGTr5haMpmT9LkP71pk54Twl2P6wlDcn
3KjkbnNtpTmzRXofuz22YGWztW/vDntIo6nm3YciXLsb2clSF5rJl+QUuko8COTTV6B07LsHyLMR
jaZfbjVzEjFokLil2HXhrqaPbYypZTVEB1nvuqC3D7wAeoU6bXHL7lCEHT9KdFAQrY/SBuFuAhdN
tIp4Q0DXY8IPhHj/aJa3hychl7gyZ+cVmE4rIYzS7oBAwCzWp6IuJqOqjwHbyNanjYdT8OqoErga
wqadgHnoslN1bTXaTFmut//rvdnYNRpAh4yXLomylksWeLnWUxjJCmBTcsgd+J/k+jr0RHbEKH6I
kBlUkeV00TTNIPl6PntUx5b2LD+55M+bjIz4h8nZco9rBm+KV1DfcJXBk1F2eXo4OA8uzkiLXef4
oieyJclqgRrFufhWMkjIWbLjUjw5NcNAU5dzL6mmBCnHxZeFIbgWoblj+3pWFXrMDvaIPlhRQTPJ
QLbhfh944i2LSzmHimCZaXKvS8QGl1WaJXp+GLyxVa+jWrkD0QwdT3OFeALEJPUiErvDL8VD4+LY
vphmSYi2rgZ05hoQTJCgMJLF8z9gtNr9nqF5aSqZBI8m1nROkCDn/eyqzVv+iSWIimhmmLefXQ5b
yqZCqMOH9WekKuXcOqPU4g13w4AFGICKDlonmHGLX7qtFTaFxVVOnRJP7qjjlwrHctnp7Xj4R4zz
CB4bx2w5U5UWYlVZ8+SmqSbOfd6DRXUa2Mhs5V2UUBWdSRGQgw+JcTfTI8ji3ILv9DLAIqaWZErt
Nf7Y34C8gcgkdSeXqAFUa0VM9vVPIkKcLl17uAHMZqHueWigEQAT/9BAhkFAn2ymM0qQVuEcOK9F
AOEaSjl9/9d479ajIUlDvBkQqnGSZFWhrRGTNAMK6LQ0j5MqfavD63f07HNzhM+q8o68XoxgcS7y
hZHgUUBPagM+NDMFkkDs8lfe2Yw8P2h/G9R2cTo2bEuQany+h4FIFW72u2lPlCr9YPq994vz0d/B
0BDwnycbpgIUKAxSDg7pqvN7qpfMte5ybekNgUyHa0WdY48P1+hKVGEaq9mddeuNIFHB0Tsjz9tl
0Birsxt9yqtu/0SIIFVghhP06Ohvbl0RDYAmWenr4pfFtY975hAuYxam1KPEq6bGLK3vSIsj7r+B
ZgHuv9xgH0qmK8Te1p2eQ113Uf9VZeU9etk2PtvWOwA2A5z1nwi/TD9mk3eQhYDnlqpZpHWOJ786
dkETlvhBx0LmVe7WSqI4aXLKCflnYuwT6GMOXTeUUqMxQ2c0XWQAnqky7mxiyR2lgOVy4lFw2/jr
QO7yc0dlmx8DFkeM8ty3md9PV6wpOwJReh4XjPrDsXtianHrtUCOVrkg4cPunjR+Yk32nFHuH71X
yJy/wAsic4uDNs7DNn6SH0YClnpBmFmkZnJ4DuTuFR7ylhDxNy/jufih4pCg4Ji8xwyxdAmHJb2w
GwdZL2dBzM4BRiHd5BBH8fDBcD+PhYe24EtPskDvyWeplPWGydpFaJURXuF7dMDLRw4LVX+uhB/e
nxSXgVOpWYjMw45/Lopb7o0wS65yKq9s8W7iEiv5oD1nt+OEe5nCvr/bcFgLAzRab1ELDCJMUEWf
I7wBO40wVP7gcm5G61gZZWUZLhNE2awqfchvs1D6h1n88XzagLcM7tbvhho2CBFe7luI5E2JfJGL
+nWCowtKNdYDF05Dtm/1gjrQpO0WiEkrzHfs4x4jJsRdHDHDLRGmYejgRSLVOuHH/r8A8INvjS/A
4Rxskv2oaqK0Z2s6P3xPEqEB4tbenBZDgWaEjX4fko3zQTvgWCxcIrosPpK3YhWAH2CFdD19t0bc
P6D2lKLM0vAv947Epx1Ktfbb4QdHbJlg50SsIkRQzzf9rJqbKAOqVu+IrU1Llyhh3dxzciIz8twl
OuFRV7AIfJRNepDdJlKGCQdDnGCF3y7utNc4nPUGIpAIeM8CwZ7Kvauu7uFHKuND4RNo1odAVsm8
1dgaR5bQHwu12NPuEguIw21QW6GAZRXOxe3naPE9VoaoX3uB21jOybFmLzQbewBk7D9lCpL6oh8j
weBU25hq5HHKVgSItnFVdC96k8X7XEKw4FRLIwmEMNMxF0s61AItklYXwdeu6edrlo6ISP204nMl
gZcI7Lz8x9hxnglUVB9xAxh1Z6lL9Ot7NfFr03V0Km9DB/vgNWgvoxPRyFAvpv7IBI4/WJN9kVnx
qR9q1X+ON1ygdon7UrS/eMLcV+/IqGmC7ylUo2PN5MA7cIb7VAqI0gH8NN6N1vnIz92O9vhZQQPc
ADstzfSafJL4XD/w+rGPd2MQhuuzkKBrDJiWwvvsFrogWrOhwI0BtrxVwG6VAUzZaGyJofKzsIBn
ufUI3OQ7TSejniXevEwLMbPBspjg52sEryrXqxnx2jJPwO8X0b4Rhzr90+3Zrsh9IAmovQVpQ7iE
lmcc4W3niXYV83OIEhMQNeT3gQdD+6huL4ZvSX5Nf/+QyBDlW6LWctH8sN2M7VHlqfRPPq+LtTu8
LhU1LQC/WoVECflNSwMzO51wrKgHcRa4uMwmb2UCOM15g4asosXWO2aH2QhUbkaqlZdROtDya6Ot
wqsBkVAr9x7Qp0T0h3A6IX890Q8apUxkLy6Uo3tva7KFHFxYYHVH1BGNgNIxlszY0caCJ9SaQWFz
yNuUmMc7G8o4wVbsVvORQx8F8whIxYRWQPeocY4zvEGmFJ8NG4aPicziQBDAf54cDpvHsgyHlMxC
d3dHEQhkuiZ+1r7wiIYh/yi1U/UzSRwgTNngWqmWHlfml+hN2VxLk3zqUC6se9fWkD1tBnulwl9X
V4x+X/w1REI07682c9pmgWqWhVyBwJ0ZixnnH2wm15qRrLf6qzJhAtAPYd2IJnVT1fRKAaXZlVQT
sDWdkVsM9XSsxCV8O73Zcl6NyL2+INDGapy6FAzkAUgLVBqr+jnGeJ8bOsNVi6B9i1S8OQnqFLst
ZuS+IWNYnd4B3oo0CAdk3HIo7a7oUWkipNf3ofdLXJ0b8MGVRxNdneVx68GV9Qtb2O3LWr9Jg4dm
cjJZWc+mvr57aBkau9oqWcwIi5katMHbUvkl2jHRVuvTLGYNqk3j7oq9G+4ULdjRC8+seDQXp7lu
GuUpBcws8c4PiyON98u+/9fDAdIHlyf6ChAfmg4NEHtyLreYnFO6jaZtUof5zxl+NGg7vG76ShLk
16YztO8Vr2+3n+v1uA9OA+GhZVenVd0GjEp4K1/0TDwApbTi7xcwa+rUbORTYeve7xJfr2jMXZRr
WFE8ewWPatYLzhn6lFXlcsDtXvW1VMtxXvh26i8ldxZvqBBxfqqNitAvTCYizYflS6tpUgDrD6lr
XWJUBgOak6P3vqwaZMDSmfcQWscklv84qANcOzjuWaFYdwPaibVyOeKjvU3L5+wA44iPL74xcI2k
4UuuJ1IcUfbCSwyq04xCC13Jz/UlFtJN1r5rAj/npwVr3k0BIE5rrIIpd6IIoxOWbL5NcYn2OqN3
IjcSknVEDdNUvmUivvS84l7MazFPe/HGPa4wTR4Lo71tzwYp9r/LLxip9rO3C35ss9SMNnYcv9FA
+mYVR4tjHcvyXmk4yhuS4/yRSESD+leNrY5lzO2gQ44O9VOVYzYYDFtUIlQ+bWDpAcQ/XOJfB6zO
iP0lZKoD10GYZdr6jR8jmVyjIM5O4LTCNAVf4V3KW0anOoVY6HzfGh+yuQNe9Up9Cny9wPqgbIKp
7DKPBx3TOrcan6WprfAl2XtcA1u4RLKVYVW5Ww799ccClHZRufBxTSXXrOv2SKG+7AzJeoIpntl0
5gHEx6YhoYM58Pa4muOZ2nOTVw2zekUUrRcXpsLc+2VhgynWeB1TafydylNnLPeM8CvtBB9V5k4p
HnuQ+POESZ/NNW4dK1dd6XE+8LmdyteCPlGYO3e9w+mIkbhNHGs50VstjmvSeWnxcy/ZQfaKZQSl
M7hcWKdgsfRZv3FyCA4TVyZK84xtQaKvP+yN99c2BWduCZP5Vf8rvGglec/7hhvkmeA3jeu7chUK
yRy2Wz8c/zZafuNY1BIXX1ftiOLw8Q4tYFD+Vhlca3KU67mnG3Dt9B0zwKbv149ZhqdDNmVLYh17
jJm2yp7CHjLJ4TLdhqhg9Q1izftph857lsx68YnaqDs4K+XQRKLiY8C9YKndFWyxF5rYFY5iNC3h
ahqKz8K9sVB7UyRIuxJYaqC6CGHCAp+sCMBKHcf7q9T0XC/1BuNJbJuzt/tbrcR9zhSrlMARuH9r
CFc4iy9jnowmTMoaBhhV0TdyxES3uSbatwnVgEA8JM03Mpvc3LSI6H6bWqem/S7jFQZaV2Ud9Vwc
xg5xQPQWyvKVc/dHEOSIBugdip57Ply1Alf6un2/f2mAuoH76WfRN/aZn/HvkqaLtnAac9Y8or11
ebBd+NsRzBkBfRZ5k9A/5blu9OMGAbIeVDVhBbxTy2L0Nyt6rS3vi0RWvk67qc8Fo8/2G84XGSN4
s2/A1UiBjLpM7wZoF3GA2puK6o+HsDkRDQENAvXcBP47cKDGNJbGinv68NGikZIXm0npymRkXGy4
qGn4VtijI/rEglih4ZFdayJP62d2yzSa8POy4bnC+6YWhdIpkC8KoqWTMCP0tLTc1YTWZb2fH/is
Y9eKDZRLfpp71dUtxvAljHyxYJI0i1EUqNRSKShTQmMpGHseFCMcg572gnaGzeUyzwvUvV2rzR3D
r00fXFwxVW1wsOCDuanZuDlAIvBIc8kLOc4puGyzmjXC85HLjyksZUL67bePcy3S6nkg2RC74rQ+
sUsIg1lMZWpzTAYI6x2+FNPq3M3A5HtdZORLOISv+K9/5sc6gQhE3w/PZ2CyMboT4scWyMELf+qa
SUNGYI+iRyTLELiaZ07xnbnd4y7z3Ghd2MNccQ/c7Uj9fueaWzbhORwarK8xyfPDflxtPKqutpdl
UzlP3/5uDER0fmpy2h1BjNry5684oCtxlDBUZqubC7K31X/qM2ZiSdtCc1g+QlUG8ChY4SZEST9o
Ju1TCF9IlmEIOthB+JofNjuOMH4DYflxlC+lKDw333sHrJtSLSRSn/xpmN4mPgMklj3coxwZL8HY
D3G7GyH+ttLBpOzvXTu1dg89rv1ujBugvTpa2F1s2BCCFVCQM5IZEYQihZOqK3USo/7ui3eM3FdN
je67J7D4uK0SgKEc2w7alvOtMjdxzHhJzR3sdn+Oj51WVJNdG/0jFXng1D7+DGmjmA61G7DcRfeF
Nka36L24CykH8S+kUfCdwwYTb/TkC3tevt5FEXfE7KZ2ifytCLdyvwf2ZIzYzWx4oaxYmQnupZxF
1UNFX8jSutxWeK2FMTPr6MENJG05H/j6BYCxultCC8xDGWUXw5v5Yp+c+LioiwllsN33KuDByS/d
AaZQP0TWYFvM6VktetF+nKFKFeKtQrqBQxSie9c7yDGAlFMaIbU6WMcBQdzX0AZGqSWY7cUwdFnR
Vufv8P/OrMcCQhCnOlnbJ+Wdr5zK+82CRt8pYh5l38x/Gt1kwDe9eSUjp5slXYYQpIaSH1w78ft0
DogcGkydZ/KqD/IRmD/F3QD0Rz8cGTJFSRKLnSdKcW7z01UngKV0dQrY6xY5+l/874P0PZeuN1Pj
SgyY5lRqgfKH6JaOTzlx5mYpFBs3XhpWYJkJXNod9z21wzDd1WN70nleQPN8lb307G+AWBG7XHmZ
k2g+KsSEopG5zsIKswb5y9IfFM43EluCjfiKBo8mZrs0Zwk3ZiLoIkxRM1Ov3Ozf3WXUhfm6HmYK
PRo8IHJaFi4tpcj/Wo/MGuSF/ODltifVrJmIbzwM0DSCeIru0znk6gS4ppxJI9eja3NH9RsNxRll
9WvZiRi+bzLozOkOhRTrJc/JeWZvcZINRAVOodbE6M8abnnXRCR2YeVa+ax0gMTz1ijAHkNPvqFf
chjKXG69LUM1Ifnrsb0ZyypzSFZo/EvePjitXMGefgenGbvUypKfUEplthGxF6pABRhxei+TnfD4
A8mXBO0+xXI3srK8jsnyJT9Li1QMufTBKwCzlfAPGAZnswKX0LxpsgObp6g1P5+BxYfSkVZo8rxg
LVervp0YBHz07Avvpj+YEQAfGQkorV0nZBzVNwUJNT3zYwdcwodrrTRXiDmvYk6XZ6JYgDio8XL4
hpq/K4MnIqL0RHsj/44kQz3KrBvUB2hcqfE4K/00jx8vTkhAfW4T6AESqu8+sqWXMLP1n29FrzCU
WVpuKVxqkLh4R+2YQZn5vqzJMi/ktIZ8jrPxbdsqp2SzEbQrosIDTKgHNnnnl6xgdjLycvB9S90i
/qDgrzcTBiuesfcAT9x1HD6RtCwIf4QE95MKVTxfImcCjyo4GM1SNXKuXr5ql6+C8HTBrtX5KhMY
w8xjygyqAkIIlONZOI1Cbtmt4rNhv92bI5HJSQnipUBveUVHlXRI5LPp1IGmQSgDwih2tCELuCgD
jo/TlgjaZmTRz4IEXb7NeYfUIdE6w4YHp+jAV2O7byDj+UE/GqXOOpnksEJCViSPn2ZyJiakkGlT
Pqgdv/9OaJuG+p2DGFG+UOZzgQQcS70SWSq1+6liaU3A5qh8gnDXWcVTAyV5iYRhjTXq39L7/uEL
IVeCaTbFM4l1aCzSchFOslpCYPbao+pAXC4OHVPZfsSw9onGAi+qVB6n7n20GvXRwUCIFWuLHreP
ZswAeHLEIDGpLDXJx/feg3seF7P1vlIsilssBJ3BrUMNE1lbB+4qT2mRJfl5a6fcgsfqg/GAPmyI
XhEbkhMtPFrBhVEahhvpk8wLl4pj5avN4NhbGqPRW4TzncOjBUJMLT9CcNQrLzBdMrtFp2/GAE3t
F2w9n7xOSXOQP8Zdy/4OC0Qw1Mde+QS1l9nOete82qyVN21BDEtavZiHd2PcubFo0a7uKgZnSjXd
5EXU8P1wXesneommXSRNlP4q7VYEFINtLRBYBBapq8WXrYZLxaqDRpHtxyGGArBhOEx71qlwc/uK
p33lrEN9zQzrPfJY0c7vkuNyZI8MfP1z4+u80XArGePpB24R+c5owkC535ihhUxOxk52re4gOJHN
jxvUtmASC7mNXyw1fRudrswQzsNlfkSySGreWvT4dEkIKDDsN1UQH3CwI99A2PRwtjjskofq8n9P
kLLuVLKd/8f0En/Yx4CsMYdFcWCepZDNem2Dl/guSRffJFwzkXyn06P71RlNLzKrb9i3dAwocPGt
xH01589vYxxLwm5nUQuAdleK68z6rWJZ8XWJXYbGxg5inEh7kkuZnKtDAtA2fkeUT6jcKlvCkTHw
enWF9ozpvvPzuy8cHRamv6Yn3OtKXjEX8GHrZU56GSbuGnzW5RxYgDTZkRwMcoovi/rEfExPf9rT
dgfVL9iMqSjRLVX/Dgsf0dFWgJhOrky7Ua5WtUUTUYc1a+SZp/Jv2MV+ixKGUwrve37wNQGknfBG
FQq/Dkgzigjum7LltN5Blti9hVkDRKp1y5cCQ8zku7lQbQioHz0dA2ai6xU=
`pragma protect end_protected
