.GT_REFCLK0(gt_refclk0),
.altclk(q1_altclk_m),
.axisclk(q1_axisclk_m),
.apb3clk(q1_apb3clk_m),
.apb3presetn(q1_apb3presetn_m),
.apb3paddr(q1_apb3paddr_m),
.apb3penable(q1_apb3penable_m),
.apb3psel(q1_apb3psel_m),
.apb3pwdata(q1_apb3pwdata_m),
.apb3pwrite(q1_apb3pwrite_m),
.apb3prdata(q1_apb3prdata_m),
.apb3pready(q1_apb3pready_m),
.apb3pslverr(q1_apb3pslverr_m),
.bgbypassb(q1_bgbypassb_m),
.bgmonitorenb(q1_bgmonitorenb_m),
.bgpdb(q1_bgpdb_m),
.bgrcalovrdenb(q1_bgrcalovrdenb_m),
.bgrcalovrd(q1_bgrcalovrd_m),
.rcalenb(q1_rcalenb_m),
.trigackout0(q1_trigackout0_m),
.trigin0(q1_trigin0_m),
.ubenable(q1_ubenable_m),
.ubiolmbrst(q1_ubiolmbrst_m),
.ubmbrst(q1_ubmbrst_m),
.ctrlrsvdin1(q1_ctrlrsvdin1_m),
.ubintr(q1_ubintr_m),
.gpi(q1_gpi_m),
.ubrxuart(q1_ubrxuart_m),
.ctrlrsvdin0(q1_ctrlrsvdin0_m),
.correcterr(q1_correcterr_m),
.debugtracetvalid(q1_debugtracetvalid_m),
.refclk0_gtrefclkpd(q1_refclk0_gtrefclkpd_m),
.refclk0_clktestsig(q1_refclk0_clktestsig_m),
.refclk1_gtrefclkpd(q1_refclk1_gtrefclkpd_m),
.refclk1_clktestsig(q1_refclk1_clktestsig_m),
.trigackin0(q1_trigackin0_m),
.trigout0(q1_trigout0_m),
.ubinterrupt(q1_ubinterrupt_m),
.ubtxuart(q1_ubtxuart_m),
.uncorrecterr(q1_uncorrecterr_m),
.gpo(q1_gpo_m),
.debugtraceclk(q1_debugtraceclk_m),
.debugtracetdata(q1_debugtracetdata_m),
.ctrlrsvdout(q1_ctrlrsvdout_m),
.ch0_clkrsvd0(ch4_clkrsvd0_m),
.ch0_clkrsvd1(ch4_clkrsvd1_m),
.ch0_loopback(ch4_loopback_m),
.ch0_gtrsvd(ch4_gtrsvd_m),
.ch0_tstin(ch4_tstin_m),
.ch0_pcsrsvdout(ch4_pcsrsvdout_m),
.ch0_pinrsvdas(ch4_pinrsvdas_m),
.ch0_dmonfiforeset(ch4_dmonfiforeset_m),
.ch0_dmonitorclk(ch4_dmonitorclk_m),
.ch0_dmonitorout(ch4_dmonitorout_m),
.ch0_resetexception(ch4_resetexception_m),
.ch0_phyready(ch4_phyready_m),
.ch0_hsdppcsreset(ch4_hsdppcsreset_m),
.ch0_phyesmadaptsave(ch4_phyesmadaptsave_m),
.ch0_iloresetmask(ch4_iloresetmask_m),
.ch0_pcsrsvdin(ch4_pcsrsvdin_m),
.ch1_clkrsvd0(ch5_clkrsvd0_m),
.ch1_clkrsvd1(ch5_clkrsvd1_m),
.ch1_loopback(ch5_loopback_m),
.ch1_gtrsvd(ch5_gtrsvd_m),
.ch1_tstin(ch5_tstin_m),
.ch1_pcsrsvdout(ch5_pcsrsvdout_m),
.ch1_pinrsvdas(ch5_pinrsvdas_m),
.ch1_dmonfiforeset(ch5_dmonfiforeset_m),
.ch1_dmonitorclk(ch5_dmonitorclk_m),
.ch1_dmonitorout(ch5_dmonitorout_m),
.ch1_resetexception(ch5_resetexception_m),
.ch1_phyready(ch5_phyready_m),
.ch1_hsdppcsreset(ch5_hsdppcsreset_m),
.ch1_phyesmadaptsave(ch5_phyesmadaptsave_m),
.ch1_iloresetmask(ch5_iloresetmask_m),
.ch1_pcsrsvdin(ch5_pcsrsvdin_m),
.ch2_clkrsvd0(ch6_clkrsvd0_m),
.ch2_clkrsvd1(ch6_clkrsvd1_m),
.ch2_loopback(ch6_loopback_m),
.ch2_gtrsvd(ch6_gtrsvd_m),
.ch2_tstin(ch6_tstin_m),
.ch2_pcsrsvdout(ch6_pcsrsvdout_m),
.ch2_pinrsvdas(ch6_pinrsvdas_m),
.ch2_dmonfiforeset(ch6_dmonfiforeset_m),
.ch2_dmonitorclk(ch6_dmonitorclk_m),
.ch2_dmonitorout(ch6_dmonitorout_m),
.ch2_resetexception(ch6_resetexception_m),
.ch2_phyready(ch6_phyready_m),
.ch2_hsdppcsreset(ch6_hsdppcsreset_m),
.ch2_phyesmadaptsave(ch6_phyesmadaptsave_m),
.ch2_iloresetmask(ch6_iloresetmask_m),
.ch2_pcsrsvdin(ch6_pcsrsvdin_m),
.ch3_clkrsvd0(ch7_clkrsvd0_m),
.ch3_clkrsvd1(ch7_clkrsvd1_m),
.ch3_loopback(ch7_loopback_m),
.ch3_gtrsvd(ch7_gtrsvd_m),
.ch3_tstin(ch7_tstin_m),
.ch3_pcsrsvdout(ch7_pcsrsvdout_m),
.ch3_pinrsvdas(ch7_pinrsvdas_m),
.ch3_dmonfiforeset(ch7_dmonfiforeset_m),
.ch3_dmonitorclk(ch7_dmonitorclk_m),
.ch3_dmonitorout(ch7_dmonitorout_m),
.ch3_resetexception(ch7_resetexception_m),
.ch3_phyready(ch7_phyready_m),
.ch3_hsdppcsreset(ch7_hsdppcsreset_m),
.ch3_phyesmadaptsave(ch7_phyesmadaptsave_m),
.ch3_iloresetmask(ch7_iloresetmask_m),
.ch3_pcsrsvdin(ch7_pcsrsvdin_m),
.ch0_iloreset(ch4_iloreset_m),
.ch0_pcierstb(ch4_pcierstb_m),
.ch0_bufgtcemask(ch4_bufgtcemask_m),
.ch0_bufgtce(ch4_bufgtce_m),
.ch0_bufgtdiv(ch4_bufgtdiv_m),
.ch0_bufgtrstmask(ch4_bufgtrstmask_m),
.ch0_bufgtrst(ch4_bufgtrst_m),
.ch1_bufgtcemask(ch5_bufgtcemask_m),
.ch1_bufgtce(ch5_bufgtce_m),
.ch1_bufgtdiv(ch5_bufgtdiv_m),
.ch1_bufgtrstmask(ch5_bufgtrstmask_m),
.ch1_bufgtrst(ch5_bufgtrst_m),
.ch2_bufgtcemask(ch6_bufgtcemask_m),
.ch2_bufgtce(ch6_bufgtce_m),
.ch2_bufgtdiv(ch6_bufgtdiv_m),
.ch2_bufgtrstmask(ch6_bufgtrstmask_m),
.ch2_bufgtrst(ch6_bufgtrst_m),
.ch3_bufgtcemask(ch7_bufgtcemask_m),
.ch3_bufgtce(ch7_bufgtce_m),
.ch3_bufgtdiv(ch7_bufgtdiv_m),
.ch3_bufgtrstmask(ch7_bufgtrstmask_m),
.ch3_bufgtrst(ch7_bufgtrst_m),
.ch0_iloresetdone(ch4_iloresetdone_m),
.ch0_phystatus(ch4_phystatus_m),
.ch0_rxcdrhold(ch4_rxcdrhold_m),
.ch0_rxcdrovrden(ch4_rxcdrovrden_m),
.ch0_rxcdrreset(ch4_rxcdrreset_m),
.ch0_rxchbondi(ch4_rxchbondi_m),
.ch0_rxdapicodeovrden(ch4_rxdapicodeovrden_m),
.ch0_rxdapicodereset(ch4_rxdapicodereset_m),
.ch0_rxdlyalignreq(ch4_rxdlyalignreq_m),
.ch0_rxeqtraining(ch4_rxeqtraining_m),
.ch0_rxgearboxslip(ch4_rxgearboxslip_m),
.ch0_rxlatclk(ch4_rxlatclk_m),
.ch0_rxlpmen(ch4_rxlpmen_m),
.ch0_rxmldchaindone(ch4_rxmldchaindone_m),
.ch0_rxmldchainreq(ch4_rxmldchainreq_m),
.ch0_rxmlfinealignreq(ch4_rxmlfinealignreq_m),
.ch0_rxoobreset(ch4_rxoobreset_m),
.ch0_rxpcsresetmask(ch4_rxpcsresetmask_m),
.ch0_rxpd(ch4_rxpd_m),
.ch0_rxphalignreq(ch4_rxphalignreq_m),
.ch0_rxphalignresetmask(ch4_rxphalignresetmask_m),
.ch0_rxphdlypd(ch4_rxphdlypd_m),
.ch0_rxphdlyreset(ch4_rxphdlyreset_m),
.ch0_rxphsetinitreq(ch4_rxphsetinitreq_m),
.ch0_rxphshift180(ch4_rxphshift180_m),
.ch0_rxpmaresetmask(ch4_rxpmaresetmask_m),
.ch0_rxpolarity(ch4_rxpolarity_m),
.ch0_rxprbscntreset(ch4_rxprbscntreset_m),
.ch0_rxprbssel(ch4_rxprbssel_m),
.ch0_rxprogdivreset(ch4_rxprogdivreset_m),
.ch0_rxrate(ch4_rxrate_m),
.ch0_rxresetmode(ch4_rxresetmode_m),
.ch0_rxslide(ch4_rxslide_m),
.ch0_rxsyncallin(ch4_rxsyncallin_m),
.ch0_rxtermination(ch4_rxtermination_m),
.ch0_rxuserrdy(ch4_rxuserrdy_m),
.ch0_rxusrclk(ch4_rxusrclk_m),
.ch0_rx10gstat(ch4_rx10gstat_m),
.ch0_rxbufstatus(ch4_rxbufstatus_m),
.ch0_rxbyteisaligned(ch4_rxbyteisaligned_m),
.ch0_rxbyterealign(ch4_rxbyterealign_m),
.ch0_rxcdrlock(ch4_rxcdrlock_m),
.ch0_rxcdrphdone(ch4_rxcdrphdone_m),
.ch0_rxchanbondseq(ch4_rxchanbondseq_m),
.ch0_rxchanisaligned(ch4_rxchanisaligned_m),
.ch0_rxchanrealign(ch4_rxchanrealign_m),
.ch0_rxchbondo(ch4_rxchbondo_m),
.ch0_rxclkcorcnt(ch4_rxclkcorcnt_m),
.ch0_rxcominitdet(ch4_rxcominitdet_m),
.ch0_rxcommadet(ch4_rxcommadet_m),
.ch0_rxcomsasdet(ch4_rxcomsasdet_m),
.ch0_rxcomwakedet(ch4_rxcomwakedet_m),
.ch0_rxctrl0(ch4_rxctrl0_m),
.ch0_rxctrl1(ch4_rxctrl1_m),
.ch0_rxctrl2(ch4_rxctrl2_m),
.ch0_rxctrl3(ch4_rxctrl3_m),
.ch0_rxdataextendrsvd(ch4_rxdataextendrsvd_m),
.ch0_rxdatavalid(ch4_rxdatavalid_m),
.ch0_rxdata(ch4_rxdata_m),
.ch0_rxdccdone(ch4_rxdccdone_m),
.ch0_rxdlyalignerr(ch4_rxdlyalignerr_m),
.ch0_rxdlyalignprog(ch4_rxdlyalignprog_m),
.ch0_rxelecidle(ch4_rxelecidle_m),
.ch0_rxfinealigndone(ch4_rxfinealigndone_m),
.ch0_rxheadervalid(ch4_rxheadervalid_m),
.ch0_rxheader(ch4_rxheader_m),
.ch0_rxosintdone(ch4_rxosintdone_m),
.ch0_rxosintstarted(ch4_rxosintstarted_m),
.ch0_rxosintstrobedone(ch4_rxosintstrobedone_m),
.ch0_rxosintstrobestarted(ch4_rxosintstrobestarted_m),
.ch0_rxoutclk(),
.ch0_txoutclk(),
.ch0_rxphaligndone(ch4_rxphaligndone_m),
.ch0_rxphalignerr(ch4_rxphalignerr_m),
.ch0_rxphdlyresetdone(ch4_rxphdlyresetdone_m),
.ch0_rxphsetinitdone(ch4_rxphsetinitdone_m),
.ch0_rxphshift180done(ch4_rxphshift180done_m),
.ch0_rxpmaresetdone(ch4_rxpmaresetdone_m),
.ch0_rxprbserr(ch4_rxprbserr_m),
.ch0_rxprbslocked(ch4_rxprbslocked_m),
.ch0_rxresetdone(ch4_rxresetdone_m),
.ch0_rxsliderdy(ch4_rxsliderdy_m),
.ch0_rxstartofseq(ch4_rxstartofseq_m),
.ch0_rxstatus(ch4_rxstatus_m),
.ch0_rxsyncdone(ch4_rxsyncdone_m),
.ch0_rxvalid(ch4_rxvalid_m),
.ch0_txcomsas(ch4_txcomsas_m),
.ch0_txcomwake(ch4_txcomwake_m),
.ch0_txctrl0(ch4_txctrl0_m),
.ch0_txctrl1(ch4_txctrl1_m),
.ch0_txctrl2(ch4_txctrl2_m),
.ch0_txdapicodeovrden(ch4_txdapicodeovrden_m),
.ch0_txdapicodereset(ch4_txdapicodereset_m),
.ch0_txdataextendrsvd(ch4_txdataextendrsvd_m),
.ch0_txdata(ch4_txdata_m),
.ch0_txdeemph(ch4_txdeemph_m),
.ch0_txdetectrx(ch4_txdetectrx_m),
.ch0_txdiffctrl(ch4_txdiffctrl_m),
.ch0_txdlyalignreq(ch4_txdlyalignreq_m),
.ch0_txelecidle(ch4_txelecidle_m),
.ch0_txheader(ch4_txheader_m),
.ch0_txinhibit(ch4_txinhibit_m),
.ch0_txlatclk(ch4_txlatclk_m),
.ch0_txmaincursor(ch4_txmaincursor_m),
.ch0_txmargin(ch4_txmargin_m),
.ch0_txmldchaindone(ch4_txmldchaindone_m),
.ch0_txmldchainreq(ch4_txmldchainreq_m),
.ch0_txoneszeros(ch4_txoneszeros_m),
.ch0_txpausedelayalign(ch4_txpausedelayalign_m),
.ch0_txpcsresetmask(ch4_txpcsresetmask_m),
.ch0_txpd(ch4_txpd_m),
.ch0_txphalignreq(ch4_txphalignreq_m),
.ch0_txphalignresetmask(ch4_txphalignresetmask_m),
.ch0_txphdlypd(ch4_txphdlypd_m),
.ch0_txphdlyreset(ch4_txphdlyreset_m),
.ch0_txphdlytstclk(ch4_txphdlytstclk_m),
.ch0_txphsetinitreq(ch4_txphsetinitreq_m),
.ch0_txphshift180(ch4_txphshift180_m),
.ch0_txpicodeovrden(ch4_txpicodeovrden_m),
.ch0_txpicodereset(ch4_txpicodereset_m),
.ch0_txpippmen(ch4_txpippmen_m),
.ch0_txpippmstepsize(ch4_txpippmstepsize_m),
.ch0_txpisopd(ch4_txpisopd_m),
.ch0_txpmaresetmask(ch4_txpmaresetmask_m),
.ch0_txpolarity(ch4_txpolarity_m),
.ch0_txpostcursor(ch4_txpostcursor_m),
.ch0_txprbsforceerr(ch4_txprbsforceerr_m),
.ch0_txprbssel(ch4_txprbssel_m),
.ch0_txprecursor(ch4_txprecursor_m),
.ch0_txprogdivreset(ch4_txprogdivreset_m),
.ch0_txrate(ch4_txrate_m),
.ch0_txresetmode(ch4_txresetmode_m),
.ch0_txsequence(ch4_txsequence_m),
.ch0_txswing(ch4_txswing_m),
.ch0_txuserrdy(ch4_txuserrdy_m),
.ch0_txusrclk(ch4_txusrclk_m),
.ch0_tx10gstat(ch4_tx10gstat_m),
.ch0_txbufstatus(ch4_txbufstatus_m),
.ch0_txcomfinish(ch4_txcomfinish_m),
.ch0_txdccdone(ch4_txdccdone_m),
.ch0_txdlyalignerr(ch4_txdlyalignerr_m),
.ch0_txdlyalignprog(ch4_txdlyalignprog_m),
.ch0_txphaligndone(ch4_txphaligndone_m),
.ch0_txphalignerr(ch4_txphalignerr_m),
.ch0_txphalignoutrsvd(ch4_txphalignoutrsvd_m),
.ch0_txphdlyresetdone(ch4_txphdlyresetdone_m),
.ch0_txphshift180done(ch4_txphshift180done_m),
.ch0_txpmaresetdone(ch4_txpmaresetdone_m),
.ch0_txresetdone(ch4_txresetdone_m),
.ch0_txsyncdone(ch4_txsyncdone_m),
.ch0_gttxreset(ch4_gttxreset_m),
.ch0_txcominit(ch4_txcominit_m),
.ch0_txphsetinitdone(ch4_txphsetinitdone_m),
.ch0_txprogdivresetdone(ch4_txprogdivresetdone_m),
.ch0_txsyncallin(ch4_txsyncallin_m),
.ch1_iloreset(ch5_iloreset_m),
.ch1_pcierstb(ch5_pcierstb_m),
.ch1_iloresetdone(ch5_iloresetdone_m),
.ch1_phystatus(ch5_phystatus_m),
.ch1_rxcdrhold(ch5_rxcdrhold_m),
.ch1_rxcdrovrden(ch5_rxcdrovrden_m),
.ch1_rxcdrreset(ch5_rxcdrreset_m),
.ch1_rxchbondi(ch5_rxchbondi_m),
.ch1_rxdapicodeovrden(ch5_rxdapicodeovrden_m),
.ch1_rxdapicodereset(ch5_rxdapicodereset_m),
.ch1_rxdlyalignreq(ch5_rxdlyalignreq_m),
.ch1_rxeqtraining(ch5_rxeqtraining_m),
.ch1_rxgearboxslip(ch5_rxgearboxslip_m),
.ch1_rxlatclk(ch5_rxlatclk_m),
.ch1_rxlpmen(ch5_rxlpmen_m),
.ch1_rxmldchaindone(ch5_rxmldchaindone_m),
.ch1_rxmldchainreq(ch5_rxmldchainreq_m),
.ch1_rxmlfinealignreq(ch5_rxmlfinealignreq_m),
.ch1_rxoobreset(ch5_rxoobreset_m),
.ch1_rxpcsresetmask(ch5_rxpcsresetmask_m),
.ch1_rxpd(ch5_rxpd_m),
.ch1_rxphalignreq(ch5_rxphalignreq_m),
.ch1_rxphalignresetmask(ch5_rxphalignresetmask_m),
.ch1_rxphdlypd(ch5_rxphdlypd_m),
.ch1_rxphdlyreset(ch5_rxphdlyreset_m),
.ch1_rxphsetinitreq(ch5_rxphsetinitreq_m),
.ch1_rxphshift180(ch5_rxphshift180_m),
.ch1_rxpmaresetmask(ch5_rxpmaresetmask_m),
.ch1_rxpolarity(ch5_rxpolarity_m),
.ch1_rxprbscntreset(ch5_rxprbscntreset_m),
.ch1_rxprbssel(ch5_rxprbssel_m),
.ch1_rxprogdivreset(ch5_rxprogdivreset_m),
.ch1_rxrate(ch5_rxrate_m),
.ch1_rxresetmode(ch5_rxresetmode_m),
.ch1_rxslide(ch5_rxslide_m),
.ch1_rxsyncallin(ch5_rxsyncallin_m),
.ch1_rxtermination(ch5_rxtermination_m),
.ch1_rxuserrdy(ch5_rxuserrdy_m),
.ch1_rxusrclk(ch5_rxusrclk_m),
.ch1_rx10gstat(ch5_rx10gstat_m),
.ch1_rxbufstatus(ch5_rxbufstatus_m),
.ch1_rxbyteisaligned(ch5_rxbyteisaligned_m),
.ch1_rxbyterealign(ch5_rxbyterealign_m),
.ch1_rxcdrlock(ch5_rxcdrlock_m),
.ch1_rxcdrphdone(ch5_rxcdrphdone_m),
.ch1_rxchanbondseq(ch5_rxchanbondseq_m),
.ch1_rxchanisaligned(ch5_rxchanisaligned_m),
.ch1_rxchanrealign(ch5_rxchanrealign_m),
.ch1_rxchbondo(ch5_rxchbondo_m),
.ch1_rxclkcorcnt(ch5_rxclkcorcnt_m),
.ch1_rxcominitdet(ch5_rxcominitdet_m),
.ch1_rxcommadet(ch5_rxcommadet_m),
.ch1_rxcomsasdet(ch5_rxcomsasdet_m),
.ch1_rxcomwakedet(ch5_rxcomwakedet_m),
.ch1_rxctrl0(ch5_rxctrl0_m),
.ch1_rxctrl1(ch5_rxctrl1_m),
.ch1_rxctrl2(ch5_rxctrl2_m),
.ch1_rxctrl3(ch5_rxctrl3_m),
.ch1_rxdataextendrsvd(ch5_rxdataextendrsvd_m),
.ch1_rxdatavalid(ch5_rxdatavalid_m),
.ch1_rxdata(ch5_rxdata_m),
.ch1_rxdccdone(ch5_rxdccdone_m),
.ch1_rxdlyalignerr(ch5_rxdlyalignerr_m),
.ch1_rxdlyalignprog(ch5_rxdlyalignprog_m),
.ch1_rxelecidle(ch5_rxelecidle_m),
.ch1_rxfinealigndone(ch5_rxfinealigndone_m),
.ch1_rxheadervalid(ch5_rxheadervalid_m),
.ch1_rxheader(ch5_rxheader_m),
.ch1_rxosintdone(ch5_rxosintdone_m),
.ch1_rxosintstarted(ch5_rxosintstarted_m),
.ch1_rxosintstrobedone(ch5_rxosintstrobedone_m),
.ch1_rxosintstrobestarted(ch5_rxosintstrobestarted_m),
.ch1_rxphaligndone(ch5_rxphaligndone_m),
.ch1_rxphalignerr(ch5_rxphalignerr_m),
.ch1_rxphdlyresetdone(ch5_rxphdlyresetdone_m),
.ch1_rxphsetinitdone(ch5_rxphsetinitdone_m),
.ch1_rxphshift180done(ch5_rxphshift180done_m),
.ch1_rxpmaresetdone(ch5_rxpmaresetdone_m),
.ch1_rxprbserr(ch5_rxprbserr_m),
.ch1_rxprbslocked(ch5_rxprbslocked_m),
.ch1_rxresetdone(ch5_rxresetdone_m),
.ch1_rxsliderdy(ch5_rxsliderdy_m),
.ch1_rxstartofseq(ch5_rxstartofseq_m),
.ch1_rxstatus(ch5_rxstatus_m),
.ch1_rxsyncdone(ch5_rxsyncdone_m),
.ch1_rxvalid(ch5_rxvalid_m),
.ch1_txcomsas(ch5_txcomsas_m),
.ch1_txcomwake(ch5_txcomwake_m),
.ch1_txctrl0(ch5_txctrl0_m),
.ch1_txctrl1(ch5_txctrl1_m),
.ch1_txctrl2(ch5_txctrl2_m),
.ch1_txdapicodeovrden(ch5_txdapicodeovrden_m),
.ch1_txdapicodereset(ch5_txdapicodereset_m),
.ch1_txdataextendrsvd(ch5_txdataextendrsvd_m),
.ch1_txdata(ch5_txdata_m),
.ch1_txdeemph(ch5_txdeemph_m),
.ch1_txdetectrx(ch5_txdetectrx_m),
.ch1_txdiffctrl(ch5_txdiffctrl_m),
.ch1_txdlyalignreq(ch5_txdlyalignreq_m),
.ch1_txelecidle(ch5_txelecidle_m),
.ch1_txheader(ch5_txheader_m),
.ch1_txinhibit(ch5_txinhibit_m),
.ch1_txlatclk(ch5_txlatclk_m),
.ch1_txmaincursor(ch5_txmaincursor_m),
.ch1_txmargin(ch5_txmargin_m),
.ch1_txmldchaindone(ch5_txmldchaindone_m),
.ch1_txmldchainreq(ch5_txmldchainreq_m),
.ch1_txoneszeros(ch5_txoneszeros_m),
.ch1_txpausedelayalign(ch5_txpausedelayalign_m),
.ch1_txpcsresetmask(ch5_txpcsresetmask_m),
.ch1_txpd(ch5_txpd_m),
.ch1_txphalignreq(ch5_txphalignreq_m),
.ch1_txphalignresetmask(ch5_txphalignresetmask_m),
.ch1_txphdlypd(ch5_txphdlypd_m),
.ch1_txphdlyreset(ch5_txphdlyreset_m),
.ch1_txphdlytstclk(ch5_txphdlytstclk_m),
.ch1_txphsetinitreq(ch5_txphsetinitreq_m),
.ch1_txphshift180(ch5_txphshift180_m),
.ch1_txpicodeovrden(ch5_txpicodeovrden_m),
.ch1_txpicodereset(ch5_txpicodereset_m),
.ch1_txpippmen(ch5_txpippmen_m),
.ch1_txpippmstepsize(ch5_txpippmstepsize_m),
.ch1_txpisopd(ch5_txpisopd_m),
.ch1_txpmaresetmask(ch5_txpmaresetmask_m),
.ch1_txpolarity(ch5_txpolarity_m),
.ch1_txpostcursor(ch5_txpostcursor_m),
.ch1_txprbsforceerr(ch5_txprbsforceerr_m),
.ch1_txprbssel(ch5_txprbssel_m),
.ch1_txprecursor(ch5_txprecursor_m),
.ch1_txprogdivreset(ch5_txprogdivreset_m),
.ch1_txrate(ch5_txrate_m),
.ch1_txresetmode(ch5_txresetmode_m),
.ch1_txsequence(ch5_txsequence_m),
.ch1_txswing(ch5_txswing_m),
.ch1_txsyncallin(ch5_txsyncallin_m),
.ch1_txuserrdy(ch5_txuserrdy_m),
.ch1_txusrclk(ch5_txusrclk_m),
.ch1_tx10gstat(ch5_tx10gstat_m),
.ch1_txbufstatus(ch5_txbufstatus_m),
.ch1_txcomfinish(ch5_txcomfinish_m),
.ch1_txdccdone(ch5_txdccdone_m),
.ch1_txdlyalignerr(ch5_txdlyalignerr_m),
.ch1_txdlyalignprog(ch5_txdlyalignprog_m),
.ch1_txphaligndone(ch5_txphaligndone_m),
.ch1_txphalignerr(ch5_txphalignerr_m),
.ch1_txphalignoutrsvd(ch5_txphalignoutrsvd_m),
.ch1_txphdlyresetdone(ch5_txphdlyresetdone_m),
.ch1_txphshift180done(ch5_txphshift180done_m),
.ch1_txpmaresetdone(ch5_txpmaresetdone_m),
.ch1_txresetdone(ch5_txresetdone_m),
.ch1_txsyncdone(ch5_txsyncdone_m),
.ch1_gttxreset(ch5_gttxreset_m),
.ch1_txcominit(ch5_txcominit_m),
.ch1_txphsetinitdone(ch5_txphsetinitdone_m),
.ch1_txprogdivresetdone(ch5_txprogdivresetdone_m),
.ch2_iloreset(ch6_iloreset_m),
.ch2_pcierstb(ch6_pcierstb_m),
.ch2_iloresetdone(ch6_iloresetdone_m),
.ch2_phystatus(ch6_phystatus_m),
.ch2_rxcdrhold(ch6_rxcdrhold_m),
.ch2_rxcdrovrden(ch6_rxcdrovrden_m),
.ch2_rxcdrreset(ch6_rxcdrreset_m),
.ch2_rxchbondi(ch6_rxchbondi_m),
.ch2_rxdapicodeovrden(ch6_rxdapicodeovrden_m),
.ch2_rxdapicodereset(ch6_rxdapicodereset_m),
.ch2_rxdlyalignreq(ch6_rxdlyalignreq_m),
.ch2_rxeqtraining(ch6_rxeqtraining_m),
.ch2_rxgearboxslip(ch6_rxgearboxslip_m),
.ch2_rxlatclk(ch6_rxlatclk_m),
.ch2_rxlpmen(ch6_rxlpmen_m),
.ch2_rxmldchaindone(ch6_rxmldchaindone_m),
.ch2_rxmldchainreq(ch6_rxmldchainreq_m),
.ch2_rxmlfinealignreq(ch6_rxmlfinealignreq_m),
.ch2_rxoobreset(ch6_rxoobreset_m),
.ch2_rxpcsresetmask(ch6_rxpcsresetmask_m),
.ch2_rxpd(ch6_rxpd_m),
.ch2_rxphalignreq(ch6_rxphalignreq_m),
.ch2_rxphalignresetmask(ch6_rxphalignresetmask_m),
.ch2_rxphdlypd(ch6_rxphdlypd_m),
.ch2_rxphdlyreset(ch6_rxphdlyreset_m),
.ch2_rxphsetinitreq(ch6_rxphsetinitreq_m),
.ch2_rxphshift180(ch6_rxphshift180_m),
.ch2_rxpmaresetmask(ch6_rxpmaresetmask_m),
.ch2_rxpolarity(ch6_rxpolarity_m),
.ch2_rxprbscntreset(ch6_rxprbscntreset_m),
.ch2_rxprbssel(ch6_rxprbssel_m),
.ch2_rxprogdivreset(ch6_rxprogdivreset_m),
.ch2_rxrate(ch6_rxrate_m),
.ch2_rxresetmode(ch6_rxresetmode_m),
.ch2_rxslide(ch6_rxslide_m),
.ch2_rxsyncallin(ch6_rxsyncallin_m),
.ch2_rxtermination(ch6_rxtermination_m),
.ch2_rxuserrdy(ch6_rxuserrdy_m),
.ch2_rxusrclk(ch6_rxusrclk_m),
.ch2_rx10gstat(ch6_rx10gstat_m),
.ch2_rxbufstatus(ch6_rxbufstatus_m),
.ch2_rxbyteisaligned(ch6_rxbyteisaligned_m),
.ch2_rxbyterealign(ch6_rxbyterealign_m),
.ch2_rxcdrlock(ch6_rxcdrlock_m),
.ch2_rxcdrphdone(ch6_rxcdrphdone_m),
.ch2_rxchanbondseq(ch6_rxchanbondseq_m),
.ch2_rxchanisaligned(ch6_rxchanisaligned_m),
.ch2_rxchanrealign(ch6_rxchanrealign_m),
.ch2_rxchbondo(ch6_rxchbondo_m),
.ch2_rxclkcorcnt(ch6_rxclkcorcnt_m),
.ch2_rxcominitdet(ch6_rxcominitdet_m),
.ch2_rxcommadet(ch6_rxcommadet_m),
.ch2_rxcomsasdet(ch6_rxcomsasdet_m),
.ch2_rxcomwakedet(ch6_rxcomwakedet_m),
.ch2_rxctrl0(ch6_rxctrl0_m),
.ch2_rxctrl1(ch6_rxctrl1_m),
.ch2_rxctrl2(ch6_rxctrl2_m),
.ch2_rxctrl3(ch6_rxctrl3_m),
.ch2_rxdataextendrsvd(ch6_rxdataextendrsvd_m),
.ch2_rxdatavalid(ch6_rxdatavalid_m),
.ch2_rxdata(ch6_rxdata_m),
.ch2_rxdccdone(ch6_rxdccdone_m),
.ch2_rxdlyalignerr(ch6_rxdlyalignerr_m),
.ch2_rxdlyalignprog(ch6_rxdlyalignprog_m),
.ch2_rxelecidle(ch6_rxelecidle_m),
.ch2_rxfinealigndone(ch6_rxfinealigndone_m),
.ch2_rxheadervalid(ch6_rxheadervalid_m),
.ch2_rxheader(ch6_rxheader_m),
.ch2_rxosintdone(ch6_rxosintdone_m),
.ch2_rxosintstarted(ch6_rxosintstarted_m),
.ch2_rxosintstrobedone(ch6_rxosintstrobedone_m),
.ch2_rxosintstrobestarted(ch6_rxosintstrobestarted_m),
.ch2_rxphaligndone(ch6_rxphaligndone_m),
.ch2_rxphalignerr(ch6_rxphalignerr_m),
.ch2_rxphdlyresetdone(ch6_rxphdlyresetdone_m),
.ch2_rxphsetinitdone(ch6_rxphsetinitdone_m),
.ch2_rxphshift180done(ch6_rxphshift180done_m),
.ch2_rxpmaresetdone(ch6_rxpmaresetdone_m),
.ch2_rxprbserr(ch6_rxprbserr_m),
.ch2_rxprbslocked(ch6_rxprbslocked_m),
.ch2_rxresetdone(ch6_rxresetdone_m),
.ch2_rxsliderdy(ch6_rxsliderdy_m),
.ch2_rxstartofseq(ch6_rxstartofseq_m),
.ch2_rxstatus(ch6_rxstatus_m),
.ch2_rxsyncdone(ch6_rxsyncdone_m),
.ch2_rxvalid(ch6_rxvalid_m),
.ch2_txcomsas(ch6_txcomsas_m),
.ch2_txcomwake(ch6_txcomwake_m),
.ch2_txctrl0(ch6_txctrl0_m),
.ch2_txctrl1(ch6_txctrl1_m),
.ch2_txctrl2(ch6_txctrl2_m),
.ch2_txdapicodeovrden(ch6_txdapicodeovrden_m),
.ch2_txdapicodereset(ch6_txdapicodereset_m),
.ch2_txdataextendrsvd(ch6_txdataextendrsvd_m),
.ch2_txdata(ch6_txdata_m),
.ch2_txdeemph(ch6_txdeemph_m),
.ch2_txdetectrx(ch6_txdetectrx_m),
.ch2_txdiffctrl(ch6_txdiffctrl_m),
.ch2_txdlyalignreq(ch6_txdlyalignreq_m),
.ch2_txelecidle(ch6_txelecidle_m),
.ch2_txheader(ch6_txheader_m),
.ch2_txinhibit(ch6_txinhibit_m),
.ch2_txlatclk(ch6_txlatclk_m),
.ch2_txmaincursor(ch6_txmaincursor_m),
.ch2_txmargin(ch6_txmargin_m),
.ch2_txmldchaindone(ch6_txmldchaindone_m),
.ch2_txmldchainreq(ch6_txmldchainreq_m),
.ch2_txoneszeros(ch6_txoneszeros_m),
.ch2_txpausedelayalign(ch6_txpausedelayalign_m),
.ch2_txpcsresetmask(ch6_txpcsresetmask_m),
.ch2_txpd(ch6_txpd_m),
.ch2_txphalignreq(ch6_txphalignreq_m),
.ch2_txphalignresetmask(ch6_txphalignresetmask_m),
.ch2_txphdlypd(ch6_txphdlypd_m),
.ch2_txphdlyreset(ch6_txphdlyreset_m),
.ch2_txphdlytstclk(ch6_txphdlytstclk_m),
.ch2_txphsetinitreq(ch6_txphsetinitreq_m),
.ch2_txphshift180(ch6_txphshift180_m),
.ch2_txpicodeovrden(ch6_txpicodeovrden_m),
.ch2_txpicodereset(ch6_txpicodereset_m),
.ch2_txpippmen(ch6_txpippmen_m),
.ch2_txpippmstepsize(ch6_txpippmstepsize_m),
.ch2_txpisopd(ch6_txpisopd_m),
.ch2_txpmaresetmask(ch6_txpmaresetmask_m),
.ch2_txpolarity(ch6_txpolarity_m),
.ch2_txpostcursor(ch6_txpostcursor_m),
.ch2_txprbsforceerr(ch6_txprbsforceerr_m),
.ch2_txprbssel(ch6_txprbssel_m),
.ch2_txprecursor(ch6_txprecursor_m),
.ch2_txprogdivreset(ch6_txprogdivreset_m),
.ch2_txrate(ch6_txrate_m),
.ch2_txresetmode(ch6_txresetmode_m),
.ch2_txsequence(ch6_txsequence_m),
.ch2_txswing(ch6_txswing_m),
.ch2_txsyncallin(ch6_txsyncallin_m),
.ch2_txuserrdy(ch6_txuserrdy_m),
.ch2_txusrclk(ch6_txusrclk_m),
.ch2_tx10gstat(ch6_tx10gstat_m),
.ch2_txbufstatus(ch6_txbufstatus_m),
.ch2_txcomfinish(ch6_txcomfinish_m),
.ch2_txdccdone(ch6_txdccdone_m),
.ch2_txdlyalignerr(ch6_txdlyalignerr_m),
.ch2_txdlyalignprog(ch6_txdlyalignprog_m),
.ch2_txphaligndone(ch6_txphaligndone_m),
.ch2_txphalignerr(ch6_txphalignerr_m),
.ch2_txphalignoutrsvd(ch6_txphalignoutrsvd_m),
.ch2_txphdlyresetdone(ch6_txphdlyresetdone_m),
.ch2_txphshift180done(ch6_txphshift180done_m),
.ch2_txpmaresetdone(ch6_txpmaresetdone_m),
.ch2_txresetdone(ch6_txresetdone_m),
.ch2_txsyncdone(ch6_txsyncdone_m),
.ch2_gttxreset(ch6_gttxreset_m),
.ch2_txcominit(ch6_txcominit_m),
.ch2_txphsetinitdone(ch6_txphsetinitdone_m),
.ch2_txprogdivresetdone(ch6_txprogdivresetdone_m),
.ch3_iloreset(ch7_iloreset_m),
.ch3_pcierstb(ch7_pcierstb_m),
.ch3_iloresetdone(ch7_iloresetdone_m),
.ch3_phystatus(ch7_phystatus_m),
.ch3_rxcdrhold(ch7_rxcdrhold_m),
.ch3_rxcdrovrden(ch7_rxcdrovrden_m),
.ch3_rxcdrreset(ch7_rxcdrreset_m),
.ch3_rxchbondi(ch7_rxchbondi_m),
.ch3_rxdapicodeovrden(ch7_rxdapicodeovrden_m),
.ch3_rxdapicodereset(ch7_rxdapicodereset_m),
.ch3_rxdlyalignreq(ch7_rxdlyalignreq_m),
.ch3_rxeqtraining(ch7_rxeqtraining_m),
.ch3_rxgearboxslip(ch7_rxgearboxslip_m),
.ch3_rxlatclk(ch7_rxlatclk_m),
.ch3_rxlpmen(ch7_rxlpmen_m),
.ch3_rxmldchaindone(ch7_rxmldchaindone_m),
.ch3_rxmldchainreq(ch7_rxmldchainreq_m),
.ch3_rxmlfinealignreq(ch7_rxmlfinealignreq_m),
.ch3_rxoobreset(ch7_rxoobreset_m),
.ch3_rxpcsresetmask(ch7_rxpcsresetmask_m),
.ch3_rxpd(ch7_rxpd_m),
.ch3_rxphalignreq(ch7_rxphalignreq_m),
.ch3_rxphalignresetmask(ch7_rxphalignresetmask_m),
.ch3_rxphdlypd(ch7_rxphdlypd_m),
.ch3_rxphdlyreset(ch7_rxphdlyreset_m),
.ch3_rxphsetinitreq(ch7_rxphsetinitreq_m),
.ch3_rxphshift180(ch7_rxphshift180_m),
.ch3_rxpmaresetmask(ch7_rxpmaresetmask_m),
.ch3_rxpolarity(ch7_rxpolarity_m),
.ch3_rxprbscntreset(ch7_rxprbscntreset_m),
.ch3_rxprbssel(ch7_rxprbssel_m),
.ch3_rxprogdivreset(ch7_rxprogdivreset_m),
.ch3_rxrate(ch7_rxrate_m),
.ch3_rxresetmode(ch7_rxresetmode_m),
.ch3_rxslide(ch7_rxslide_m),
.ch3_rxsyncallin(ch7_rxsyncallin_m),
.ch3_rxtermination(ch7_rxtermination_m),
.ch3_rxuserrdy(ch7_rxuserrdy_m),
.ch3_rxusrclk(ch7_rxusrclk_m),
.ch3_rx10gstat(ch7_rx10gstat_m),
.ch3_rxbufstatus(ch7_rxbufstatus_m),
.ch3_rxbyteisaligned(ch7_rxbyteisaligned_m),
.ch3_rxbyterealign(ch7_rxbyterealign_m),
.ch3_rxcdrlock(ch7_rxcdrlock_m),
.ch3_rxcdrphdone(ch7_rxcdrphdone_m),
.ch3_rxchanbondseq(ch7_rxchanbondseq_m),
.ch3_rxchanisaligned(ch7_rxchanisaligned_m),
.ch3_rxchanrealign(ch7_rxchanrealign_m),
.ch3_rxchbondo(ch7_rxchbondo_m),
.ch3_rxclkcorcnt(ch7_rxclkcorcnt_m),
.ch3_rxcominitdet(ch7_rxcominitdet_m),
.ch3_rxcommadet(ch7_rxcommadet_m),
.ch3_rxcomsasdet(ch7_rxcomsasdet_m),
.ch3_rxcomwakedet(ch7_rxcomwakedet_m),
.ch3_rxctrl0(ch7_rxctrl0_m),
.ch3_rxctrl1(ch7_rxctrl1_m),
.ch3_rxctrl2(ch7_rxctrl2_m),
.ch3_rxctrl3(ch7_rxctrl3_m),
.ch3_rxdataextendrsvd(ch7_rxdataextendrsvd_m),
.ch3_rxdatavalid(ch7_rxdatavalid_m),
.ch3_rxdata(ch7_rxdata_m),
.ch3_rxdccdone(ch7_rxdccdone_m),
.ch3_rxdlyalignerr(ch7_rxdlyalignerr_m),
.ch3_rxdlyalignprog(ch7_rxdlyalignprog_m),
.ch3_rxelecidle(ch7_rxelecidle_m),
.ch3_rxfinealigndone(ch7_rxfinealigndone_m),
.ch3_rxheadervalid(ch7_rxheadervalid_m),
.ch3_rxheader(ch7_rxheader_m),
.ch3_rxosintdone(ch7_rxosintdone_m),
.ch3_rxosintstarted(ch7_rxosintstarted_m),
.ch3_rxosintstrobedone(ch7_rxosintstrobedone_m),
.ch3_rxosintstrobestarted(ch7_rxosintstrobestarted_m),
.ch3_rxphaligndone(ch7_rxphaligndone_m),
.ch3_rxphalignerr(ch7_rxphalignerr_m),
.ch3_rxphdlyresetdone(ch7_rxphdlyresetdone_m),
.ch3_rxphsetinitdone(ch7_rxphsetinitdone_m),
.ch3_rxphshift180done(ch7_rxphshift180done_m),
.ch3_rxpmaresetdone(ch7_rxpmaresetdone_m),
.ch3_rxprbserr(ch7_rxprbserr_m),
.ch3_rxprbslocked(ch7_rxprbslocked_m),
.ch3_rxresetdone(ch7_rxresetdone_m),
.ch3_rxsliderdy(ch7_rxsliderdy_m),
.ch3_rxstartofseq(ch7_rxstartofseq_m),
.ch3_rxstatus(ch7_rxstatus_m),
.ch3_rxsyncdone(ch7_rxsyncdone_m),
.ch3_rxvalid(ch7_rxvalid_m),
.ch3_txcomsas(ch7_txcomsas_m),
.ch3_txcomwake(ch7_txcomwake_m),
.ch3_txctrl0(ch7_txctrl0_m),
.ch3_txctrl1(ch7_txctrl1_m),
.ch3_txctrl2(ch7_txctrl2_m),
.ch3_txdapicodeovrden(ch7_txdapicodeovrden_m),
.ch3_txdapicodereset(ch7_txdapicodereset_m),
.ch3_txdataextendrsvd(ch7_txdataextendrsvd_m),
.ch3_txdata(ch7_txdata_m),
.ch3_txdeemph(ch7_txdeemph_m),
.ch3_txdetectrx(ch7_txdetectrx_m),
.ch3_txdiffctrl(ch7_txdiffctrl_m),
.ch3_txdlyalignreq(ch7_txdlyalignreq_m),
.ch3_txelecidle(ch7_txelecidle_m),
.ch3_txheader(ch7_txheader_m),
.ch3_txinhibit(ch7_txinhibit_m),
.ch3_txlatclk(ch7_txlatclk_m),
.ch3_txmaincursor(ch7_txmaincursor_m),
.ch3_txmargin(ch7_txmargin_m),
.ch3_txmldchaindone(ch7_txmldchaindone_m),
.ch3_txmldchainreq(ch7_txmldchainreq_m),
.ch3_txoneszeros(ch7_txoneszeros_m),
.ch3_txpausedelayalign(ch7_txpausedelayalign_m),
.ch3_txpcsresetmask(ch7_txpcsresetmask_m),
.ch3_txpd(ch7_txpd_m),
.ch3_txphalignreq(ch7_txphalignreq_m),
.ch3_txphalignresetmask(ch7_txphalignresetmask_m),
.ch3_txphdlypd(ch7_txphdlypd_m),
.ch3_txphdlyreset(ch7_txphdlyreset_m),
.ch3_txphdlytstclk(ch7_txphdlytstclk_m),
.ch3_txphsetinitreq(ch7_txphsetinitreq_m),
.ch3_txphshift180(ch7_txphshift180_m),
.ch3_txpicodeovrden(ch7_txpicodeovrden_m),
.ch3_txpicodereset(ch7_txpicodereset_m),
.ch3_txpippmen(ch7_txpippmen_m),
.ch3_txpippmstepsize(ch7_txpippmstepsize_m),
.ch3_txpisopd(ch7_txpisopd_m),
.ch3_txpmaresetmask(ch7_txpmaresetmask_m),
.ch3_txpolarity(ch7_txpolarity_m),
.ch3_txpostcursor(ch7_txpostcursor_m),
.ch3_txprbsforceerr(ch7_txprbsforceerr_m),
.ch3_txprbssel(ch7_txprbssel_m),
.ch3_txprecursor(ch7_txprecursor_m),
.ch3_txprogdivreset(ch7_txprogdivreset_m),
.ch3_txrate(ch7_txrate_m),
.ch3_txresetmode(ch7_txresetmode_m),
.ch3_txsequence(ch7_txsequence_m),
.ch3_txswing(ch7_txswing_m),
.ch3_txsyncallin(ch7_txsyncallin_m),
.ch3_txuserrdy(ch7_txuserrdy_m),
.ch3_txusrclk(ch7_txusrclk_m),
.ch3_tx10gstat(ch7_tx10gstat_m),
.ch3_txbufstatus(ch7_txbufstatus_m),
.ch3_txcomfinish(ch7_txcomfinish_m),
.ch3_txdccdone(ch7_txdccdone_m),
.ch3_txdlyalignerr(ch7_txdlyalignerr_m),
.ch3_txdlyalignprog(ch7_txdlyalignprog_m),
.ch3_txphaligndone(ch7_txphaligndone_m),
.ch3_txphalignerr(ch7_txphalignerr_m),
.ch3_txphalignoutrsvd(ch7_txphalignoutrsvd_m),
.ch3_txphdlyresetdone(ch7_txphdlyresetdone_m),
.ch3_txphshift180done(ch7_txphshift180done_m),
.ch3_txpmaresetdone(ch7_txpmaresetdone_m),
.ch3_txresetdone(ch7_txresetdone_m),
.ch3_txsyncdone(ch7_txsyncdone_m),
.ch3_gttxreset(ch7_gttxreset_m),
.ch3_txcominit(ch7_txcominit_m),
.ch3_txphsetinitdone(ch7_txphsetinitdone_m),
.ch3_txprogdivresetdone(ch7_txprogdivresetdone_m),
.hsclk0_lcpllclkrsvd0(q1_hsclk0_lcpllclkrsvd0_m),
.hsclk0_lcpllclkrsvd1(q1_hsclk0_lcpllclkrsvd1_m),
.hsclk0_lcpllfbdiv(q1_hsclk0_lcpllfbdiv_m),
.hsclk0_lcpllpd(q1_hsclk0_lcpllpd_m),
.hsclk0_lcpllrefclksel(q1_hsclk0_lcpllrefclksel_m),
.hsclk0_lcpllresetbypassmode(q1_hsclk0_lcpllresetbypassmode_m),
.hsclk0_lcpllresetmask(q1_hsclk0_lcpllresetmask_m),
.hsclk0_lcpllreset(q1_hsclk0_lcpllreset_m),
.hsclk0_lcpllrsvd0(q1_hsclk0_lcpllrsvd0_m),
.hsclk0_lcpllrsvd1(q1_hsclk0_lcpllrsvd1_m),
.hsclk0_lcpllsdmdata(q1_hsclk0_lcpllsdmdata_m),
.hsclk0_lcpllsdmtoggle(q1_hsclk0_lcpllsdmtoggle_m),
.hsclk0_rpllclkrsvd0(q1_hsclk0_rpllclkrsvd0_m),
.hsclk0_rpllclkrsvd1(q1_hsclk0_rpllclkrsvd1_m),
.hsclk0_rpllfbdiv(q1_hsclk0_rpllfbdiv_m),
.hsclk0_rpllpd(q1_hsclk0_rpllpd_m),
.hsclk0_rpllrefclksel(q1_hsclk0_rpllrefclksel_m),
.hsclk0_rpllresetbypassmode(q1_hsclk0_rpllresetbypassmode_m),
.hsclk0_rpllresetmask(q1_hsclk0_rpllresetmask_m),
.hsclk0_rpllreset(q1_hsclk0_rpllreset_m),
.hsclk0_rpllrsvd0(q1_hsclk0_rpllrsvd0_m),
.hsclk0_rpllrsvd1(q1_hsclk0_rpllrsvd1_m),
.hsclk0_rpllsdmdata(q1_hsclk0_rpllsdmdata_m),
.hsclk0_rpllsdmtoggle(q1_hsclk0_rpllsdmtoggle_m),
.hsclk0_lcpllfbclklost(q1_hsclk0_lcpllfbclklost_m),
.hsclk0_lcpllrefclklost(q1_hsclk0_lcpllrefclklost_m),
.hsclk0_rpllfbclklost(q1_hsclk0_rpllfbclklost_m),
.hsclk0_rpllrefclklost(q1_hsclk0_rpllrefclklost_m),
.hsclk0_lcpllrefclkmonitor(q1_hsclk0_lcpllrefclkmonitor_m),
.hsclk0_rpllrefclkmonitor(q1_hsclk0_rpllrefclkmonitor_m),
.hsclk0_lcpllrsvdout(q1_hsclk0_lcpllrsvdout_m),
.hsclk0_rpllrsvdout(q1_hsclk0_rpllrsvdout_m),
.hsclk1_lcpllclkrsvd0(q1_hsclk1_lcpllclkrsvd0_m),
.hsclk1_lcpllclkrsvd1(q1_hsclk1_lcpllclkrsvd1_m),
.hsclk1_lcpllfbdiv(q1_hsclk1_lcpllfbdiv_m),
.hsclk1_lcpllpd(q1_hsclk1_lcpllpd_m),
.hsclk1_lcpllrefclksel(q1_hsclk1_lcpllrefclksel_m),
.hsclk1_lcpllresetbypassmode(q1_hsclk1_lcpllresetbypassmode_m),
.hsclk1_lcpllresetmask(q1_hsclk1_lcpllresetmask_m),
.hsclk1_lcpllreset(q1_hsclk1_lcpllreset_m),
.hsclk1_lcpllrsvd0(q1_hsclk1_lcpllrsvd0_m),
.hsclk1_lcpllrsvd1(q1_hsclk1_lcpllrsvd1_m),
.hsclk1_lcpllsdmdata(q1_hsclk1_lcpllsdmdata_m),
.hsclk1_lcpllsdmtoggle(q1_hsclk1_lcpllsdmtoggle_m),
.hsclk1_rpllclkrsvd0(q1_hsclk1_rpllclkrsvd0_m),
.hsclk1_rpllclkrsvd1(q1_hsclk1_rpllclkrsvd1_m),
.hsclk1_rpllfbdiv(q1_hsclk1_rpllfbdiv_m),
.hsclk1_rpllpd(q1_hsclk1_rpllpd_m),
.hsclk1_rpllrefclksel(q1_hsclk1_rpllrefclksel_m),
.hsclk1_rpllresetbypassmode(q1_hsclk1_rpllresetbypassmode_m),
.hsclk1_rpllresetmask(q1_hsclk1_rpllresetmask_m),
.hsclk1_rpllreset(q1_hsclk1_rpllreset_m),
.hsclk1_rpllrsvd0(q1_hsclk1_rpllrsvd0_m),
.hsclk1_rpllrsvd1(q1_hsclk1_rpllrsvd1_m),
.hsclk1_rpllsdmdata(q1_hsclk1_rpllsdmdata_m),
.hsclk1_rpllsdmtoggle(q1_hsclk1_rpllsdmtoggle_m),
.hsclk1_lcpllfbclklost(q1_hsclk1_lcpllfbclklost_m),
.hsclk1_lcpllrefclklost(q1_hsclk1_lcpllrefclklost_m),
.hsclk1_rpllfbclklost(q1_hsclk1_rpllfbclklost_m),
.hsclk1_rpllrefclklost(q1_hsclk1_rpllrefclklost_m),
.hsclk1_lcpllrefclkmonitor(q1_hsclk1_lcpllrefclkmonitor_m),
.hsclk1_rpllrefclkmonitor(q1_hsclk1_rpllrefclkmonitor_m),
.hsclk1_lcpllrsvdout(q1_hsclk1_lcpllrsvdout_m),
.hsclk1_rpllrsvdout(q1_hsclk1_rpllrsvdout_m),
.s0_axis_tready(m3_axis_tready_m),
.s0_axis_tdata(m3_axis_tdata_m),
.s0_axis_tlast(m3_axis_tlast_m),
.s0_axis_tvalid(m3_axis_tvalid_m),
.s1_axis_tready(m4_axis_tready_m),
.s1_axis_tdata(m4_axis_tdata_m),
.s1_axis_tlast(m4_axis_tlast_m),
.s1_axis_tvalid(m4_axis_tvalid_m),
.s2_axis_tready(m5_axis_tready_m),
.s2_axis_tdata(m5_axis_tdata_m),
.s2_axis_tlast(m5_axis_tlast_m),
.s2_axis_tvalid(m5_axis_tvalid_m),
.pcielinkreachtarget(q1_pcielinkreachtarget_m),
.pcieltssm(q1_pcieltssm_m),
.rxmarginclk(q1_rxmarginclk_m),
.rxmarginreqcmd(q1_rxmarginreqcmd_m),
.rxmarginreqlanenum(q1_rxmarginreqlanenum_m),
.rxmarginreqpayld(q1_rxmarginreqpayld_m),
.rxmarginreqreq(q1_rxmarginreqreq_m),
.rxmarginresack(q1_rxmarginresack_m),
.rxmarginresreq(q1_rxmarginresreq_m),
.rxmarginreqack(q1_rxmarginreqack_m),
.rxmarginrescmd(q1_rxmarginrescmd_m),
.rxmarginreslanenum(q1_rxmarginreslanenum_m),
.rxmarginrespayld(q1_rxmarginrespayld_m),
.m0_axis_tready(s3_axis_tready_m),
.m0_axis_tdata(s3_axis_tdata_m),
.m0_axis_tlast(s3_axis_tlast_m),
.m0_axis_tvalid(s3_axis_tvalid_m),
.m1_axis_tready(s4_axis_tready_m),
.m1_axis_tdata(s4_axis_tdata_m),
.m1_axis_tlast(s4_axis_tlast_m),
.m1_axis_tvalid(s4_axis_tvalid_m),
.m2_axis_tready(s5_axis_tready_m),
.m2_axis_tdata(s5_axis_tdata_m),
.m2_axis_tlast(s5_axis_tlast_m),
.m2_axis_tvalid(s5_axis_tvalid_m),
.gtpowergood(q1_gtpowergood_m),
.ch0_rxprogdivresetdone(ch4_rxprogdivresetdone_m),
.ch0_gtrxreset(ch4_gtrxreset_m),
.ch0_cdrbmcdrreq(ch4_cdrbmcdrreq_m),
.ch0_cdrfreqos(ch4_cdrfreqos_m),
.ch0_cdrincpctrl(ch4_cdrincpctrl_m),
.ch0_cdrstepdir(ch4_cdrstepdir_m),
.ch0_cdrstepsq(ch4_cdrstepsq_m),
.ch0_cdrstepsx(ch4_cdrstepsx_m),
.ch0_cfokovrdfinish(ch4_cfokovrdfinish_m),
.ch0_cfokovrdpulse(ch4_cfokovrdpulse_m),
.ch0_cfokovrdstart(ch4_cfokovrdstart_m),
.ch0_eyescanreset(ch4_eyescanreset_m),
.ch0_eyescantrigger(ch4_eyescantrigger_m),
.ch0_eyescandataerror(ch4_eyescandataerror_m),
.ch0_cfokovrdrdy0(ch4_cfokovrdrdy0_m),
.ch0_cfokovrdrdy1(ch4_cfokovrdrdy1_m),
.ch1_rxprogdivresetdone(ch5_rxprogdivresetdone_m),
.ch1_gtrxreset(ch5_gtrxreset_m),
.ch1_cdrbmcdrreq(ch5_cdrbmcdrreq_m),
.ch1_cdrfreqos(ch5_cdrfreqos_m),
.ch1_cdrincpctrl(ch5_cdrincpctrl_m),
.ch1_cdrstepdir(ch5_cdrstepdir_m),
.ch1_cdrstepsq(ch5_cdrstepsq_m),
.ch1_cdrstepsx(ch5_cdrstepsx_m),
.ch1_cfokovrdfinish(ch5_cfokovrdfinish_m),
.ch1_cfokovrdpulse(ch5_cfokovrdpulse_m),
.ch1_cfokovrdstart(ch5_cfokovrdstart_m),
.ch1_eyescanreset(ch5_eyescanreset_m),
.ch1_eyescantrigger(ch5_eyescantrigger_m),
.ch1_eyescandataerror(ch5_eyescandataerror_m),
.ch1_cfokovrdrdy0(ch5_cfokovrdrdy0_m),
.ch1_cfokovrdrdy1(ch5_cfokovrdrdy1_m),
.ch2_rxprogdivresetdone(ch6_rxprogdivresetdone_m),
.ch2_gtrxreset(ch6_gtrxreset_m),
.ch2_cdrbmcdrreq(ch6_cdrbmcdrreq_m),
.ch2_cdrfreqos(ch6_cdrfreqos_m),
.ch2_cdrincpctrl(ch6_cdrincpctrl_m),
.ch2_cdrstepdir(ch6_cdrstepdir_m),
.ch2_cdrstepsq(ch6_cdrstepsq_m),
.ch2_cdrstepsx(ch6_cdrstepsx_m),
.ch2_cfokovrdfinish(ch6_cfokovrdfinish_m),
.ch2_cfokovrdpulse(ch6_cfokovrdpulse_m),
.ch2_cfokovrdstart(ch6_cfokovrdstart_m),
.ch2_eyescanreset(ch6_eyescanreset_m),
.ch2_eyescantrigger(ch6_eyescantrigger_m),
.ch2_eyescandataerror(ch6_eyescandataerror_m),
.ch2_cfokovrdrdy0(ch6_cfokovrdrdy0_m),
.ch2_cfokovrdrdy1(ch6_cfokovrdrdy1_m),
.ch3_rxprogdivresetdone(ch7_rxprogdivresetdone_m),
.ch3_gtrxreset(ch7_gtrxreset_m),
.ch3_cdrbmcdrreq(ch7_cdrbmcdrreq_m),
.ch3_cdrfreqos(ch7_cdrfreqos_m),
.ch3_cdrincpctrl(ch7_cdrincpctrl_m),
.ch3_cdrstepdir(ch7_cdrstepdir_m),
.ch3_cdrstepsq(ch7_cdrstepsq_m),
.ch3_cdrstepsx(ch7_cdrstepsx_m),
.ch3_cfokovrdfinish(ch7_cfokovrdfinish_m),
.ch3_cfokovrdpulse(ch7_cfokovrdpulse_m),
.ch3_cfokovrdstart(ch7_cfokovrdstart_m),
.ch3_eyescanreset(ch7_eyescanreset_m),
.ch3_eyescantrigger(ch7_eyescantrigger_m),
.ch3_eyescandataerror(ch7_eyescandataerror_m),
.ch3_cfokovrdrdy0(ch7_cfokovrdrdy0_m),
.ch3_cfokovrdrdy1(ch7_cfokovrdrdy1_m),
.hsclk0_lcplllock(q1_hsclk0_lcplllock_m),
.hsclk0_rplllock(q1_hsclk0_rplllock_m),
.hsclk1_lcplllock(q1_hsclk1_lcplllock_m),
.hsclk1_rplllock(q1_hsclk1_rplllock_m),
.debugtraceready(q1_debugtracetready_m),
.ch0_txmstreset     (ch4_msttxreset_m),
.ch0_txmstresetdone (ch4_msttxresetdone_m),
.ch1_txmstreset     (ch5_msttxreset_m),
.ch1_txmstresetdone (ch5_msttxresetdone_m),
.ch2_txmstreset     (ch6_msttxreset_m),
.ch2_txmstresetdone (ch6_msttxresetdone_m),
.ch3_txmstreset     (ch7_msttxreset_m),
.ch3_txmstresetdone (ch7_msttxresetdone_m),
.ch0_rxmstreset      ( ch4_mstrxreset_m ),
.ch0_rxmstresetdone  ( ch4_mstrxresetdone_m),
.ch1_rxmstreset      ( ch5_mstrxreset_m),
.ch1_rxmstresetdone  ( ch5_mstrxresetdone_m),
.ch2_rxmstreset      ( ch6_mstrxreset_m),
.ch2_rxmstresetdone  ( ch6_mstrxresetdone_m),
.ch3_rxmstreset      ( ch7_mstrxreset_m),
.ch3_rxmstresetdone  ( ch7_mstrxresetdone_m),
.rxn(q1_gt_quad_base_serial_rxn),
.rxp(q1_gt_quad_base_serial_rxp),
.txn(q1_gt_quad_base_serial_txn),
.txp(q1_gt_quad_base_serial_txp),
.refclk0_gtrefclkpdint(q1_refclk0_gtrefclkpdint),
.pipenorthin(pipenorthoutq0_to_pipenorthinq1),
.resetdone_northin(resetdone_northout_q0_to_resetdone_northin_q1), 
.rxpinorthin(rxpinorthout_q0_to_rxpinorthin_q1), 
.txpinorthin(txpinorthout_q0_to_txpinorthin_q1), 
.pipesouthout( pipesouthin_q0_to_pipesouthout_q1),  
.resetdone_southout(resetdone_southin_q0_to_resetdone_southout_q1), 
.rxpisouthout(rxpisouthin_to_rxpsouthout_q1), 
.txpisouthout(txpisouthin_to_txpsouthout_q1)
