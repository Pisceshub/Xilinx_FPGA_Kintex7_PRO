`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16448)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEHcA42TsmOWkHd+n/5aa09U3CiYLGZjf5V9NYmJa0+VL5XX9cGnsX377
azdXTTjyZaopwVQ3kwkZvUHs8mHLTbD1EeNTp+nfmmkd1saNzXkFEEfyTfQJ/fuUsWD2yM4JgQzX
1kTMs2iA9qOFT7qgUA4PcnAL6jXWwAhAMEQU0sdUKR2VYIS9+j3YT+kNGYFhWBmoVqj4KFxAcZgw
NlyyinXuMdiwT7VdKlKuQBlPuUE4vq+RA3kS4WJXWrawGqfA8OzCWqmV04t7QgN2475cJMPwzAZa
ffN8m81DIYADncQrPufrKQnBPwVN7tt/Q7mUv0LGPG1YcG9YGaZ9FDPi8zLOdNOMJZfdmnpjgKJL
uuIVLOIgVQllKGafFYYfFHpdf9Qe/tqpCmRPbgsNC/eUg4FAXoRA3fYPJ2LdF8TBg/8IDc39r4rW
qtyMxUWjG/IMI5OI5CS3DfT7s6enbfncb23BCktRF3GzY2i7rwM9wCZuWA4NgIV8bNfjtCGbp34H
e4TDpNVCqggcQwZcbMQYQcjP1OccbodopFmSuCVff1t16ariK8FWYo0QKj+AP/4eiOynMegYcrmo
L2OyTr95W/Y+Dvwd5IkukWl2gDFYbtWLziTfsodD9gnsJxmvAmiaM+xm9Du6Skh1LaRFC34X/anv
5YnK4PGMZmQxCK8JOkk8ERQYES0zX3US3wdaYdJ7BDRfN4zn2wcDzt72epJhunMqZA7VBu4woHHT
V4Ya4G3Pj6MODsl8Te1Q3su42yJarkVt5yEuAw5yzSu0/zo6eAmSR4M/HfUbkS+l6O6gjwOk69Rk
qne4IE4Glz5KKAIrvgt65eBhYHwCBK14v3J+a0qslh+K+IwR01xz+PSZqf+I+p8Ujt2x8ZDzfj5n
PxIUa1kjAMt8YBy+QmJnt+TVGgdbJLrlpfzi321mMBY85LO3DY12XrcOyRpJCfFlN5TpmHJtplJA
M9cILVY1Ev6K7oZHqD+DYmLiMs2YyYH64sDsHcnw0SZTo4/Spwvb3yoxuJLz1Ua/ragMwklCOmyC
FTLPV646cPiNwz4rzWtU0lFWeKCBxV7+ZhbLjSmMp+/xqosjfwlqJcXGDndzCMcaRtbCOLXji46s
mkh7ee9F+gvaX7zeHo/IJ3iVzftdk0lUrUMlStJglh1Kf4yv3NZvOZUCXGMKU+tFdIZifCD7jDy/
B/R3d6+075nfsQn+QyujZdKe4T+Ltt3lg6DAnGkkPzhdh1CMeJos1Bi896X170eR3vY351Sqh7A2
5q4V5MMWazS8vu8rXYiGyRmUQ6N4MojBL9ITiwiIU4GJkz+bEBLkWPukLn0A9FsDhYTmxSyDVOvW
YUHCVv8vOSYF0gUeptr+HpLGJOpo8knBt+8iX9+1XEbQ+gcYbeyqF6cX8n+nvA65ERgw3O6ZqXoC
05y5qNLW1b8NlY2c6eyU2RPK7LB3mBmwmcyzSskUL8NG4WaOVX0SCOjLOvfIYqaOOA6vVvEwWa9/
iOGfm7oM3bt+qIUODkOZGQLGMGowUq9xAbu3pdrAOuiBmTU5CIRpBaYCcnPBuq3Dqf6cVshbgxmq
koVC2Wpz60dQnsuC+Gpu2ZO47ly4WLeebt/Ri05Gjaj2zDIKFt4XNg/wdOra/Moxna5G+H3uh3YW
Qs45MwcM7W25XfW2zPyBYvrNSRPehVsTzCcx/q8mUbr4bMN+jRrV8RU25ydHyWY79CNKMhSRPjRX
XCgsLK5+VbJbSQ4LvBRpVcKaAX34aevk9nox4UihKLlG4sru/dYV1hA3X49cl5gTTgyyecumCfk4
ZKW7SrmuNdfA5UhawqnhWtsDf4QeSWXfhYIwdYuuxQHowY1ZxDl0g2E2Lt7piQtCUHpzEoiOSG/Y
bWR7vzByh4dxs4jdqkMURZiseKyAZlSjB7Drs0hmd/pwkOwm0gGxuhs5ZHOJqiIZYQp4XAloM51a
v4KjcjTCsNoIjWGkd3rDElEX+OJzoaqlbUU8OvBpfuO6WCXybG1K3LPFWhHim5ua8dz/AIDvRKUY
1ZYAeIHwIlW5YKYzbFTvfUtEqudY1e0p7tpOc/j0iuKrg+SOIyx7qoaLpbKv2u7Mx1vL+7squ4EF
w1oXbeodF6PUAnX+vqqWhWFBf7RAPLEZ666bQNsEiqFTod8rMAsUizccaslcTr0Qe1r9++OhRR9Q
YFrcsZpm2c4ZsfsMIeerKIi9r0QBU4arS3pFmekyMv5CbGkmNUoEv4ynpr34gvuu+xGoaH3xry3T
JbjZ8SsSXG+YUKz9lQMcwGoiagFSR7ikYYlRZE7z82q1rDO/7SWeA/LfVJs8CbEzPwTQEPlM3j42
HUlqUTX7DE7qe4nhL5V6h7LsGMwFS+YqfytAtx/S2RSV+RXDSwpBTLVzT8ebNH2d46yJVgJ3Gkc2
WKigP3TcvNG0Z+VzL2IALLCm0tf8An2NBZZ+0vjNKdacf4NZaodlR6idsXbMJAbWJmQLex3ULT4B
muEMPaLXkMphiZI8q8jVjkU8p2eIgnn9wV2wwYXQDczk20uSUNT1O0dvLMO6lqir8JIbG+dPO5VQ
d9h2Hy9GDJI/Wm2sbUqiIPXOOFvdad8HkhPWIbqj9qAa8XEEfai4D0PmRgm4Rfd6DvIs3XE4Y61U
1sZgVS7xMbMfvVw/ZDLFuQxPcFsnXVGDbG0B9d6RAvqRAJ0KRtqd4Ui7jgl/5PK26621o2Y2c/cS
UHXQKzXJMD2L8Fxy8wraagmDKnm9hT4y6g26o5mYsWIvbp4uX9/HWQFyF1DX7ac9s0TLKzXWi/TB
NiT54At8qPFbCJXuD8YkCiApVnIe9TMl16/EF7YPJtQegOjg/D+Yd/jbErvaGStdbBs/ZAsRxCBx
1TnrrLdz4bthyJoVtzYbZO0Fgef6dGp+QorMxL30Sw7UoMAphdypfEY2RzWVX5k2vHXe6TfVzVJU
ufsQXhdWke+Kmp/bDpCmKsKE2gAnk1FRjeVoteWQcy0gfa0UBT09scWm8Z7IhmuOoDyGlJSobKrT
ct2Z16hI1GfgX7PTngwkrVrXgzEmLl72z69Bb3KNQBdfG15WlWPcuCYuoYNH2uP6zhCYeviv/WK7
kYEzWPloX9RjQQzQVOoNbhyniBVGY30CxpFqlLyX0y8QXnOOCy7ty8xWtzT8oYxxYTp7/kQVsZf5
P4hXhkKdxOv1UG6nleU6kyAwzyaE+HZXFH156faAL9s2uqzxZjijA62eh1UEfQeezIDc18JzSy5T
QgrJ0RCC21zJa58/x1HRSKaVMeVyLoQ7oajxwk6SU4LjO25JiU52VYgxBa+0nKQnT6T2fGe+zDNP
gaeqvk38qTjB91OLovxyplhqvMJRyVGoN9pLE4IR3dYjsdJVnrhIcsFODX5Fi+3yL8hsRNdlXcWk
R+8u7T0S/q+v3DSofiAv4ibghlOgd0EChOFe4VJZfQbbDW64z/KpwpMEB671I+Lt9z8v9zjXXD3t
rTVgciRtmBhDeWUZSZ5hBZfIg8an7mdz5VP+P6XqrC4MLYiKhZe/RTlUvI8Wq6ZQ792IA6nQbZgR
+4vBjvq9srj+6W6qk1LwxBb6FI7sp956zc5wGefrhg3iLx9pWs/DBQZb7Ix6upeBBQ/M+0zWHv4S
YXnkztt9lQ1dhynx/n9FvHJAHz2aN6dx2OMy8u/XY2NbdViG8nbu0js7XeZ/iwkzTRjpLRhwMyl+
RGqBK8w8NWVxLnnxTqHgubOv2pWI5wRbk/7r7RBjij9pAa+AtXqZugmYu57jX8UBaAUZthaUYOvx
jCYuzco93okhK3y5oNYR7i6N0M19+YQvPIFS2tZw93KGuTPxIl+QDKBLkbQ/2H+io1kc12IpKAI0
V/z5DGSTeb5jzz14ScAEuWXh45uUpqBDYG1/0OwTUWZWNc9oEIrJ49nTkd85tpyxlK4FmyFPhDyZ
RXBb1z5kTEBYitpKN71W6VcuzE5KcruZBGI277H5wZtXRjgjoe6Q1lHJ+ryYOzZzBoUev5j71wGQ
SOS3Gh3IcFJcqJeueDAvjQzF0o7Au1TiDKUh90t2gxbcpb6PS3XbS9KIVtVQBO+qLDmHM5tBBODm
CfqG6STZwTubXSA5vq6sQDNhvXo2chz22kJAWdac6IuyuBNuFrx0Mv7p8t8Z+CFz+t2Yf2h+Q7Eu
wb8ciURrHib3WSDaVdtXaLkgHkmt3ysDHV8nTAOY1a7gI6E22M10ZB3cqsyakfFCX9zO9ERaYwvm
gPgO/ifvDY5C0O1tV4Id90obElxDQstfVvQT3VlhGag5JQbEacR616u7ts7rNQDtKmdMWM60kCKM
aM4t2rghmd6E5WjS9Ehl0bUpNza1lFgiY9XTfQ3TtOS75sJV8g4YcT7cKpQw9Kj8SmeV1DkvtPss
Co8mxwvucwlJhYGN1LWhE3KDIzkdzi2RX2YlTm5L/RxLRCo8RKqmPWb5ErZCK66ukUqMKOrl3Xov
sClkFyy7wRc1KEoMpyjCai7cIZuQnDUxHT/J2vF1Gq9If0u0JKMMmEqKLSVu3QNps0jWI4BdDTJx
vXDuGQ4aXN7LSxYW2VBfm2iB2tYQ3Egq6gBfciWJizRcvbTsClA7kQf7aVEJwZGkY3M/M9GEaLbl
EEuJB5fmSBdEWJhqnfw+QOPLnbWwRsxVqeFn1Mica829rOe3Fm28F6c9PxFwQpC+T9z/m7NcL4CO
yhqoAtOQNR3ws0LeQMouW8hDmbLdTCZsHJRBuLJVqPXsNDDSln/RHH/9X5gwNpSJXVnOeJjU2O1h
bHwfIe3V11/iwEy6F6ogeKT+EwkJz3xABmzm1ZnA5GfRS+Q/Nl4iNxzrnBWyXNIcn4fK/8njJ9dZ
ItE67HqKZWnQ241uFiEtdabJrZE4lbrk13OBmAgOdgfBCeI59Cy8QunJ321Rtm23Ed74qcOoVjf4
XSHUOFWxhDzgZwoyhcgRN9wHGnEGOPs08Rq9K/CoXjdO3kpYfHagA9AjChK0TT/ZsUlOmoRHl+ky
wLA2fJzQyNwv0zeN575MixUEmR0yFIn3X2zSsVr8G9EpqhcX5YSIpbMMURbjvhGZK8AMN6aS4HrK
bpbqkrsf4PvlfRFjKqISTb8n1Nwh9JXTkIjBfN5IhgnvbIbU/n1ZGk7waAczkp/LmQnvOFVZLIMo
rzXezhgdABswgZdTqR7QamFCuuZGTSJbKc5FZoeczdtNfm/NeZqyUFxL8vD653uhfLoxLwpQgDSu
eq4pKAFmorcW2YDARmXpLaOFcuQNmt650dAfSc1/eMM0fLHcevNZzbvCyo5pV4oOrPMXmpkM9lrW
c8INKZz0RPIWmHAzo4LAuq7nBMZX0BWPkXMC5lwwJPtwJmJU61pZa3xcEbhuYJbs/FsCVRVscQce
Zm0rNj1eJ/nlGs0CDGP4/ZRYg2NCX9niSxUdvpgK8uCqkzKI7CjyXix+mgHfXxMhnq/Q1uBfxEgc
d/edu1ULu8GB7tz+Vm7snfzhYzI1717McCl95m+/YM/GER+DTckRPIWjoK2/gXS+nLoiPpaKcgb/
VlAKP5hqM/IScBWTRQNknx1srqs3dBD5NvpvUjyT4lRNpp4uKjscdaCWfNgpzfR5Qhy83xM75UK7
805SoF9JLPDAbLtWGvN7/9hrjXwpkSbCqcmXgT6mPpvzoEqKMkHx3NTYA8/EGqmTVpSCHS5rTcdV
uPT5KXmu1oLO/KXL8FfEgpb96mfXk5/j5GjIpUb5ZOmxuVVXPhONfud6bhPEaGYXKaz1HbkOiFp5
bVfoY5BpwsyhvY30iU7cyz3b5YG6HOVrRqJhMpHq+ITbzohQiz0MF1QaTSFMQ22lVwGUVtoBGk4O
tVy3oMuVN0XDiKzyP/AML8otrsvt+CpRZRKosDK74vHe5s/vpluF2nNoMnK8+m0hC8iTcsnqaxLm
Nl73m7mr3Y2nAO0aoCJSer1f8tUYhCJqcRKH1r1KBmqNB4CKEDP8pxiQorWv9TFaQMmIOna4cqJh
zRTT8+PKnLPMK/lC6Lc+ygUOtKJpiM8uqke2wbSljHfeVhO7qtYo6KkOIEhsd/mdKKs/pIGzAxgp
sjlmyWCuTeQS7veN8xT6PQEN+M40RRfku24jTS+isW63vsPZwcstTZIdVbhZt1PN5lrKaQ4C9LEq
3la+KKrVE9gXepxJ6fubHVzXDqsGZXvlKxJ3dv2lzEANU4BDm+aON81AEh5QIEy0ogTSeEhJH6Oe
4f0Lav1qO4e1QV5rcHPaHEQOrmL5VahlbsmoBHyGsf/lhSYcEtCaHxUuufeAnpEueImsWIyiSrwe
A5Uo3qcYPEMG6KGFl2iahpoEh+ltWIywyjIS0rlXgoHKZFzgkdcP+OPrisNPK1Z9aLCCP8wZstsD
fOcZ3xgSMcj9PcuzqWMN+3sb5T9Cpof2yIsmjCPYznlUozAEAiVpZNC147Wkwgf76sG5yNgEic+7
FDqbSVxZqH/0TfmmbeHOwA6wCg47UhGgXCEU2BqYxP4iVui+VA3O0/euGuKO3BpweKYYhBalu7gw
fIcmlYDrFv6rYrOdoxDhhklc/DV+zo7eFty9bR09TEBzptPFleLj3rg/ragQXcreHcgI4deWeo+H
M5O9ApJCsnO3zOHQRGZZ2NUKvsV/rC84OI31yP4g8dc+ZQYGsWsBscmgtv06EdsGMWZ1N6nZUk9j
4tZJdcgkXKKqU9Xtdl7Z2AazY1MFad480RCZ1zqWIg6/94C3y7QbkVuXNrfK1EbMH6c6OIobJx7I
B0dMNiv8dkf7Oq9B6C65UMbpNUZGBW6d62qMnG138msJ2mEGMDIYaKQebjJmNSPmCBCigCw5psJE
dzDAwV1m2ogPlorwhorJ+OlwbJVESRm8HtPgRdjn/KBMa+2RFRmTcnbBg28FQ7ciLJZWRukWGM1G
T/6BlL/dOTcIN8mT09R/cyVdpkX2m8kpvOVwfW2EqTiDe5IxnjU9Frhct0PPXbHI/ZtnCGrESNra
1gmeBTQMYHbcvXlibyd+KXHAj6uuI0wxUm48c0H1heuvXOYnvhxUwATR1MTmVAT3GtrTIqIVZcYj
qlJ3+b1Vtxrzk4MTDEZ/7vmXWJ1xcb6vpsLDdQ/Gdo7ESxZ/PODFGpGwYnNshqBod68cL9d4youc
62A8q/65Kx1Cfn4VxKT2n2fbYVfA7bN0ngl6CuXPr0G2oJl9w743kYxRdlt2z+HyXysyvp0cu3lJ
Aglwn3yCJ66QCMi/mNG6w8ejzp4qPza6HcqddJEC/WqOCiKiY8nKokDZci67FUdfl5yAwrwoD9LH
L3aXNziFXr9dcrGYbIx3B177JUHuLp1FK9Lqrr0Cr6ovSM1jdZWc7WUvmYiNsbediNbVh6xRY/HT
WmjZ8QjVjhoOaf40diyLY6pJ0TgeitECxvSiVWpBXBNJIptwJPYer9XgCHWfWuv2G4uLN4Bnpd4Y
roHz5njLIt+c/hP3y2vCXo8wkBl8P1stqTSpuAFfBywZaC686r4F1hiD7//0KzszILSzlZqy8rrG
gAtdb7MzX0EqnpRg8tfkO+knDFdLN+NxxJ+hN41O//vsDgdRXYFKVzbI4SjCxsbZBuW6698xq1U7
NYyie70tyhh2u0AziL7vMo46oRUEGgzs1QV5XsMOELV/rDTm3DMFFD+53bzigeYGA4nU9BcR6ja5
4br9CFah/8QbcrFoVbYt33/JxppB0hIwRND/K5E79k4OQGhfr78Mnd+CRpPPDBwPoQzSOmkFXyNM
irbNZkykmpS6JozqnV3WaFs6DhKhx8lGTPLeDvFCbz9mpmeIOTZ//osVitYqvBUchiG7X4lSUs4s
Hsrk4mw85p9GVNAwoXPfDSO3wocnimHq+kF/TEheEyaZEnQ1ldYfbIo9c3zUbcUZBvwaXDyBopom
tSYAaUsjWx2BgPkM2qznejlGZkisCXW3JU2dS1fyJ179gzMaQvZVk4VRfcf5Aki/A7nTN/V50Sxd
HFp7BZK1I/EemGv4zrOdpMGkneZe6wx2Dx0Z/swiaLO7GMpcDPv+u+GNVs8ycffqT2PlQK+Ruukw
974lrSNI9uykFmGzia5DBh3Qcgk98Za3MqqRNjEXuhEfYBvSAtdZfzMLEXTkDeIjGrFf6Xq5Zkn4
QQvDDNTdwWlhedgLw0yRr2PA79lWc4WKsbWjPIPwqcpr1Sn+4ciBtg4KdpSvQFlXTfQ5qYg6hOlh
vRea0qaZSByypRurv42NjqLydPFzQ3B2ShT1GxNTw6TJopEguidBqkolJIJFtfYRM4E4L8kdOxDG
Hn8UwiT1p3thGg8jkLqJE/jNMPFfe2sBzV59wq0VmTBJgWopZCiECzkf5/GLjiSspwT3+P0Uq/lp
GgrSF8Yx7uiy6zxbZ/8j4JA795vXlgvMOR2rynEP6BdHTGPQDpUovgCrfiJ9mRjgC/GugarOscry
m6tkQneibS95pUmpXgE1lvDtlKgkrNxgi0iTv0BCZqsLTM0yAW7IzvFMTSmsFNiQhiCAzb/esMWW
5qmGP5HPRhHiguY2Js/Npn2XlvvrNn3smhsdMlDwTJGceeoEyOD009o3bQDDNxpWoxRgXKPmm5in
X561KbSiU38zhLb+9Uo8sw2SYJYUepkUdZgXPMUhdNnTe5EcMMnfr83RWYeDDyVgDtU8778ZMtO+
hlXAq23A5z/uG1IzXmvHSAg+llV/mAI/xKImxPURsFbmocwctGjwRX5IT3LvSkKOMj6aGukZW9m+
L25AOAVqzDrlPhSUY36+GM5qs+EiH3+4DNZ1kmD7ue5KjFBXmQ8mSAbllQ2Xxuo7y5ZojpVtYo8y
nTZfyDCSoX7R515DwTNt0dbXrQNKEaPHTgabwC2XrZwnWci3RkmiTgxgDicrCGrcNd+AnhN2IPWq
CZzhStuGoYGRDsdNqcNRc3HBtokJcFZZw2Woqb4hhli/HQ+YW4ndKTAWRWNByTNIUzqDmClot+7v
k0soLpwXTcJY2zhdjjlopYxjtByqfmDBXw7jtaHPOERKC7pGnLKiQ/J3hjZL5Hnu6dS9HqS7GCzE
vt5jGH0STnVqqDoD+6rLNw/aQWmCj3VAoUevCoLLqByKdXV6tq5eX06s+ivognlYD9i3qbYdT1Hm
aear1cSPUsA287y2AZORhuq0rlm/sYe1+zK2Y9YkHzVKzTBUlVqHk2Imsqx3VtzvZpEn3HOIUG0l
oGVOQN8lBTTzm/6BdSeoBOINyB9GGnitPs5aCR1QJ2p7g/FHYlBcpl7Fxt72vDDDmprjqpeNsUAx
/V6vnoqeYK+atS3ePWe8KqSpBkamxem0xzO8U0YrwtFzZZalBfWjmZNLPPAasQPOe/y6vElvx+Lw
h+uYFT4rGSdAHzI1rnTi2qqbPk8Isfx8ezGpYTsmzlBsyQHGzR2xB7gZtZn2Zhrsj1AwhJqkNzbQ
gzh/d5O/6vF8VPWIl0+Jc5ANu9rZBypKFtNa+ul+3vD9d3+q4MR+qyrMNTCHeVlC115g7pGfcAVf
I+pWp9sRQvpXImkeRdAupoths9TANRtN2eR7T4jxggWg3v0NO11czGVEep83B1HtTdAn0rfJZP7J
hsH7rU9rrWFOJiaeQozXZkcNIBMCuKgFq81RrMzf7OQKU6d/EpjXs09aJb2H8TkQuZb6lDh/+aiV
Tjr2iJvoMWy4XFLejyLCWTU+1R02dGDkYZSkuNLJgOejCFgIYXMh6NoglMnSorWsAOn1f9RLp7z1
Vg7siMwZgVZIdqvA2ob6XTOXlacaOmpgMU+KDoOm3FKLxONqx+A+fjeq1EnvCwaId9V+k++NhYq1
SQu4803L+u4KzUXiGHDqcARjGxQC8NKdsLozLlcTW/edfDaQMmULl4FrjZPkcVhAdJ/Mnib1OBQG
ZO4oP7wput52hfxiNtEKv4fejwSSxpYi7pUaLFh/5WmDNMmLRcfXY44Mi9YsQaiZk658811S1YZW
hSCw7OZlDwwfGqfb4xHsuDJfohDu7ds6KwxtcHxMVpAxZqcjN0TXeJ24+XfY8VwgAZyZu7f+S7Qw
8sC2IztYFpGncYezbqFr4cSCwIYSEN3jEsgSXHCTbFVmVcfhk+I3WjO5FMbp8QwHEWlFRv2ycIK5
fo13r8d8iKL/Kn4cEfd3PR8qSVZCwZbuaDOd6fDVwJhDuBqB2hOD/2WrD29fozuMkpSdRAkT9+DX
JpdOQj0+cUMVHgBSgqF8UJ9odO54Q45wmXr5OKblcrX7qkg1/YgOOtEy5vKRHqqn+iaKsC/DG91u
qF1rgNXRTLtt9K8amECQI4FEzmoMU+AxRpHSs+lJ1VxF8U9Hn2TrhPmxlo8zs1fOFrRGmdE7rFiC
MPfXKJWdFAQ/WpMGoEYyoiHFgykwY3wA+DXqckqQTnxjipNG2ATLMupL+z3ocHaf4n/elaRy/5KE
aaEWlzeESJID4XVEUfkLKU7uX/g+K2k8+PpLoFXQvcfg4lUdUpaPU29sJa73dk13FORUXAxem8ec
ctcJMF4rlzyz41LpcNvlrR8+0Gw6fwyPsWx9pnltHsJct657a65lgw2CLOQgJSfHHPW6IrbUmAsk
u5BUQ4FHNjU21aRfXn9hCIjCrGCpsBzZaPSUuWLDjrzl2WLo/uL1gcqe8ei6ZUbO2x+LSnOWWDpA
l6OpSLe0WemkR846NPHVYPAQ1SI5YQfiChZtvE3WZtw9hb5R9jQJv55TcNWSk3bNvKu9BYQ/Ap+W
ZT3xghAbAYk3/OeR9Laj22xnUBvcQRCr7+mluJblZoxk2WQTnRNETdnVnVdR1lLbfJZjy6qxySvv
Ejdt6qA2HTbUtn40nYCX3LQiyTR5euz96L7UgaqPNb/lirrud3NBbhsmH5gMIy0h3l7n0VQUGTwz
HZgtkoq9BhqtNqn1TtstWrziJNy41BbIfO3FJveHY3jyklyv0W0z4RAmInOWO2uvfGv4YdBNUQ31
j+7MyMAchsppat7cpcZOyOFHlLvG1s1KOTUkN+oaYm1sOyBEgxUtoByTYb9VnXwsnfXCR9srzkzS
EcF4ndSXR6jI35ZPcBKEuu3ER+4j4egz4A9ho39g8QFrEqsgB1ca5z1RsafEW11vm5e3LCr6T5IH
CRxibrufgXxyRr4J78eWYwoeq3QsZBoAMxj3K6CWYG6AYLlTvX5/gOWlJJujxPoFc9DZsd2tOrWw
S8o3BqPaf4eiHJNi6rv7JtzWlLY7VTdCtOmhMPDG24FvvS/gqboGO4xxhCFJzl1cFDcejraZb7qm
EeRut5clj/1QiVLvlThmzE4gVtd3SKhy5cUMP1oUX06qcgzITKpmbO+x71cjffHRR9YuUXkq8kTd
VMnvo5gcTBtlKw/6dPl0uhPvABrXb1kWgkD7Iez72mFA7mSrRSu+PS87Vme/dYO1gd+Up1+9mmtY
UYMkYLzqsXbsmiCF/hHon4VgmqWiTRSDY4uwUrDFBDnNnXZmiUNQH678Ejp53wWDL5lT2ostOBD0
JtonBEXMegtSLvi26OpwYIgCbi91J8uTZyxMYGUNZ1jlUeHigLcLZsrYqNWbVuxcO39JfEuCEQNK
8oPyYNsO6Gd2PupEM969ZXgXC6LYotv1AcOw2ljmVg7VD0v4Ug/wa7MVEIvJX6wkrzVbHBO4bLj+
WvUbrkOV+d6moRJMQ3AYkThSMYmUDggDSR4feJNI65lv6F1HM1G/EDYGMsIa9NcuWQOn1MBBMawI
JmqB1sZWVXDZhd2ZozBZ16dOD7oEos7y9cjR+/mzh4s/BXJmWlnJMWTogOHSbcgqke5YXs/QgB8n
CGF9WFt9osCvRVEumeSmcvR3ykpeql+oN43nX9i2bcgvF22+pLnmMMyMWOz/1GF2qnq0drqEhFiD
6RV6ddwOtkC9WParBHCzVzA2nH/GXTL+vEbJP8ORYp6z2E1m0rNfBe/zlZec11VmSZogD0e+Aiva
rHVmEnIKGoXgWdvF64t+KQA4/NwUbCynWE6SpVHq1q2SED1UEqsEWl6a6fe3TBI2MPf5ws0QWaJu
nepCCPS13+wIqyP/SZ3LEgj5FV+3tdjcT9Mi1SlhEoL5xiP3aAbmHd2X4PPlEMS5knBAs3TmrPyV
0Dux30Ouod3HkEWNFDhgWZmdM3UrrsxSqI7Pf8P+MN0gM7qOewiDzNOom6YKno90hGEaHktHcjCF
vfJo8nHNl5l4hdihyybWIFuPaRNY0HhP441NGEdulRmL4zVAxgX07I0x2kPZvNkV0PxnjFCfvFC2
cWgdvQJeqWXzatd3q8KG1pfnM6tZJzNp9ueDQPJDc08o/8fWjPa1T6a9IxukGT7jintfsrnp4Hqg
BEJqiLZ2dWHqOqL2CqdgVgXSqbvSB4edGOaQSlX19Ezfphip5tlxIYX/6IFlHO4jTgaTziJNGz5c
S7/C09HsS4nqSTzKY/GXfLIkMjL60H3K6P4pW7kVbolu2dtoRXTuaNrzSNpk0Y5mygWvQJitfBqV
i5T4Y/PR3DyWujpAziwKp30+6Ah7eRjrUWOySqpO+5FzxoOCWOsFEqz0M0t38rCIl36mAwjEwqFE
oTj/lGeNZQmxpzwMfzG2OiYLRbiCSpJSCCgh+qY20zG3Yt5ey5zhvQuvB3T5AhWO/yWAOnEMaqTr
Adeyvhiqfx6bCFTmaZeogx2E4P1g6bjP8s5luT6en0AKLwz5XDH6YzaYYkrgfRXotz9/rd3FX5sD
glTjvUWQCkG1MCvKMLEkF5s7f0CpgKi3IMlTfXFDqzpMS3AvAuzNYhm3pccWjQQHv74VA7NWbZ3n
YEijCsBWLG86YBqaC33P7uhJoARDc2FrGbhHbcbtJOgeumLWdmuRDM7llJbs8gU0fyk5TrkYK+Sh
E0glDM6rVx00JTu9n9kvIx2T2W03gm5TSC+KBArDrDkpanqLBafryC911F1O5bRs57hLvtuTIO+4
sVRx8mOInFrePY6uJVfoQnsWoQ4G+/Cv0CWlzCCWGytNka4fuM+cJBYzDSQfkKhWuvuME6Z9j7rf
m+Ll+4WirmWCNINPdFKCcj++sF2yKQxEREYKQn4PFGqq2JNrJmw6YD9IynZ6g6Lpo6xYzUfATr1M
e8MW5o9HScqhAIxjJiuWI/HqSlNt/L96hRW0vgamwOvR8tcsrhg66avBhoF3kVqTmpG8Za6jhNB0
TtKwcKtfYk+bUoGTI/XQTIH+YfkR5BXjxYJC1r3+ob5yaG27Bz6UeONTCJcfKwEXTlBDfcll87ac
jy/8ScizWTKag4+aGlqMPRki/Mik4+7DyWcqF8YIr5Qt9Clly/rNy5U3yP3fVQknKL+y1YNMpm7x
e7lgoObVLmTum5Z1bW04zeL/pdBPjopsyPpelcGC/sZPvPwNFYdQzihOEOytCr6sqXb24zfMtu+x
cwxY3Mx/ryDzxtlnUI1ZrlQ7ULKBoX7OPsFTpbAC3E3k6aDaU6S0ESzp+jSESMJAwUweteWuFTq0
OxDer1xFgzwf85dmmPKkiBnKrv7tdjHDdzII71F95d4II/Ye2yc7Yc1FBMw4VfRr4eJvv1k19uYQ
z7CJMIGId+R5I0qypLEf09YdbanICUfdp8Qv7VT7VpM1zXn0LIK5mppK4udIa23yWbXW7NF3BD2O
IekSYcEyJDp68HpHvUnfb1WXp7hBu3h3vFPmHAERveUdsFKDAYBwZ81GWyagJrRDI6uY2zPQVBCR
Wi/4nkwZPWbjpYbv4HaQK/HqTdJuMegPn4gyrocBHvXI+kb+Ki9gocUt1cCzVFaguEeIeNN0WgKU
0Lbxx5V1VA4Hy5ORl8jmC3Rf85Oj0SxmGRVDW42ds1HBJJwacLHsRv/8iKFHDer9gQTAZeDn5HU2
Q7iTxElaHUukHDAY1JAXeBig27A9hQ9RbquQpHRA2ZATj6uSN/wqmdn0+zEBj/SAVzHN0YPfmQPi
11Kim0N5+uMkdst0pbXgJ5z7Gz0QskeqrSdEkfoTIlJe1qMa1qd0v2/pPPD2R2fhlOGTnwKbW2ea
0TRPpyYuz7BTBPPqIf1d4WQeyO9W58BrkIfR2tEP581WYbHyWTxlZd3D9gzKjUbKY35PiYkLmdDE
Bwb6Y6d3af1wghH7mx+TbLw3w9IchRv6kItAlJE45CZxVFzDUmKkBW1N83ODDdi4E9jCX8pu8wGT
bSPSIKbDlhirUxCRWTDnhT1UXluvM2tiOKKZtJDb2zKwXXQhcTKEt3wbdH3OZ0l6cQSibFPiVM1l
0CWz6Lbd2IDxi184aXFBMFcDazcID8Edicw6NxCdjzQ8AuK6ltFtrjTiCX88rzViOn9hR/7n9n9K
YOBnAmfxg5owjOlqfTS1sLVDcct6i5wpHEvr7L038i4LMB1rsVgp+dwEIm743lFi7Q2GwqHreWIF
goUquzzeuA90DQsRExOXxlSUGy79C416keKgNQUehkN4EqKuTNQ8b3q6SRZNslHKPBnhDtGX3QGJ
q/ET7nc9NGxMB2R4m/OTm1ZUHGFfJusnlYdTWjfzDRRETogeN5o+G0m2VCRf/Mx9CBcd7Rf169Bz
UBNOF7UhUaakom0lkSdUJlmaYMo3NUim97rpdAfwNMuHoPfDXz6yGc7mYVdoW8yjJsJzlA4PCVrD
5EzJLynk5vcxYqqDO497HHH+Gqm3uwFXpPhlNRfBBFiRl+nt2R8WmVuXUfJG20Ej6BOs3U+OLonz
7YofuVIapR0pCsh6ycgwdyhIVGG2+/z2/b0EU8Kqkw2s1+mhCsdnmB57qV0xQJruFSJLJERTIAsu
IHAM6TKc/whGpIqDS4CEyDUGb4rtWqxXUlEmBkKSt/yWCxJhSzQNwrCMuwh1sua4yROIJoe40lXt
nW/HdoXpnPIz/c9zteVCJ1J+ZFe6yVHeJtQZcohr0DVlvypb9nbKQqZ8p0M/e/C4aesPIw/P3by1
fDooXRlOVJ7NMjfGbysPjicIEOIbhjXv2XsRKqPPah8Xbkw6EHKY0Yf53SVrnrKSbDnx8TYKS7LL
vjzXau+MZK9P73j6rSLj0GjvDzIe+57EJgDSxfovM5YE9uEZNrfIVs9VoZ+2LpGF7sgYhxSZT5Xj
0T46lI60uWL5Qct1NfqpmJ7IglH/zZ3tFvBzfLymr7qT7Xz5mLjfVV2m2Zkm/LZAU+X02RO3Bfaw
7ZQfdDKx4u3+3zUB4v+yElWYIrv0YoOuXByD5rrUOOXLWbtInaFrdko5mnr+wsdEuzFpUL2KtuDF
Kxj8hdeqjsWueHrzxlXmnlp4WbXJDRLg2vWSYdK5vKsx8iKpkBOXjxHajtn8xpUhDOEPnUyeKme9
IoXOg8yFlVEjMh7i0cfqVtoL5UBvr5V770FC3dpu+vOGsTvhzDAq6Cc3UFRS7cjL3Nk/PA4w59hs
dsPgWLMsFk1htCqatGbH0CLABvlI/EdlPvBF7pSUtMjW+wiFBkY0QJyQJ4QxwqZMPJUTE1GO3KfU
ikwxzG8a0W3BqIWSY6ulVvT91sQ+j8sKXccD7ysIusLBi72uShD3Jj4IBb0qzWs36sclUoT3bj4e
qxdTDhtl+WJeIerjZvzi7ymju6up3jUV0J5/UH7wtnB/bD5FlcqQZsZDbpcrfpXd5X2mytF7u81N
mNc8i9Z2OvbHommChVp6hXmcSYyW7sDyUbLGOgWzppSXjkbtGN0hlbBJWLYGNVVAmdv2wL+Ubqzn
mP8DJJhtAdJTGzQcw0Q3OHmyvv2wu4JhAwqRgdehfo4lzdlVc1eRU+O0NiwkiWYTg0PZwYg2ETH+
YxpYNo8D11CxzwXK36i0Zpq0nlThmFCOZ2y7vL+2y7OJ4XJ1jNUssyxSQ/DwzwKQnkRRwNo2cCKa
EUGstOESXQ9YpFKR87U3i+3XasSh4wBJU79GnSRk8NZ/dcLToDmT1kvcOTm81EQMEbWcssi27ptw
WrWnN6/ZmjqJoklL3PX1iVtBTyZFyYeM8ql9AS+CAs1CETzscwlamSdpwL2YhrTWrl2ZSP6P0ODP
wMwKZ5AZIPUgwVOG8Sj3MVfpc/VhdXK93a/Hsc7yurGcadVi2qh5dvCAnw6fSLWniNPnvCh92fn+
0kKSv5TlYAwvTwPl2jiPladW4+1MEqY1iMmeW9tS5LFs9mxZR0jC7UuAt09q2BxMmGvhNHvZW1zT
QjF3mq3UDP2Gy/DiStWGdZHIbxzs/n4JsP9ySmbyicls6DJaTSlot9BQKPXur8v35PSuAAh56HoX
4Rf4zCg6LMNeUGxHIO7/xhC5v4vLGWTfRm+DmfgYHao8tQVq/YtT2YsOTt0+B52m/xl2XTwC6sOY
TUn5HT3hW6FY5M8DWevdITOsEso7MNwDZ9WVr0P0/VwZrltbhUqpoOdj4q3cNAXXYC0lM2fl+8Nl
5kTWBqjR/zXFttqCy6z5JvhjX5FUFUl4OunXLrnFDXWYL9WKU+ZQR/MnIymWxIPwz5GtRrpys7ZT
30PyCF9rNREnf/NkMJTiZzDcRw0VInwq1DjCTTJaaKWhRSzKg3jHTWubQ7Snp1vyI68JFMCSHs6o
0M9ZY1ABrU/pp+a60CJnS+oy6MoT/yv2ntRg33FQILhMSt/jprH9reeeE3/CD0chg+IXoiyof2wE
OFNJW7CuMt8Mku6xTYf8rJI32qLPYZLn3j7uglPwZPYkBeBmHoVXS9l/j2fD0eFkLjIczD2CNAlt
ggrBFy9dH6yH15D3Zy7Sfr9L1UBOgLmvZvz7pl3uK8w2THB7ZYws0UidUEjfW7sWOVLQtVuToUdi
Wo4KzMZIobuIWgAfpwLRc0zhuINp7yK95PJjw5gjPiZB52fnE+yAmg6DqyYSYX1pWiw1W5VgLOd/
Dgi+mXtv9T7kbNHCwa6c32XaAK1HRsa1BtvjodMeE18ao9TSLyzdWSrCqjMxtSSS/76hAhnQ/ulU
OmS8PRsD6CYRy3DUYmZ9tRHT5yt4vE7DShtzqPSQ34kxr10Xb0esuFQiU1ArCOWtXnyTE/+GP7NK
3ETh51CXgv53kn4k2Wr4Xgx95nppxWgPhHw2UQFWNKJNw5FWatXbOD9rQwX8hWcKUpA2pGfmXTY/
GpkR8u0q+NxbfA0VghMy3nQmX3NmCyCi+DJsz7NKVWhmKuXppUf4AGOfzbQRWGn0bndANJ/CDQ19
EEXmdYIvJ5VCq/VFvPaw2O5VliAZ04nS+VxTqI3SYX7kpES083b0AHgXXL3ZT0uoqs/zCQQ26ceD
YKy6le6fUXS7mZ1wrljc3Wl4oR5gYomJL9ktv9AnW4dpLjiSf3UtlzfTejVu1q1I2JuQ0t7rVlpB
STLjn6bnya5pXauj35uYxeqvhdcFnoe6xSgk+vsLV88zfiaUOJq9uT/9R6lmkeB3WVWH4zjXuEs2
pwCWR3ggMZiscelrkOnJbZeGHZ/V8KspqK4ZtvzQgk9r/b4QSNXU1Y6+N4/CiihEF0tbWppJ0jXX
aOgs0MVXewRHwGldzu4FPSqmmF5z331Lt64Fv/es/h/y4VIGf4o4g0DT105hJK0wmlo7pENaTnx7
VGxWzm9LGNfsP5/QgUndcLUnejI4j5MGqthI4nr0lb1vVd20NvDPRcuyMYcuzi02SUrIve1kqolg
LfLimi1oxOWifB/TGwrtDnlAi0oHuIJ7q3DHUdUWir7kz1RYYg86WTBI10eIgIQ6IweSvERVICnJ
VCkfM2EgXhxvHz47k0K6LxccfMZupnGI8VzFF5AVrap6Di+Kx6z/TIxPFegLRzTixRTTuBUVGIzc
YHN9nuDjekEbNrLnVefdjFHHNU50cOWOaOQ1Lb5b1742Y+S+lvF7Y8KnVnEvtfK/fJzcrF/tk63C
VTVk5/Llyn9LAg3jHsCi/EML1t/8M7y4oT1ElouJDVE+mSAWnx+9VJQ8jOeniCQp7mIpivwwCmx8
4dP20ysW0r806N2aH4SNwjMDx19+zAC6gksHAFFAm+/nUhuVEkAytX+1c2NhXkidwDu+7YJIPMMA
Q8BaAHmweXxcUbaLH7dooyCCZiH4qLUnjd0DVefeV4c0UzMap7LtNO58sBoUpgujIlvaPO0Smh5m
67TiaMiHlqTdepdoGvewhosbflGFdD0GgJNLZntUAHIK8bYLGFygaDfeiA02oYxMd2cM0kClCJbC
/tnWNLFmtvzaYwBkBNwKZHAgFkHMCz8owBEltKrLsbwJ+ZFMd751w7blgtFwxH4j8ickPrX+LXTF
eZk0g4hz5hVcUhSRoF0tOnOcPrrER6T/StGI4X+rhhBS09tYpkk6tC7su4q3j2pbAMeyg0ijMFSG
ELVE8BdjJFgKaPvpJqPRSk9yKCQJ6BocK6Ek+6nGKqemo4FnFMyJ7fO2IcyOrNy++0+lqs6L95Do
t+cNF/E5fpOfoTO3SL0edweTG1n2MvSD/sNWF4x5U9jDvKxGP3X+sxxkEFQPqWryHuJB2ZEUMYfB
oGUo0GajNJgbf/7AMICjy91+fEkChz1a4O/U/xLbrKBt8AhHEHwfQSrt9eC1c5n4DjjbIrxGIMaG
dU/xCk2vwQoN8KqNXTLR6+4Agbr4TIQzQ6V0MsQmArp5VdSOcjTHr4GqLTswQouL78LKlVxcmEzg
roxZU+sawbdzVLIRKbnbNLtA3eIoUPy6rT/K+41CqnkWGytZxUHLlwQhJ/3o9VzqLFEbF+ETPIfS
aRr5oXgdA1CWJSKWZKp6t93c3HrIeVtY0+jiJV4e3SiZiKx+jmTsmNMIAdewjobOAiDyonNUnGBT
K5C6SvrCtb372nBwe3pswVmTrfvQd7HV5Qgi3Gh8vyxaKjRd5fTMD+39U+HgYkBpfVnPiDm7zW5u
Kh8sdEvSb45Zut1d7jI+WQ5yhwVINcnRsmrfb0ftk2aXJLI/cW2NDWT21ZOoPrdHkZ+xUfgE1hrC
F9V1bQpC5zfKIas9xeILIl2TtxUV6rZEfwxlEO8Ldx4+uBCLmrvx1yPUFuKOj9PQGjY0rkpkaphP
UzkbKrrRkABMsWBZJRzpU8dwjLEZKm1EMqw1AqAL0ov8ncVApg3mwruMfzu0L0vInP64dSPGfq9L
M1V9R7Sf7tLIMc2deaV25kXJGOwHz7mz4lO5p7WL7ZHl3ucMqYepOgg/jjN70e0LEhsu4rYblfZA
3iC3vGdwtgRguWpVxHiQ4glYzZyl/l0equK/Dw3sSI9IoOJ9Uxe1rtHLxPMRXpEq4t0Fsp+PGKvT
kDv6tVdoxSDhHlxwL47kj0O1BJAbFUsKE85rnP+YhbNEImeQwFqfZR5rBeuGtJ/XzI/rJjhiWrqx
u8q2CuflzxF1eF+51YzMRcGrTeEuduYCxq175pLYGXnb7L17GaQfya9lC8IdHmSzDydjQRVy9x0k
yWF2dala8qS217ilOkIHOgMdAcG/VLjgnE1A3G5nyZ+uaOpSIbUsbEDvWHx6kMfW8aylf0uBt76V
sCwjMol5KAl/XM5llwKAK3YJRNplKwny9QMnerMZ0Nmx7Arce5ZzUFP9x+ba50dz2Z8dmgcZYt4e
5HUHSoFUrGe18e+frcR7+oXAqJc0is13l/Jf5fVUnKVvw3dr/u/uRMsO17dmu0AOfROsYaQiGCsi
3bxqM+kZ/MOuPrKSUTxHTFhapIrDFgPgz8zANNh+m0PQ+5eOmpOjWb+CvLIPNNS9D7WblwFEjzYH
O2Yh7TbCRFhcv1RIKOm+a6UJ3SuSWeqitmzw+o1e6WYKA4s1pLpKTjzIf3a9iZOwk4Lvu4hyg6jj
1z59p1RTg/tcm6BEY5le7Z7tZDYHz1kOnhxPt63k/g1t8zo9/hN/6xFcpbyVbDZunvPiDzRnRXHO
n2scbRfc2yycaspPbFhVGRaYE7tBH/5h0xMOuK9LJ6YKGRy+I7B3gD3y8mgKASYTZzi4+2DXgBgI
a1MWlV66f+cibGuzo6ltOsLVnnNQcdNPYVgYmrf5BqZUuKTutN699p4WXnXcimqmBIs97fXSZpLr
jwbaFZGW8SDhs1EyEJbW4evJyE3WfjqWnMOWk5QOp7dploOih9wV8+vQurveNaPYSbo2SYXrdL9O
qVuvHkQ/r9LRvfyHL0qjExNrII7M9SrSA5B8OZCdCeWJpASavNK390NMGIvMhsnOFu+85W22VRjB
LDxNturPrZzZ/UdC9i22Pm0MJheFnQwn2k00XqBZpOU1s6dhY5vWsBmyQla/qX5aCPf5iaoPPL8a
so+kWSGunIsfR+UtMmHMtA9BGjzHczczJzLEseYAkKT65ihIVdq5Ej5MaYz9Yc34lB1ZOKY6tWlW
BRUeaOFRoMoBmu4omVRjCGwQfK9KV9nVV4Fy9okp676ujrHa1GW6vNICSxpglk5aoXOcbppoU03I
gUSEvq8M1FdBD7rGnOlNpPjKMFM5JqDjQVffyqLDib98ZpD5Eok+9dKgqvw4en1J8EvpPItaRYj5
Hsmx2cQCH8//J1MBqmWUPF1wqtb9HcWl0xmJldNg6UMTmUw18Hr2TxWG05Zj5GcDqbB9dp85dwKa
fyia8blbuZRrMcrqYuzAv45Mza4gK6OlupW+yiIC1erd8uYi5Ag7giMNYAGSYNV6flS91duFbOq5
lViJJ+xTHp4prMCcigvNRhWdaP6g8oWU9XySGsaJths7ehCr/2Xu8u3MCydVQtiZoMDrJdWJ02/K
9Q5EWGm79Zy+s41m/GRO7DS5uxdNgU9dzHYWxXH7y0l2CY8qIFspGoLKu3ToiJO2ruJFXxPuOrIz
oy+74TTIDOKTgfc+W4ae3wPVx9ckMNcQyS9dHlrXpOev9KI8HwJAnxPCeXEhNF/Sdxr05rKoeBY2
Jt1608qgUR9tGvRIjZuis0kdjIyqhQN8l+ZkaITTlsdJXOKKBzvUGvRPCNRSF2xgX3DFE+eTAwGe
Aj08T0QugKw9E3OZQHqMxszdqUDh+1eYYZLYnxQ6Bre7rTrBxtWqE+hjFz7LShBOjjqsTVT6H+L8
FrVIN9JMc/Utde98X0G2qtl1cWwYvmk9VVJoKXA5ZWW2bf6TmWm+LR2OiMFMfnAnPm1RZRG4IExQ
rQAYGfy4xzROG+9X7pM7o4ATCGa6pv7i02sgYkGN63bPQQK3+JCgdI+R9H/df8siCWU5dNSzI+j7
s9cJ3dfLjjioG31ZuixicjSGsXgPqEfDvtmrG48eooNkWP/KqBpfKDZefXS+bSA/GRSgsYMUt7lG
USAABdp65DtCrrQXbye8cfE3V4cIITarj4AnzmTSpbibDuXsUNijTmYGdShY5yYaIvwd1VU2y/cf
TpI6xUjhDkUSApsKUAacVHnG2ivK5PXmlABMigNfK3mfLqV60gG7YiDHtApVJjKOTAdHXi8q+bnH
u9WmLvWW3o4YcIHGs54T81a2Z2uzzrcgtbVEnWiN5fWYnJsJBvqidUvSOZRe2kNL4zRvIWJVK7MK
Nyj+B7Fwc6CMYWE+y4XtBws+fKBVLvO8p95SuxgckJUW2Cmw0t910NUJYXPGrq/c+gb5j89uK2sW
pduNs91YcRlSWifJF6akcrUQHTdQZ2vAeRxgT4v+Wge2dfeSKyKr4pDosFdpY3rb7Xj2wvTzbtg2
6+1pOUNbV69yXMWAPS0B792pPZM/CcIFmw31oHsOfFZb/PPYa/WRBrxQeg4K1h0rG8NrgQSaZOzi
scbIJ9F1qLpaQvI/zrIc8+xtf91POJmuSIzamdyocWE396O5VQFamBmqYCvRQQ9gGVsw88wJabDm
Brcs3zqYVTdixDOLcGZ/zYDOOFst1VIl6knMfz23Sdp+tgXsAe/Njli2Si0uWtu7MgF8PHX19PZy
O9V8zAkqpTVZA1a3xW1PXETWPOA2hPwF9MyaD9x8WAe9ZT0DqFb+4KdnYHgwe25XjQOzuuEWO8/F
v7T594EmivoeTwC6ffLIHztF0avjCBcqsPfHrT085kWCiBo8iUr2LljUpGWin26XNAJolmmpewHY
ueROFdrt6bQ+VxqxJ/wl93qWslJffxpA9SzrGg/kYsA=
`pragma protect end_protected
