`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7568)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEH1cHPlahAeeD6n06w4uaJMxNgyqKJHatxFMHzNCptc9re995aHTFELR
EG7g6NbBSopK5XoQnXQR5qIQZuUOSj4Guekq78o4eWo7FeEoSy/8+Ks/PG9QeN2JWnKykf9OAVIW
0LK4BKF7NEyZBwpBil4EJ5ia31Addk51ty/EoERBrfUhcT5JH1TMLmldF1uDzfcBqxdGjDcV3jrj
6kSEM1m9s5V6ybWIxgVFikA5Fvm2BN4JuAY0b/8tNyxy75MMFkiJq1dM5AeQWsLN+u2piq9fKGA2
KITanCiyzHvU3LokKYWqpTp8TjX1ZgB5R2QaNmO43OsR7FExsQhvbBOQF3dsKtpg3F7f7zFSQzFD
jx9KWlEZIAL0mTN4ZLvoyz/HOT6oRZVKF5BPs5laZ390opC6PxB+0mKXmsiBId14vgShau6JjQ+q
SsXFc5aMzkRvWCjG3kaRJ56owC0Z6ksAn9JRQlgj05XZJw3CmU1D4/lZ2gD0mY8SRLsaHGRomgz1
h7Hi/wTMvrgQIz2F6yHSKrM+B7lwefA+DHfp5hI3PipuFQVDV2t+WVfFa0ogQPAav/+t58FbPMKU
jWR5LWHvrZtDtaMgQewXuCLW4YzSXaKFbbou8BB+CbgJoopndwxZxuMl8ntSRFiNPV2sfHdD9CmQ
t0hzAOf1hLYqCvBzoJnckEvsS6iN35r8u+KSjhe7R8MA7bzyPXk+ULXqNdrrvrLGk6EXXBI3BJcf
O/etzb+YukPdL7kHL1nWrw+i8NOWg0U0rC0HCEu7b9v5jJnP2ly7V4S613SbBLjndfoeaUxJKPVC
RkDi0vNGSJETS4yjFCO9HA6ZaXp+sYAu0HTKxQi1LQOibD+AjWGnbdhMgPiRt5xUP/rT6Bv+1gdh
oW7ft44DVQ7P2r1w3/bRm/orD2BL6wfO230V2+SZ/yHNBtzvkVuMNtLxlKoPe24AWamo1/nFyCC1
CI20Cql0PZ+ZI+5VJQVUGrflLjx7r2xRLXgeqIS30/eyL5MvZJZSSti+aJxT/qVAPS1gMpKTKAzv
A4B1tdy+UkVlHm73SHUGQgKiYf7X2PXQdtI6zpwJTba75su58nx8LD7soX6yDxRg+kCFhbg2JWGE
bfA1YStg6dp+FmgF/iUlg3DMfih268eNY8HiNq67bfa52dmTe19t+2eUqOmJS82PVT8p41Aur3OX
W6O7nRCJiIv12CrWs60kXBUng+528aMRlEUXxq6F7dJh2BAAB04oq6XXJaXZsJN7Wj7x33W04rmu
mpGWKVZEblzJe/L26Rzt75ICC/K45Z75ZtkQcbBHp8Zv7GdtX1Jqek4562Q+s3+9IO405hdjB4BH
4fE1yba0lOzVcyzrgXyl8idLBcmyjn/N51UGLjzqFggdjdqPHmMktEyZ4bgUbd1h14zhtt0Wokuy
8lYfrjxmUjTMPibbOuOuZbMQ9iHWb/7VmPSrD8+IrNe7jsB9OFrxidM5lWE6W2VuI42bCs/xmPjx
ktqFliktA3FNRzELHRReGC5zpt8Umur/K8Oirl1bYl9davP6E18JsoMHvVtiisJsVorRz0/PZqD6
FQhGbo4JvUc6VbWXZ82BpQvohf7xWI39lQi+1iXop/fceuk+WK1DoS31hcX/7uRZ5OPJHLAvEpM4
cy9EKugcvV9RKPZTspETiUQ3jlFrMz9vvevUulhpkzaLUvphGLhJNfvgqBlm/Ksz/l3uG0ewcTi1
IDBnt5/v8uHtpZ66JRr+PMgd7Kabd74gZke/sp8DLDvXQx0qa45Ho2Ar/v8e1ZsHZ8xSXU9KXJeN
xXSx8wJcVcQKi6X7sK1RXHWmTRcz7Z3A+qORbV4AnwokegO0k3jbKVHwV3T9SguIqq+qjGo/Xtls
aTMr/wqw+LYvoEQw74dHYJXHuTA7cd+QMNfnicRgYp4pFn/n9x2SAWBs/hLdycjhUHaxJF93V8nT
fCxAksm8qzRaIvd5YYZs5WnMukdaJRHsC3LgU/V6bDa5fPZW6w9fj6PKjPdb+V9Nt/lVyVkJdc0H
WBM2h3ekDoLsiY0o2iY3b6srWkStJE3VQ84hGpJHxfu1r4VUJyvyKqxsCmY0DtBCv+I1HZmytcyD
4UnjzD28q8ZhhvSrkVyqAlsyDhzm2g8l1xCUkogfwJlUH9tSrSmiuvdJ6aU06JiT37wOiVv+rpiI
kSA6KxCuQ/0K9QvoPrxEp+QWogPdc4stdZKngFisZhapmFE90lRZ4CvkknDJ8jj3H3jkHmZdlfFT
kQ7HJJ6BqJTa02metcvqeHt4ln97yQmqoaXIMXlzJp5kQ2VS8NEVw/M6FgDW3ppmSzo8vhK/iOu2
960VKOd0LUlNz56yZkik/mi1y+9aIUUuTNyKnKTwyskQhQOxo0BcaznJY42VOP7YFNew25XkDKpq
EN6CGKfJmKs/V6jLYTINJmr5w5BCMQRFhuCZxkZQKErj15CSzgGD0V29Qf7oxYW/92kJRC4uENQf
1kvnmqNOefHRdhwH3hhOrh7587u9/bAiyji8SjDu98b1M2WlJ8KRfCXKqP6wboJaz6RscjYzY47L
oTBgCGrRP0mKADizyaztc0aicNhmdmG+bEoULjZLucAn4BczL+rreDzjrnHaprFtnsyZRvQlzWP/
N/y1oUeEGmNr1zFDdKBdnfDDasszzNDkJxISkfBoaKU8K0+nQySPzwgk1OH6JQfdylpKA1MtG+Eh
CWWlNwUTzhqxCLS477YWvjilvI30HhrkJgq86QGJEazMdgQN7EDyquAq/lKPOaiGHgsONFoM7FZ+
+pSdNLDWxLgEJ6ougI2IcMWo6pOhsPANXCn6NKOQoNCqn/M5zy/rCQffEaChq1fYYTmuDxIh0Abf
gwJ1bL6j5YGqc9pwHeJQKbgCd829fSZmhtPg14OcLYomZ+O5tfWXJjLDFvLK6VfsAyIf6uVZIg08
FdlYncjneFojxZDtlMrIYH8InMwfpvL0Q2siDFq5gzlVjNd4brLYLUdpgweHymUqKpM3kJUlVZuB
7WQMGkuudvHWthFPem5x0trh6c9IDE5GN2rDMrJlLxLgNCC/X+K+WxiQVOXK6/clw08jZgb73za3
RgvwvbPpFFBieWkMOej2VaDK0TWxLPYS27IvQJM+sGJEJAl8mgJoQWp0fuPrRFguKt0aewyMow0M
2KLxu3zJQPjyzjP7XqgNoFb7dhlYZ14/qt0uaM3P7Sz0EGZJjCn1FYMpZMrhm8W8KbuajJMIBQy+
ChKSaQWuKTofCjFDJi/cyfC69zsrlIQfJor13hLv4ABIfBx0eohFiCfsWxZxAYhD8tkIdXTImNFg
7+oz82oogwZWNES6qqlIPVqh73PVho+sG2qPmb8vCNGDuADMqesyOPxDz3Wn37sg2bu3cJz6vMmY
Cyr0oQ0s4K22zaLdAVkharfco2/Qh5CRKEmQDWnMDSoeg1y3R16srt0jRXk9XuM0A9P/+wv3061y
Vu1XaCuUvxLPw4iicBBBgFapEEVCMi16MaHgTLvs8xQeA1eCiK1xlsXLsDn/iNmQQ/VyzD20fDx0
wtw18gATBbnUtculicN6kdy7eJOAfJ3CSGSNl82+eDwxED/AJbFx923pdO4kaYL8wvn3inWJSsaV
uV/T4EiY+2/R+u53TNbtU5fStmWJuJIlba26JJt+ahSPaBKEd1iWktAbTKnDxkJh1k+Ig8Ch38TR
tEbUMSpDPTOWG+lBUwV9VNoxDc7eXM3umX/i4XUeEY5SAyqoie0el30HkOtuXzwa8UQiQ1XiKO6C
ShxmchxMQ5yCqqccqwq+UQPtstrzST17U8ziidreGKRAwRMhIGYFXZomfh2Ka6Vv30e1MqH6G6i0
aXzN8U+WiSHORKexWM/wsnefXHzss6OR6cmux+RsPDveQlnVm/v7qISmIFUqPXF11/nDObkhyihj
JESzjUHYNDJ7zc/ViomA29AE2l939NEfa4ue4sRPKrGThcGyrwoVjgdPIDsljte3bHSNr7iutyFO
W/GfvFb1whuC07ljiOUfsWHTmwPWU625OHcdkio8LRvQ6UhnDfM3b+SrUWJZlCOJ08TyUIzCMAZB
2/sjQKEYWtc3xkp0iOk5Lok53R9ZsA0xk+nB8Hjqh1UZVzAQPxA8zHVxV4v7oAvSCZQc0DRoHozB
f+Rm8lNQCSh/4Qtu+vjEy/QCfY7oF04doMERJEAfRXeIkDdPQgvANFCmqIJPxvuv36AWHVLuts4k
GdU77PW3rW50Vf7fdxy9qjZrbxQN8qq4INJ1DUdCk94uqNKD8j17YFfq2GXaaC4tYbyk2Tt5dROu
recdsHhUAuaK/qlHiYqGbkeJxC1kMLakgYjDBYisR/vVaGbFABHBfqxZGvsPv4yAiQXh189rGaR4
sxysDf7jrUeeD/Gmw2i3ulxomkUM3mKLd90QYUeVm2vkmyVpYWNMCkX7M3EY2fj8GSnLQ6ukfnc3
o40xnhy3OBq9o4NkOTJFez8hgVl9lcumJMKkR47nK9C3AZUUnUArbGqDHdHn3bknPoQcObVzy7pJ
Y3OGy2Z3THlfM1ha4bGV4m359V6A1BUODLv9eXP6YpGrWQjdJwsym+lkvD6vzfkMbcmtwQ8q5IyS
wFohmRe1Czg41oNFEjU1JdoT2eGLSZgje1xo/cJwDPLnAkbyfmjlVt3fupAgvNGeZS6SBMQmexIr
ELYcpaMsXzALi8sPSouEsRu0hIQRTRGnJjBx9K1Sr1UBckYRdie3tHx2yObuqb5EPnYAzqOuS5Dy
CJ6igb/AyNojHLtQePOGmeZWPrUhKPG02ckg4xriOI2CjTgM808IhoJEhpZI25UWnhVo999jeSRa
THfI1Tjf9D07Va+MFYC+kLBLNM7sNyZfCUXP12LqpkboqO8MSvo/NR2uopBNwozHjGt9TdcXhhKC
z2BicQZI0Z+Uq6wnD2kWn3ryCSsN+xCoIJPqUkdua8a0lnWFoDw7NdpRzEuPPnl0foaJRYieSVuX
JfDjco/LOODbsefaHx1C11rXrqh3xOg75dpbQIcKtSn9HEiUQ5In4lJXP2mqvunFHeqUbRKwWPuL
bXhH394MkVFYpcWBo5YzWNaCddd93vjvxpZCIzXdXCOgPjgcVPD84LFPcl41hap1I/d2USslCNMM
vEOgrFjY1ViiLYwC/PknL3L7E7xsPcm25nHl2r5oWuc1jafg2i6yI20O3a0PgZfNG5yy45TOU183
mpP5cFDKnqrqWhQ9T6CoAQPExXTAnChJvyyIdxSjWnX4/mZXG1lEHKhERg7kRzHVTKBWvn6uClXK
IqFa72SaaHubbebGgQapNhPoIusTbEXuqMWGhv3Qjd4egWYEweO1tOSd1O4pGSJuWoJwKRtP9iK6
rZij4MZBW8pZdtjGetIA9ARhuYUX27qUIcE5WtEJLXguE2LN/yrLs5Cz88S2jNKgH2VgM34yNkDg
XUal+Hv/vETdGC5t9EPXsLApqO0S7qsOfecrq50gbF1VKElEujG4b7m3YoABuyg9knhbpuyn6sy+
cMds3/P6B9nwI0TY8klQQtRaN1AVfszNOEBUDGIMhUxvcnty3leldl7n0Y6t/MurGrZ/CiVX1WyR
CK8x7Hwmdwp2yELCs1x/aQLVb8K5Aq8GhfzsZzIz+zwktO0sZPE5JutXqWe60vc1x57Y7gL/pKtT
cw/6yyo1zrbnsy8V3y0DOZ47QyBjGXQoVscQWY8//DP72JGayN2bkzcPuMd+A9hxySNg0wn7INgX
o3FEdvWRfZbo+i6J5Wgb7ksfcV6b1gFBjGyBXWutr8kty5hRBLKzDqgtdL4J6NqAl+vy5eU3nVgE
ljcn15ua8z/quDSjvuMSMz9AJupUqy3cCHqhbl5Pxn4cVkTCtBGFB0vbskwOHr1YOeulF/e50hTC
Zyu5sZc69phJhDs41bYfyje36xvLT9F9R6VlmrTWMih5PGa5PL0Ce5QMLVSvTekkmj5ua6MwDbU1
+k9elXiWSNGGprTXA7iDpNvgZAB4ePMtqyZ03/osvlRkPafyqktJJvZ6q0fW0gde3ULr7r106QtO
Sw1ZaP69fK6pD1lWFHmm7GdIZDM2pTR6x0tpPpWwrsUNEG+huasVNfzoLk42OulQ1ZNWJ7nh8c4I
VR/rBHF6WJynAm4WTgHKV5J4NuCeb46Shu0YazWVvQanm0bsDUjUf/CzpJMHiPVsrIYoQnh8WoLa
ADezoZZk4qzezH8lmrzzIbknRak6Mjs7MqySPr6hUuenW6HFNoKweZVDOeCh+chdNA+o/OUlsNRB
55IShRA6g+ZyOMp9wmu9pJt5Ixv1eAEyf6gr1pjx9x2bYvrAV07nVGMuHRcTSiVArvYoLp4XlYip
p3XxrVlqcvyFQt1p+9rItfO8+x6TkfJ4zVnVotYuq77Mf/BthJ059ATUtdpJIEx14+F7OPBlCaB2
aJ0eSBLGAqjUKoda6YTnFSeoP25dln+KkFUpDIneMxLmOWERt3LQ/FVmAHWIg7NY9QgHyn3IdMOQ
N8Nej/pxnJhV2CSI6MbYbx0QyPJAY3zyMvy/1ncey8TYtAqdPIkx8jL5/v+WLLwzbUzYNakELF2B
AvsUndOQlfI9YUFl4tFTypxuxoVXHws/4qUHwvXml27ku5kZFK/XDi5S793AQi343yac2vLiKwUJ
ZQAd0Gh10Zpco+UkWyYpOpV+8ErFAsODB43K54QADxAQ0C5bklWEOTyPVsjyvmkkD5oqVw2wpffu
vR+NzRXXZITvr9BQP+N6eXtSqGk0KOE76zwQ0K6Ot9thEne5rQM1XsLif09dIYwlFL/HYxv03E2R
B4sj9f/sO6YsU2myq0VeeEFzgb1+Ap28IbWB9kTTbPSiINPIcw8XfXCkftli8kN8T6WjJ0Xa8Np1
U1wUBODao8YVp9RiamlQBLaueqLhKCvrERrwz4YG2ASioI8A95n6iBsDn5oakN9p7hGG0aIvUUqv
4yI6Gp8TZaoe+7VSskax4iaLysos42z9lgYpYOI9zM9h6VidcDAbfeRBy0T9yLsALQIUiZHIAVsT
bd8+pGSUpghaeYZLVaVtYexokG0M8FuqTg/apoUqCqeYvBt8UPkU3QMjOKMs1o0ciX4aRhjIp85l
MU4sfVxcJkEMMyGuZoUhURd8imQ1VpxMrjnkhQH141PgO1A4C4dm0KqYBSbapNqZhSQt6o37LEFX
z8t6GriPlNON4zKFNCKoSLRZrPlcfHwJD1F1f9Bp0adwgbAZ4mdYU+IPYXzEK7/DwhlTYA6gfoLx
ulExkGTAFNQ4+baGqznmul/mZ9rTnDMOCJG2nDTWsfC3s9za1MnpyTeFEtw5sd54fHWgbArlYR6c
PosUJkgALeXKmQqNKnkGz+bFNM6njSYI+I+PQHHTxJoASPYBgT20WBnmeF1DKp5RsWvdzRxINz4E
w8N3Hq1mpDlarlu+TOcczuGupgJgUQkP94tEQC2zGXSFLkuin/FPAGbbRAGT0Z23R40pRApQoE86
a7JAOZQGhXNygHumt7cZdgVH6qrF58Niv5ZMiAk0m6WtrpAqqlVSkD+pBG35NIau2MW+3W9MfHQk
hq745b5MKIvJSoxyD3W1ysx+0If7mYlL/Cx7Q83pOwIp9wPvSTQDKPX3N6BWVUlgArC1tAE1Dt5A
2SNcJiTy2WCF/tpSrBxGFVGQ30YBvYuGu//SCszbA9vm0MlcBUGkdVyUi6MF7zHiOzPzJYe94FGG
my3ul7KhJXHM7Qw7ODxQlBuDsdtOaN+rrYPcJSObbSnkri4qzl0Rk5hGAzKII/Tjrr7v5aWP7aw4
eYwVYLjx7EgVEAY9Afv7tu+6vB/HR23Q9fRfGARsZxRunpSuBKqIhEjKfvxKKv2V8q93P4hS1VXy
MtwpqUtnkKp2+NL2+R3K51fF5fUPCCXXZlUKD/KCiz4m4ajOMVDYQbYRslWvICWhMIPriLqURyQo
4ky4McECekoPOfL24jztU40lyiFlSrAUUr50R0XHC3rUIfBUBbiBjKiGSdD9QQSyNrZoDStdKgdl
4joHwTokNXiX6CCHKKq0VDBTpubPfn64yoR+Hdltin1H30Tdi5IlR25liTBHQeehpRwNrKajx9Bo
TyipJdNNsSU1sLlPfCodgow2R5SkFZ9rK7iO3EAeEktKz1/BUVgf1Ma/M+7q4/CV5yThP7Hmrbld
wuZkoOEg0I/vrz6nkXMrx/twB9FhP2ZOZqTSvXybeMglrsAPSZnqrLUd7/XK+LAnkJmhnIeA+Y0P
XcUZyk6F6sSUj7oGsiZPhDGmV51YkdoXexzu1D/6ARdBMTybMzIudaX7nM2B2nMxyQ8QgvUlXFcg
ohUFFzICPBZADrjbpNPEdTSu1shb3egL7qcOT9fPxfk80gxnwjLM9XlM2fonGOaeEaN4ZDetGilC
pzJyoI8xNikHcCdA/gyA2a6tDARLytsLDG3cnYWCT8x9olJgVFhQj4ZH3n63WSveeg+/n7EARRzZ
3mdMX96SykyOgS/RKcw3bbiWarAJdbA3ud0nW8qJmN0mrJn80USDrdC8F5beRL3SI+iyXFpmah96
YBXw5XJm2CBCJl3wQz09ea3OAEHbDX3p9jtqZlSgrhx6HvoBYSyCuC1nfls39IRsPREGkmUU/pkZ
2TtIM9Vkn78T/pot3qepGGbo7lASzk6sW3OUljkKncmQKWt7r5bbeEc5MgENa9DOSqDJB86tzuI1
ZYcMSfHREeWPUR4JY1e5khkNShDiMmphgIQU0K2pi6NH0h6n0b6MHtsb/q6ubGwTFzGYgD0ptqxx
7tjE6FxRRbyTMdZW3ks6UeoONV3QS1uiTq2BIJ/iB8fXDxtVcbf10ZnpkCxgzUiA8IlB3QrEwlmv
aPXrKxKKtn03b5eoBhlJk7YxcYu7wuOA74EMwMKukaqxQz8hg4GuPHUjAY8f302xL37ulpRL9f49
EHSMEsoDIJLEB/q6xOWKFBra8DCA/p/yb9rOuNwRzWocXY/IUa+TFpHXfQg0YfguJFFbWGvTJtfx
60pkGkVGYRdjL3gN6HKZS5X+BA/1iI+ytUW4aH/SG/uJUE+FtrxdPgvf68lz/Jc8BtqyRglqXiBm
pss3iBrCUIDP3jDRbtEC9Sd5EKzN2p6BfwJBl2AdC2/8QyxiH8xMcGHE7TIWBNcMn0B7pWMhjtwu
6lureSRkGw4+AfepzoIl0Ym0B2A3oiAAlBCfmkkb/9HpWoUsDvudfyi5y9moIj0jCggKAeQ1UmA0
t+l3BVfrofIqrMeVFuLTHQItEhma/XVJfx0PbAi4Z3yiXbjj89Qlbq+wt7VdR9oQNwuQD0Dlw4RK
od+U0VOxtajNu6yUkj1OJJH1WsAlcFpLvTD8EtW7LEgmMPR129TCl7L68gID4UaCV9oj+ug08O6C
HZZ6B0mT/Npj4cjQ5MV4xzdBZyRVWaDf0W3amNBz+p/pZfgfbH/Gzvh8Lx0aieDvj9uGboQhwg4T
uWUcIBaa2/Bd1GH5pvcHtJHYnMn1Lwn5zxTubEApbKEZZPVwVx0OO8zqPVoH9ZE5p0V2jVkNFqev
olENC6ho2rbbv2tO4ALq4HDXrnLz11/qXgSM43ytvZDujlkjVmuFjC0wPo6T+SUL3JtHAcbLXet5
mHRio+5vXnLYfsPNJAdh2p4Bcn82mz/NebcxAt7SCkhFSsH8iwcBa8ocrKgJZcsbJryIamtNIcwb
W0g/Rp/fvmkvpRk5IKWJo6DDRIU7ISJa4pRw3jqFZrZT4juqx9p1bSEwAu/148Uy07NcHW/+8oJN
1t/xItLoMY/7Ba0Zth+1AYpdYzgRWy627ZummEMMoThOKfd6DZDR9CdV57Raga0vqdgs4hgIyYiS
0sN5M1xC8zJ0TJzIcps0nb1W6qePEqkHqKN2tiSQLCrOFeQChkotgQSSLcXu4rZ6aJeMgMWdWRZd
qfGwd0meRMX5TSbpZijz3XuTvEhBDypnU1PXQDEc67SwIic+okvpSDsDOzZcx8ync9eJnQW8KXwK
RchRGzqxZ6Nt8GDiU0Da7gkeo2ysoBiTfPQ73I0YjFnvYXoxYqYwYvPgMRs=
`pragma protect end_protected
