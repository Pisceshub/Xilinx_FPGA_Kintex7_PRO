
// XPIPE_quad0  ports
wire gt_refclk0;
wire  altclk_m;
wire [31:0] apb3prdata_m;
wire  apb3pready_m;
wire  apb3pslverr_m;
wire [15:0] apb3paddr_m;
wire  apb3clk_m;
wire axisclk_m;
wire  apb3penable_m;
wire  apb3presetn_m;
wire  apb3psel_m;
wire [31:0] apb3pwdata_m;
wire  apb3pwrite_m;
wire  bgbypassb_m;
wire  bgmonitorenb_m;
wire  bgpdb_m;
wire  bgrcalovrdenb_m;
wire [4:0] bgrcalovrd_m;
wire  scanclkb_m;
wire  scancntrlin_m;
wire  scanenb_m;
wire [3:0] scanin_m;
wire  scanrstb_m;
wire  xpscanclk_m;
wire  xpscanenb_m;
wire [15:0] xpscanin_m;
wire  xpscanmodeb_m;
wire  xpscanrstb_m;
wire  cssdrstb_m;
wire  cssdstopclk_m;
wire  edtupdateb_m;

wire  ch0_rxoutclk_m;
wire  ch0_txoutclk_m;
wire  ch0_bufgtce_m;
wire [3:0] ch0_bufgtcemask_m;
wire [11:0] ch0_bufgtdiv_m;
wire  ch0_bufgtrst_m;
wire [3:0] ch0_bufgtrstmask_m;
wire [31:0] ch0_dmonitorout_m;
wire  ch0_eyescandataerror_m;
wire  ch0_iloresetdone_m;
wire [15:0] ch0_pcsrsvdout_m;
wire [15:0] ch0_pinrsvdas_m;
wire  ch0_phyready_m;
wire  ch0_phystatus_m;
wire  ch0_resetexception_m;
wire [7:0] ch0_rx10gstat_m;
wire [2:0] ch0_rxbufstatus_m;
wire  ch0_rxbyteisaligned_m;
wire  ch0_rxbyterealign_m;
wire  ch0_rxcdrlock_m;
wire  ch0_rxcdrphdone_m;
wire  ch0_rxchanbondseq_m;
wire  ch0_rxchanisaligned_m;
wire  ch0_rxchanrealign_m;
wire [4:0] ch0_rxchbondo_m;
wire [1:0] ch0_rxclkcorcnt_m;
wire  ch0_rxcominitdet_m;
wire  ch0_rxcommadet_m;
wire  ch0_rxcomsasdet_m;
wire  ch0_rxcomwakedet_m;
wire [15:0] ch0_rxctrl0_m;
wire [15:0] ch0_rxctrl1_m;
wire [7:0] ch0_rxctrl2_m;
wire [7:0] ch0_rxctrl3_m;
wire [127:0] ch0_rxdata_m;
wire [7:0] ch0_rxdataextendrsvd_m;
wire [1:0] ch0_rxdatavalid_m;
wire  ch0_rxdccdone_m;
wire  ch0_rxdlyalignerr_m;
wire  ch0_rxdlyalignprog_m;
wire  ch0_rxelecidle_m;
wire  ch0_rxfinealigndone_m;
wire [5:0] ch0_rxheader_m;
wire [1:0] ch0_rxheadervalid_m;
wire  ch0_rxosintdone_m;
wire  ch0_rxosintstarted_m;
wire  ch0_rxosintstrobedone_m;
wire  ch0_rxosintstrobestarted_m;
wire  ch0_rxphaligndone_m;
wire  ch0_rxphalignerr_m;
wire  ch0_rxphdlyresetdone_m;
wire  ch0_rxphsetinitdone_m;
wire  ch0_rxphshift180done_m;
wire  ch0_rxpmaresetdone_m;
wire  ch0_rxprbserr_m;
wire  ch0_rxprbslocked_m;
wire  ch0_rxresetdone_m;
wire  ch0_rxsliderdy_m;
wire [1:0] ch0_rxstartofseq_m;
wire [2:0] ch0_rxstatus_m;
wire  ch0_rxsyncdone_m;
wire  ch0_rxvalid_m;
wire  ch0_tx10gstat_m;
wire [1:0] ch0_txbufstatus_m;
wire  ch0_txcomfinish_m;
wire  ch0_txdccdone_m;
wire  ch0_txdlyalignerr_m;
wire  ch0_txdlyalignprog_m;
wire  ch0_txphaligndone_m;
wire  ch0_txphalignerr_m;
wire  ch0_txphalignoutrsvd_m;
wire  ch0_txphdlyresetdone_m;
wire  ch0_txphshift180done_m;
wire  ch0_txpmaresetdone_m;
wire  ch0_txresetdone_m;
wire  ch0_txsyncdone_m;
wire  ch0_cdrbmcdrreq_m;
wire  ch0_cdrfreqos_m;
wire  ch0_cdrincpctrl_m;
wire  ch0_cdrstepdir_m;
wire  ch0_cdrstepsq_m;
wire  ch0_cdrstepsx_m;
wire  ch0_clkrsvd0_m;
wire  ch0_clkrsvd1_m;
wire  ch0_cssdrstb_m;
wire  ch0_cssdstopclk_m;
wire  ch0_edtupdateb_m;
wire  ch0_dmonfiforeset_m;
wire  ch0_dmonitorclk_m;
wire  ch0_eyescanreset_m;
wire  ch0_eyescantrigger_m;
wire [15:0] ch0_gtrsvd_m;
wire  ch0_gtrxreset_m;
wire  ch0_gttxreset_m;
wire  ch0_hsdppcsreset_m;
wire  ch0_iloreset_m;
wire  ch0_iloresetmask_m;
wire [2:0] ch0_loopback_m;
wire  ch0_pcierstb_m;
wire [15:0] ch0_pcsrsvdin_m;
wire  ch0_phyesmadaptsave_m;
wire  ch0_rxcdrhold_m;
wire  ch0_rxcdrovrden_m;
wire  ch0_rxcdrreset_m;
wire [4:0] ch0_rxchbondi_m;
wire  ch0_rxdapicodeovrden_m;
wire  ch0_rxdapicodereset_m;
wire  ch0_rxdlyalignreq_m;
wire  ch0_rxeqtraining_m;
wire  ch0_rxgearboxslip_m;
wire  ch0_rxlatclk_m;
wire  ch0_rxlpmen_m;
wire  ch0_rxmldchaindone_m;
wire  ch0_rxmldchainreq_m;
wire  ch0_rxmlfinealignreq_m;
wire  ch0_rxoobreset_m;
wire [4:0] ch0_rxpcsresetmask_m;
wire [1:0] ch0_rxpd_m;
wire  ch0_rxphalignreq_m;
wire [1:0] ch0_rxphalignresetmask_m;
wire  ch0_rxphdlypd_m;
wire  ch0_rxphdlyreset_m;
wire  ch0_rxphsetinitreq_m;
wire  ch0_rxphshift180_m;
wire [6:0] ch0_rxpmaresetmask_m;
wire  ch0_rxpolarity_m;
wire  ch0_rxprbscntreset_m;
wire [3:0] ch0_rxprbssel_m;
wire  ch0_rxprogdivreset_m;
wire [7:0] ch0_rxrate_m;
wire [1:0] ch0_rxresetmode_m;
wire  ch0_rxslide_m;
wire  ch0_rxsyncallin_m;
wire  ch0_rxtermination_m;
wire  ch0_rxuserrdy_m;
wire  ch0_rxusrclk_m;
wire [19:0] ch0_tstin_m;
wire  ch0_txcominit_m;
wire ch0_txphsetinitdone_m;
wire ch1_txphsetinitdone_m;
wire ch2_txphsetinitdone_m;
wire ch3_txphsetinitdone_m;
wire ch4_txphsetinitdone_m;
wire ch5_txphsetinitdone_m;
wire ch6_txphsetinitdone_m;
wire ch7_txphsetinitdone_m;
wire ch8_txphsetinitdone_m;
wire ch9_txphsetinitdone_m;
wire ch10_txphsetinitdone_m;
wire ch11_txphsetinitdone_m;
wire ch12_txphsetinitdone_m;
wire ch13_txphsetinitdone_m;
wire ch14_txphsetinitdone_m;
wire ch15_txphsetinitdone_m;

wire ch0_cfokovrdfinish_m;
wire ch1_cfokovrdfinish_m;
wire ch2_cfokovrdfinish_m;
wire ch3_cfokovrdfinish_m;
wire ch4_cfokovrdfinish_m;
wire ch5_cfokovrdfinish_m;
wire ch6_cfokovrdfinish_m;
wire ch7_cfokovrdfinish_m;
wire ch8_cfokovrdfinish_m;
wire ch9_cfokovrdfinish_m;
wire ch10_cfokovrdfinish_m;
wire ch11_cfokovrdfinish_m;
wire ch12_cfokovrdfinish_m;
wire ch13_cfokovrdfinish_m;
wire ch14_cfokovrdfinish_m;
wire ch15_cfokovrdfinish_m;

wire ch0_cfokovrdstart_m;
wire ch1_cfokovrdstart_m;
wire ch2_cfokovrdstart_m;
wire ch3_cfokovrdstart_m;
wire ch4_cfokovrdstart_m;
wire ch5_cfokovrdstart_m;
wire ch6_cfokovrdstart_m;
wire ch7_cfokovrdstart_m;
wire ch8_cfokovrdstart_m;
wire ch9_cfokovrdstart_m;
wire ch10_cfokovrdstart_m;
wire ch11_cfokovrdstart_m;
wire ch12_cfokovrdstart_m;
wire ch13_cfokovrdstart_m;
wire ch14_cfokovrdstart_m;
wire ch15_cfokovrdstart_m;

wire ch0_cfokovrdpulse_m;
wire ch1_cfokovrdpulse_m;
wire ch2_cfokovrdpulse_m;
wire ch3_cfokovrdpulse_m;
wire ch4_cfokovrdpulse_m;
wire ch5_cfokovrdpulse_m;
wire ch6_cfokovrdpulse_m;
wire ch7_cfokovrdpulse_m;
wire ch8_cfokovrdpulse_m;
wire ch9_cfokovrdpulse_m;
wire ch10_cfokovrdpulse_m;
wire ch11_cfokovrdpulse_m;
wire ch12_cfokovrdpulse_m;
wire ch13_cfokovrdpulse_m;
wire ch14_cfokovrdpulse_m;
wire ch15_cfokovrdpulse_m;

wire ch0_cfokovrdrdy0_m;
wire ch1_cfokovrdrdy0_m;
wire ch2_cfokovrdrdy0_m;
wire ch3_cfokovrdrdy0_m;
wire ch4_cfokovrdrdy0_m;
wire ch5_cfokovrdrdy0_m;
wire ch6_cfokovrdrdy0_m;
wire ch7_cfokovrdrdy0_m;
wire ch8_cfokovrdrdy0_m;
wire ch9_cfokovrdrdy0_m;
wire ch10_cfokovrdrdy0_m;
wire ch11_cfokovrdrdy0_m;
wire ch12_cfokovrdrdy0_m;
wire ch13_cfokovrdrdy0_m;
wire ch14_cfokovrdrdy0_m;
wire ch15_cfokovrdrdy0_m;

wire ch0_cfokovrdrdy1_m;
wire ch1_cfokovrdrdy1_m;
wire ch2_cfokovrdrdy1_m;
wire ch3_cfokovrdrdy1_m;
wire ch4_cfokovrdrdy1_m;
wire ch5_cfokovrdrdy1_m;
wire ch6_cfokovrdrdy1_m;
wire ch7_cfokovrdrdy1_m;
wire ch8_cfokovrdrdy1_m;
wire ch9_cfokovrdrdy1_m;
wire ch10_cfokovrdrdy1_m;
wire ch11_cfokovrdrdy1_m;
wire ch12_cfokovrdrdy1_m;
wire ch13_cfokovrdrdy1_m;
wire ch14_cfokovrdrdy1_m;
wire ch15_cfokovrdrdy1_m;
wire  ch0_txcomsas_m;
wire  ch0_txcomwake_m;
wire [15:0] ch0_txctrl0_m;
wire [15:0] ch0_txctrl1_m;
wire [7:0] ch0_txctrl2_m;
wire  ch0_txdapicodeovrden_m;
wire  ch0_txdapicodereset_m;
wire [127:0] ch0_txdata_m;
wire [7:0] ch0_txdataextendrsvd_m;
wire [1:0] ch0_txdeemph_m;
wire  ch0_txdetectrx_m;
wire [4:0] ch0_txdiffctrl_m;
wire  ch0_txdlyalignreq_m;
wire  ch0_txelecidle_m;
wire [5:0] ch0_txheader_m;
wire  ch0_txinhibit_m;
wire  ch0_txlatclk_m;
wire [6:0] ch0_txmaincursor_m;
wire [2:0] ch0_txmargin_m;
wire  ch0_txmldchaindone_m;
wire  ch0_txmldchainreq_m;
wire  ch0_txoneszeros_m;
wire  ch0_txpausedelayalign_m;
wire  ch0_txpcsresetmask_m;
wire [1:0] ch0_txpd_m;
wire  ch0_txphalignreq_m;
wire [1:0] ch0_txphalignresetmask_m;
wire  ch0_txphdlypd_m;
wire  ch0_txphdlyreset_m;
wire  ch0_txphdlytstclk_m;
wire  ch0_txphsetinitreq_m;
wire  ch0_txphshift180_m;
wire  ch0_txpicodeovrden_m;
wire  ch0_txpicodereset_m;
wire  ch0_txpippmen_m;
wire [4:0] ch0_txpippmstepsize_m;
wire  ch0_txpisopd_m;
wire [2:0] ch0_txpmaresetmask_m;
wire  ch0_txpolarity_m;
wire [4:0] ch0_txpostcursor_m;
wire  ch0_txprbsforceerr_m;
wire [3:0] ch0_txprbssel_m;
wire [4:0] ch0_txprecursor_m;
wire  ch0_txprogdivreset_m;
wire [7:0] ch0_txrate_m;
wire [1:0] ch0_txresetmode_m;
wire [6:0] ch0_txsequence_m;
wire  ch0_txswing_m;
wire  ch0_txsyncallin_m;
wire  ch0_txuserrdy_m;
wire  ch0_txusrclk_m;
wire  ch0_scanclkb_m;
wire  ch0_scancntrlin_m;
wire  ch0_scanenb_m;
wire [3:0] ch0_scanin_m;
wire  ch0_scanrstb_m;

wire  ch1_bufgtce_m;
wire [3:0] ch1_bufgtcemask_m;
wire [11:0] ch1_bufgtdiv_m;
wire  ch1_bufgtrst_m;
wire [3:0] ch1_bufgtrstmask_m;
wire [31:0] ch1_dmonitorout_m;
wire  ch1_eyescandataerror_m;
wire  ch1_iloresetdone_m;
wire [15:0] ch1_pcsrsvdout_m;
wire [15:0] ch1_pinrsvdas_m;
wire  ch1_phyready_m;
wire  ch1_phystatus_m;
wire  ch1_resetexception_m;
wire [7:0] ch1_rx10gstat_m;
wire [2:0] ch1_rxbufstatus_m;
wire  ch1_rxbyteisaligned_m;
wire  ch1_rxbyterealign_m;
wire  ch1_rxcdrlock_m;
wire  ch1_rxcdrphdone_m;
wire  ch1_rxchanbondseq_m;
wire  ch1_rxchanisaligned_m;
wire  ch1_rxchanrealign_m;
wire [4:0] ch1_rxchbondo_m;
wire [1:0] ch1_rxclkcorcnt_m;
wire  ch1_rxcominitdet_m;
wire  ch1_rxcommadet_m;
wire  ch1_rxcomsasdet_m;
wire  ch1_rxcomwakedet_m;
wire [15:0] ch1_rxctrl0_m;
wire [15:0] ch1_rxctrl1_m;
wire [7:0] ch1_rxctrl2_m;
wire [7:0] ch1_rxctrl3_m;
wire [127:0] ch1_rxdata_m;
wire [7:0] ch1_rxdataextendrsvd_m;
wire [1:0] ch1_rxdatavalid_m;
wire  ch1_rxdccdone_m;
wire  ch1_rxdlyalignerr_m;
wire  ch1_rxdlyalignprog_m;
wire  ch1_rxelecidle_m;
wire  ch1_rxfinealigndone_m;
wire [5:0] ch1_rxheader_m;
wire [1:0] ch1_rxheadervalid_m;
wire  ch1_rxosintdone_m;
wire  ch1_rxosintstarted_m;
wire  ch1_rxosintstrobedone_m;
wire  ch1_rxosintstrobestarted_m;
wire  ch1_rxphaligndone_m;
wire  ch1_rxphalignerr_m;
wire  ch1_rxphdlyresetdone_m;
wire  ch1_rxphsetinitdone_m;
wire  ch1_rxphshift180done_m;
wire  ch1_rxpmaresetdone_m;
wire  ch1_rxprbserr_m;
wire  ch1_rxprbslocked_m;
wire  ch1_rxresetdone_m;
wire  ch1_rxsliderdy_m;
wire [1:0] ch1_rxstartofseq_m;
wire [2:0] ch1_rxstatus_m;
wire  ch1_rxsyncdone_m;
wire  ch1_rxvalid_m;
wire  ch1_tx10gstat_m;
wire [1:0] ch1_txbufstatus_m;
wire  ch1_txcomfinish_m;
wire  ch1_txdccdone_m;
wire  ch1_txdlyalignerr_m;
wire  ch1_txdlyalignprog_m;
wire  ch1_txphaligndone_m;
wire  ch1_txphalignerr_m;
wire  ch1_txphalignoutrsvd_m;
wire  ch1_txphdlyresetdone_m;
wire  ch1_txphshift180done_m;
wire  ch1_txpmaresetdone_m;
wire  ch1_txresetdone_m;
wire  ch1_txsyncdone_m;
wire  ch1_cdrbmcdrreq_m;
wire  ch1_cdrfreqos_m;
wire  ch1_cdrincpctrl_m;
wire  ch1_cdrstepdir_m;
wire  ch1_cdrstepsq_m;
wire  ch1_cdrstepsx_m;
wire  ch1_clkrsvd0_m;
wire  ch1_clkrsvd1_m;
wire  ch1_cssdrstb_m;
wire  ch1_cssdstopclk_m;
wire  ch1_edtupdateb_m;
wire  ch1_dmonfiforeset_m;
wire  ch1_dmonitorclk_m;
wire  ch1_eyescanreset_m;
wire  ch1_eyescantrigger_m;
wire [15:0] ch1_gtrsvd_m;
wire  ch1_gtrxreset_m;
wire  ch1_gttxreset_m;
wire  ch1_hsdppcsreset_m;
wire  ch1_iloreset_m;
wire  ch1_iloresetmask_m;
wire [2:0] ch1_loopback_m;
wire  ch1_pcierstb_m;
wire [15:0] ch1_pcsrsvdin_m;
wire  ch1_phyesmadaptsave_m;
wire  ch1_rxcdrhold_m;
wire  ch1_rxcdrovrden_m;
wire  ch1_rxcdrreset_m;
wire [4:0] ch1_rxchbondi_m;
wire  ch1_rxdapicodeovrden_m;
wire  ch1_rxdapicodereset_m;
wire  ch1_rxdlyalignreq_m;
wire  ch1_rxeqtraining_m;
wire  ch1_rxgearboxslip_m;
wire  ch1_rxlatclk_m;
wire  ch1_rxlpmen_m;
wire  ch1_rxmldchaindone_m;
wire  ch1_rxmldchainreq_m;
wire  ch1_rxmlfinealignreq_m;
wire  ch1_rxoobreset_m;
wire [4:0] ch1_rxpcsresetmask_m;
wire [1:0] ch1_rxpd_m;
wire  ch1_rxphalignreq_m;
wire [1:0] ch1_rxphalignresetmask_m;
wire  ch1_rxphdlypd_m;
wire  ch1_rxphdlyreset_m;
wire  ch1_rxphsetinitreq_m;
wire  ch1_rxphshift180_m;
wire [6:0] ch1_rxpmaresetmask_m;
wire  ch1_rxpolarity_m;
wire  ch1_rxprbscntreset_m;
wire [3:0] ch1_rxprbssel_m;
wire  ch1_rxprogdivreset_m;
wire [7:0] ch1_rxrate_m;
wire [1:0] ch1_rxresetmode_m;
wire  ch1_rxslide_m;
wire  ch1_rxsyncallin_m;
wire  ch1_rxtermination_m;
wire  ch1_rxuserrdy_m;
wire  ch1_rxusrclk_m;
wire [19:0] ch1_tstin_m;
wire  ch1_txcominit_m;
wire  ch1_txcomsas_m;
wire  ch1_txcomwake_m;
wire [15:0] ch1_txctrl0_m;
wire [15:0] ch1_txctrl1_m;
wire [7:0] ch1_txctrl2_m;
wire  ch1_txdapicodeovrden_m;
wire  ch1_txdapicodereset_m;
wire [127:0] ch1_txdata_m;
wire [7:0] ch1_txdataextendrsvd_m;
wire [1:0] ch1_txdeemph_m;
wire  ch1_txdetectrx_m;
wire [4:0] ch1_txdiffctrl_m;
wire  ch1_txdlyalignreq_m;
wire  ch1_txelecidle_m;
wire [5:0] ch1_txheader_m;
wire  ch1_txinhibit_m;
wire  ch1_txlatclk_m;
wire [6:0] ch1_txmaincursor_m;
wire [2:0] ch1_txmargin_m;
wire  ch1_txmldchaindone_m;
wire  ch1_txmldchainreq_m;
wire  ch1_txoneszeros_m;
wire  ch1_txpausedelayalign_m;
wire  ch1_txpcsresetmask_m;
wire [1:0] ch1_txpd_m;
wire  ch1_txphalignreq_m;
wire [1:0] ch1_txphalignresetmask_m;
wire  ch1_txphdlypd_m;
wire  ch1_txphdlyreset_m;
wire  ch1_txphdlytstclk_m;
wire  ch1_txphsetinitreq_m;
wire  ch1_txphshift180_m;
wire  ch1_txpicodeovrden_m;
wire  ch1_txpicodereset_m;
wire  ch1_txpippmen_m;
wire [4:0] ch1_txpippmstepsize_m;
wire  ch1_txpisopd_m;
wire [2:0] ch1_txpmaresetmask_m;
wire  ch1_txpolarity_m;
wire [4:0] ch1_txpostcursor_m;
wire  ch1_txprbsforceerr_m;
wire [3:0] ch1_txprbssel_m;
wire [4:0] ch1_txprecursor_m;
wire  ch1_txprogdivreset_m;
wire [7:0] ch1_txrate_m;
wire [1:0] ch1_txresetmode_m;
wire [6:0] ch1_txsequence_m;
wire  ch1_txswing_m;
wire  ch1_txsyncallin_m;
wire  ch1_txuserrdy_m;
wire  ch1_txusrclk_m;
wire  ch1_scanclkb_m;
wire  ch1_scancntrlin_m;
wire  ch1_scanenb_m;
wire [3:0] ch1_scanin_m;
wire  ch1_scanrstb_m;

wire  ch2_bufgtce_m;
wire [3:0] ch2_bufgtcemask_m;
wire [11:0] ch2_bufgtdiv_m;
wire  ch2_bufgtrst_m;
wire [3:0] ch2_bufgtrstmask_m;
wire [31:0] ch2_dmonitorout_m;
wire  ch2_eyescandataerror_m;
wire  ch2_iloresetdone_m;
wire [15:0] ch2_pcsrsvdout_m;
wire [15:0] ch2_pinrsvdas_m;
wire  ch2_phyready_m;
wire  ch2_phystatus_m;
wire  ch2_resetexception_m;
wire [7:0] ch2_rx10gstat_m;
wire [2:0] ch2_rxbufstatus_m;
wire  ch2_rxbyteisaligned_m;
wire  ch2_rxbyterealign_m;
wire  ch2_rxcdrlock_m;
wire  ch2_rxcdrphdone_m;
wire  ch2_rxchanbondseq_m;
wire  ch2_rxchanisaligned_m;
wire  ch2_rxchanrealign_m;
wire [4:0] ch2_rxchbondo_m;
wire [1:0] ch2_rxclkcorcnt_m;
wire  ch2_rxcominitdet_m;
wire  ch2_rxcommadet_m;
wire  ch2_rxcomsasdet_m;
wire  ch2_rxcomwakedet_m;
wire [15:0] ch2_rxctrl0_m;
wire [15:0] ch2_rxctrl1_m;
wire [7:0] ch2_rxctrl2_m;
wire [7:0] ch2_rxctrl3_m;
wire [127:0] ch2_rxdata_m;
wire [7:0] ch2_rxdataextendrsvd_m;
wire [1:0] ch2_rxdatavalid_m;
wire  ch2_rxdccdone_m;
wire  ch2_rxdlyalignerr_m;
wire  ch2_rxdlyalignprog_m;
wire  ch2_rxelecidle_m;
wire  ch2_rxfinealigndone_m;
wire [5:0] ch2_rxheader_m;
wire [1:0] ch2_rxheadervalid_m;
wire  ch2_rxosintdone_m;
wire  ch2_rxosintstarted_m;
wire  ch2_rxosintstrobedone_m;
wire  ch2_rxosintstrobestarted_m;
wire  ch2_rxphaligndone_m;
wire  ch2_rxphalignerr_m;
wire  ch2_rxphdlyresetdone_m;
wire  ch2_rxphsetinitdone_m;
wire  ch2_rxphshift180done_m;
wire  ch2_rxpmaresetdone_m;
wire  ch2_rxprbserr_m;
wire  ch2_rxprbslocked_m;
wire  ch2_rxresetdone_m;
wire  ch2_rxsliderdy_m;
wire [1:0] ch2_rxstartofseq_m;
wire [2:0] ch2_rxstatus_m;
wire  ch2_rxsyncdone_m;
wire  ch2_rxvalid_m;
wire  ch2_tx10gstat_m;
wire [1:0] ch2_txbufstatus_m;
wire  ch2_txcomfinish_m;
wire  ch2_txdccdone_m;
wire  ch2_txdlyalignerr_m;
wire  ch2_txdlyalignprog_m;
wire  ch2_txphaligndone_m;
wire  ch2_txphalignerr_m;
wire  ch2_txphalignoutrsvd_m;
wire  ch2_txphdlyresetdone_m;
wire  ch2_txphshift180done_m;
wire  ch2_txpmaresetdone_m;
wire  ch2_txresetdone_m;
wire  ch2_txsyncdone_m;
wire  ch2_cdrbmcdrreq_m;
wire  ch2_cdrfreqos_m;
wire  ch2_cdrincpctrl_m;
wire  ch2_cdrstepdir_m;
wire  ch2_cdrstepsq_m;
wire  ch2_cdrstepsx_m;
wire  ch2_clkrsvd0_m;
wire  ch2_clkrsvd1_m;
wire  ch2_cssdrstb_m;
wire  ch2_cssdstopclk_m;
wire  ch2_edtupdateb_m;
wire  ch2_dmonfiforeset_m;
wire  ch2_dmonitorclk_m;
wire  ch2_eyescanreset_m;
wire  ch2_eyescantrigger_m;
wire [15:0] ch2_gtrsvd_m;
wire  ch2_gtrxreset_m;
wire  ch2_gttxreset_m;
wire  ch2_hsdppcsreset_m;
wire  ch2_iloreset_m;
wire  ch2_iloresetmask_m;
wire [2:0] ch2_loopback_m;
wire  ch2_pcierstb_m;
wire [15:0] ch2_pcsrsvdin_m;
wire  ch2_phyesmadaptsave_m;
wire  ch2_rxcdrhold_m;
wire  ch2_rxcdrovrden_m;
wire  ch2_rxcdrreset_m;
wire [4:0] ch2_rxchbondi_m;
wire  ch2_rxdapicodeovrden_m;
wire  ch2_rxdapicodereset_m;
wire  ch2_rxdlyalignreq_m;
wire  ch2_rxeqtraining_m;
wire  ch2_rxgearboxslip_m;
wire  ch2_rxlatclk_m;
wire  ch2_rxlpmen_m;
wire  ch2_rxmldchaindone_m;
wire  ch2_rxmldchainreq_m;
wire  ch2_rxmlfinealignreq_m;
wire  ch2_rxoobreset_m;
wire [4:0] ch2_rxpcsresetmask_m;
wire [1:0] ch2_rxpd_m;
wire  ch2_rxphalignreq_m;
wire [1:0] ch2_rxphalignresetmask_m;
wire  ch2_rxphdlypd_m;
wire  ch2_rxphdlyreset_m;
wire  ch2_rxphsetinitreq_m;
wire  ch2_rxphshift180_m;
wire [6:0] ch2_rxpmaresetmask_m;
wire  ch2_rxpolarity_m;
wire  ch2_rxprbscntreset_m;
wire [3:0] ch2_rxprbssel_m;
wire  ch2_rxprogdivreset_m;
wire [7:0] ch2_rxrate_m;
wire [1:0] ch2_rxresetmode_m;
wire  ch2_rxslide_m;
wire  ch2_rxsyncallin_m;
wire  ch2_rxtermination_m;
wire  ch2_rxuserrdy_m;
wire  ch2_rxusrclk_m;
wire [19:0] ch2_tstin_m;
wire  ch2_txcominit_m;
wire  ch2_txcomsas_m;
wire  ch2_txcomwake_m;
wire [15:0] ch2_txctrl0_m;
wire [15:0] ch2_txctrl1_m;
wire [7:0] ch2_txctrl2_m;
wire  ch2_txdapicodeovrden_m;
wire  ch2_txdapicodereset_m;
wire [127:0] ch2_txdata_m;
wire [7:0] ch2_txdataextendrsvd_m;
wire [1:0] ch2_txdeemph_m;
wire  ch2_txdetectrx_m;
wire [4:0] ch2_txdiffctrl_m;
wire  ch2_txdlyalignreq_m;
wire  ch2_txelecidle_m;
wire [5:0] ch2_txheader_m;
wire  ch2_txinhibit_m;
wire  ch2_txlatclk_m;
wire [6:0] ch2_txmaincursor_m;
wire [2:0] ch2_txmargin_m;
wire  ch2_txmldchaindone_m;
wire  ch2_txmldchainreq_m;
wire  ch2_txoneszeros_m;
wire  ch2_txpausedelayalign_m;
wire  ch2_txpcsresetmask_m;
wire [1:0] ch2_txpd_m;
wire  ch2_txphalignreq_m;
wire [1:0] ch2_txphalignresetmask_m;
wire  ch2_txphdlypd_m;
wire  ch2_txphdlyreset_m;
wire  ch2_txphdlytstclk_m;
wire  ch2_txphsetinitreq_m;
wire  ch2_txphshift180_m;
wire  ch2_txpicodeovrden_m;
wire  ch2_txpicodereset_m;
wire  ch2_txpippmen_m;
wire [4:0] ch2_txpippmstepsize_m;
wire  ch2_txpisopd_m;
wire [2:0] ch2_txpmaresetmask_m;
wire  ch2_txpolarity_m;
wire [4:0] ch2_txpostcursor_m;
wire  ch2_txprbsforceerr_m;
wire [3:0] ch2_txprbssel_m;
wire [4:0] ch2_txprecursor_m;
wire  ch2_txprogdivreset_m;
wire [7:0] ch2_txrate_m;
wire [1:0] ch2_txresetmode_m;
wire [6:0] ch2_txsequence_m;
wire  ch2_txswing_m;
wire  ch2_txsyncallin_m;
wire  ch2_txuserrdy_m;
wire  ch2_txusrclk_m;
wire  ch2_scanclkb_m;
wire  ch2_scancntrlin_m;
wire  ch2_scanenb_m;
wire [3:0] ch2_scanin_m;
wire  ch2_scanrstb_m;

wire  ch3_bufgtce_m;
wire [3:0] ch3_bufgtcemask_m;
wire [11:0] ch3_bufgtdiv_m;
wire  ch3_bufgtrst_m;
wire [3:0] ch3_bufgtrstmask_m;
wire [31:0] ch3_dmonitorout_m;
wire  ch3_eyescandataerror_m;
wire  ch3_iloresetdone_m;
wire [15:0] ch3_pcsrsvdout_m;
wire [15:0] ch3_pinrsvdas_m;
wire  ch3_phyready_m;
wire  ch3_phystatus_m;
wire  ch3_resetexception_m;
wire [7:0] ch3_rx10gstat_m;
wire [2:0] ch3_rxbufstatus_m;
wire  ch3_rxbyteisaligned_m;
wire  ch3_rxbyterealign_m;
wire  ch3_rxcdrlock_m;
wire  ch3_rxcdrphdone_m;
wire  ch3_rxchanbondseq_m;
wire  ch3_rxchanisaligned_m;
wire  ch3_rxchanrealign_m;
wire [4:0] ch3_rxchbondo_m;
wire [1:0] ch3_rxclkcorcnt_m;
wire  ch3_rxcominitdet_m;
wire  ch3_rxcommadet_m;
wire  ch3_rxcomsasdet_m;
wire  ch3_rxcomwakedet_m;
wire [15:0] ch3_rxctrl0_m;
wire [15:0] ch3_rxctrl1_m;
wire [7:0] ch3_rxctrl2_m;
wire [7:0] ch3_rxctrl3_m;
wire [127:0] ch3_rxdata_m;
wire [7:0] ch3_rxdataextendrsvd_m;
wire [1:0] ch3_rxdatavalid_m;
wire  ch3_rxdccdone_m;
wire  ch3_rxdlyalignerr_m;
wire  ch3_rxdlyalignprog_m;
wire  ch3_rxelecidle_m;
wire  ch3_rxfinealigndone_m;
wire [5:0] ch3_rxheader_m;
wire [1:0] ch3_rxheadervalid_m;
wire  ch3_rxosintdone_m;
wire  ch3_rxosintstarted_m;
wire  ch3_rxosintstrobedone_m;
wire  ch3_rxosintstrobestarted_m;
wire  ch3_rxphaligndone_m;
wire  ch3_rxphalignerr_m;
wire  ch3_rxphdlyresetdone_m;
wire  ch3_rxphsetinitdone_m;
wire  ch3_rxphshift180done_m;
wire  ch3_rxpmaresetdone_m;
wire  ch3_rxprbserr_m;
wire  ch3_rxprbslocked_m;
wire  ch3_rxresetdone_m;
wire  ch3_rxsliderdy_m;
wire [1:0] ch3_rxstartofseq_m;
wire [2:0] ch3_rxstatus_m;
wire  ch3_rxsyncdone_m;
wire  ch3_rxvalid_m;
wire  ch3_tx10gstat_m;
wire [1:0] ch3_txbufstatus_m;
wire  ch3_txcomfinish_m;
wire  ch3_txdccdone_m;
wire  ch3_txdlyalignerr_m;
wire  ch3_txdlyalignprog_m;
wire  ch3_txphaligndone_m;
wire  ch3_txphalignerr_m;
wire  ch3_txphalignoutrsvd_m;
wire  ch3_txphdlyresetdone_m;
wire  ch3_txphshift180done_m;
wire  ch3_txpmaresetdone_m;
wire  ch3_txresetdone_m;
wire  ch3_txsyncdone_m;
wire  ch3_cdrbmcdrreq_m;
wire  ch3_cdrfreqos_m;
wire  ch3_cdrincpctrl_m;
wire  ch3_cdrstepdir_m;
wire  ch3_cdrstepsq_m;
wire  ch3_cdrstepsx_m;
wire  ch3_clkrsvd0_m;
wire  ch3_clkrsvd1_m;
wire  ch3_cssdrstb_m;
wire  ch3_cssdstopclk_m;
wire  ch3_edtupdateb_m;
wire  ch3_dmonfiforeset_m;
wire  ch3_dmonitorclk_m;
wire  ch3_eyescanreset_m;
wire  ch3_eyescantrigger_m;
wire [15:0] ch3_gtrsvd_m;
wire  ch3_gtrxreset_m;
wire  ch3_gttxreset_m;
wire  ch3_hsdppcsreset_m;
wire  ch3_iloreset_m;
wire  ch3_iloresetmask_m;
wire [2:0] ch3_loopback_m;
wire  ch3_pcierstb_m;
wire [15:0] ch3_pcsrsvdin_m;
wire  ch3_phyesmadaptsave_m;
wire  ch3_rxcdrhold_m;
wire  ch3_rxcdrovrden_m;
wire  ch3_rxcdrreset_m;
wire [4:0] ch3_rxchbondi_m;
wire  ch3_rxdapicodeovrden_m;
wire  ch3_rxdapicodereset_m;
wire  ch3_rxdlyalignreq_m;
wire  ch3_rxeqtraining_m;
wire  ch3_rxgearboxslip_m;
wire  ch3_rxlatclk_m;
wire  ch3_rxlpmen_m;
wire  ch3_rxmldchaindone_m;
wire  ch3_rxmldchainreq_m;
wire  ch3_rxmlfinealignreq_m;
wire  ch3_rxoobreset_m;
wire [4:0] ch3_rxpcsresetmask_m;
wire [1:0] ch3_rxpd_m;
wire  ch3_rxphalignreq_m;
wire [1:0] ch3_rxphalignresetmask_m;
wire  ch3_rxphdlypd_m;
wire  ch3_rxphdlyreset_m;
wire  ch3_rxphsetinitreq_m;
wire  ch3_rxphshift180_m;
wire [6:0] ch3_rxpmaresetmask_m;
wire  ch3_rxpolarity_m;
wire  ch3_rxprbscntreset_m;
wire [3:0] ch3_rxprbssel_m;
wire  ch3_rxprogdivreset_m;
wire [7:0] ch3_rxrate_m;
wire [1:0] ch3_rxresetmode_m;
wire  ch3_rxslide_m;
wire  ch3_rxsyncallin_m;
wire  ch3_rxtermination_m;
wire  ch3_rxuserrdy_m;
wire  ch3_rxusrclk_m;
wire [19:0] ch3_tstin_m;
wire  ch3_txcominit_m;
wire  ch3_txcomsas_m;
wire  ch3_txcomwake_m;
wire [15:0] ch3_txctrl0_m;
wire [15:0] ch3_txctrl1_m;
wire [7:0] ch3_txctrl2_m;
wire  ch3_txdapicodeovrden_m;
wire  ch3_txdapicodereset_m;
wire [127:0] ch3_txdata_m;
wire [7:0] ch3_txdataextendrsvd_m;
wire [1:0] ch3_txdeemph_m;
wire  ch3_txdetectrx_m;
wire [4:0] ch3_txdiffctrl_m;
wire  ch3_txdlyalignreq_m;
wire  ch3_txelecidle_m;
wire [5:0] ch3_txheader_m;
wire  ch3_txinhibit_m;
wire  ch3_txlatclk_m;
wire [6:0] ch3_txmaincursor_m;
wire [2:0] ch3_txmargin_m;
wire  ch3_txmldchaindone_m;
wire  ch3_txmldchainreq_m;
wire  ch3_txoneszeros_m;
wire  ch3_txpausedelayalign_m;
wire  ch3_txpcsresetmask_m;
wire [1:0] ch3_txpd_m;
wire  ch3_txphalignreq_m;
wire [1:0] ch3_txphalignresetmask_m;
wire  ch3_txphdlypd_m;
wire  ch3_txphdlyreset_m;
wire  ch3_txphdlytstclk_m;
wire  ch3_txphsetinitreq_m;
wire  ch3_txphshift180_m;
wire  ch3_txpicodeovrden_m;
wire  ch3_txpicodereset_m;
wire  ch3_txpippmen_m;
wire [4:0] ch3_txpippmstepsize_m;
wire  ch3_txpisopd_m;
wire [2:0] ch3_txpmaresetmask_m;
wire  ch3_txpolarity_m;
wire [4:0] ch3_txpostcursor_m;
wire  ch3_txprbsforceerr_m;
wire [3:0] ch3_txprbssel_m;
wire [4:0] ch3_txprecursor_m;
wire  ch3_txprogdivreset_m;
wire [7:0] ch3_txrate_m;
wire [1:0] ch3_txresetmode_m;
wire [6:0] ch3_txsequence_m;
wire  ch3_txswing_m;
wire  ch3_txsyncallin_m;
wire  ch3_txuserrdy_m;
wire  ch3_txusrclk_m;
wire  ch3_scanclkb_m;
wire  ch3_scancntrlin_m;
wire  ch3_scanenb_m;
wire [3:0] ch3_scanin_m;
wire  ch3_scanrstb_m;

wire  correcterr_m;
wire [31:0] ctrlrsvdout_m;
wire [15:0] debugtracetdata_m;
wire  debugtracetvalid_m;
wire  uncorrecterr_m;
wire  xpipe_bufgtce_m;
wire [15:0] gpo_m;
wire  gtpowergood_m;
wire  hsclk0_lcpllfbclklost_m;
wire  hsclk0_lcplllock_m;
wire  hsclk0_lcpllrefclklost_m;
wire  hsclk0_lcpllrefclkmonitor_m;
wire [7:0] hsclk0_lcpllrsvdout_m;
wire  hsclk0_rpllfbclklost_m;
wire  hsclk0_rplllock_m;
wire  hsclk0_rpllrefclklost_m;
wire  hsclk0_rpllrefclkmonitor_m;
wire [7:0] hsclk0_rpllrsvdout_m;
wire  hsclk1_lcpllfbclklost_m;
wire  hsclk1_lcplllock_m;
wire  hsclk1_lcpllrefclklost_m;
wire  hsclk1_lcpllrefclkmonitor_m;

wire [7:0] hsclk1_lcpllrsvdout_m;
wire  hsclk1_rpllfbclklost_m;
wire  hsclk1_rplllock_m;
wire  hsclk1_rpllrefclklost_m;
wire  hsclk1_rpllrefclkmonitor_m;
wire [7:0] hsclk1_rpllrsvdout_m;
wire [15:0] ctrlrsvdin0_m;
wire [13:0] ctrlrsvdin1_m;
wire  debugtraceclk_m;
wire  debugtracetready_m;
wire [15:0] gpi_m;
wire  hsclk0_lcpllclkrsvd0_m;
wire  hsclk0_lcpllclkrsvd1_m;
wire [7:0] hsclk0_lcpllfbdiv_m;
wire  hsclk0_lcpllpd_m;
wire [2:0] hsclk0_lcpllrefclksel_m;
wire  hsclk0_lcpllreset_m;
wire  hsclk0_lcpllresetbypassmode_m;
wire [1:0] hsclk0_lcpllresetmask_m;
wire [7:0] hsclk0_lcpllrsvd0_m;
wire [7:0] hsclk0_lcpllrsvd1_m;
wire [25:0] hsclk0_lcpllsdmdata_m;
wire  hsclk0_lcpllsdmtoggle_m;
wire  hsclk0_rpllclkrsvd0_m;
wire  hsclk0_rpllclkrsvd1_m;
wire [7:0] hsclk0_rpllfbdiv_m;
wire  hsclk0_rpllpd_m;
wire [2:0] hsclk0_rpllrefclksel_m;
wire  hsclk0_rpllreset_m;
wire  hsclk0_rpllresetbypassmode_m;
wire [1:0] hsclk0_rpllresetmask_m;
wire [7:0] hsclk0_rpllrsvd0_m;
wire [7:0] hsclk0_rpllrsvd1_m;
wire [25:0] hsclk0_rpllsdmdata_m;
wire  hsclk0_rpllsdmtoggle_m;
wire  hsclk1_lcpllclkrsvd0_m;
wire  hsclk1_lcpllclkrsvd1_m;
wire [7:0] hsclk1_lcpllfbdiv_m;
wire  hsclk1_lcpllpd_m;
wire [2:0] hsclk1_lcpllrefclksel_m;
wire  hsclk1_lcpllreset_m;
wire  hsclk1_lcpllresetbypassmode_m;
wire [1:0] hsclk1_lcpllresetmask_m;
wire [7:0] hsclk1_lcpllrsvd0_m;
wire [7:0] hsclk1_lcpllrsvd1_m;
wire [25:0] hsclk1_lcpllsdmdata_m;
wire  hsclk1_lcpllsdmtoggle_m;
wire  hsclk1_rpllclkrsvd0_m;
wire  hsclk1_rpllclkrsvd1_m;
wire [7:0] hsclk1_rpllfbdiv_m;
wire  hsclk1_rpllpd_m;
wire [2:0] hsclk1_rpllrefclksel_m;
wire  hsclk1_rpllreset_m;
wire  hsclk1_rpllresetbypassmode_m;
wire [1:0] hsclk1_rpllresetmask_m;
wire [7:0] hsclk1_rpllrsvd0_m;
wire [7:0] hsclk1_rpllrsvd1_m;
wire [25:0] hsclk1_rpllsdmdata_m;
wire  hsclk1_rpllsdmtoggle_m;
wire  s0_axis_tready_m;
wire [31:0] s0_axis_tdata_m;
wire  s0_axis_tlast_m;
wire  s0_axis_tvalid_m;
wire  s1_axis_tready_m;
wire [31:0] s1_axis_tdata_m;
wire  s1_axis_tlast_m;
wire  s1_axis_tvalid_m;
wire  s2_axis_tready_m;
wire [31:0] s2_axis_tdata_m;
wire  s2_axis_tlast_m;
wire  s2_axis_tvalid_m;

wire ch0_rxprogdivresetdone_m;
wire ch1_rxprogdivresetdone_m;
wire ch2_rxprogdivresetdone_m;
wire ch3_rxprogdivresetdone_m;

wire ch4_rxprogdivresetdone_m;
wire ch5_rxprogdivresetdone_m;
wire ch6_rxprogdivresetdone_m;
wire ch7_rxprogdivresetdone_m;

wire ch8_rxprogdivresetdone_m;
wire ch9_rxprogdivresetdone_m;
wire ch10_rxprogdivresetdone_m;
wire ch11_rxprogdivresetdone_m;

wire ch12_rxprogdivresetdone_m;
wire ch13_rxprogdivresetdone_m;
wire ch14_rxprogdivresetdone_m;
wire ch15_rxprogdivresetdone_m;

wire ch0_txprogdivresetdone_m;
wire ch1_txprogdivresetdone_m;
wire ch2_txprogdivresetdone_m;
wire ch3_txprogdivresetdone_m;

wire ch4_txprogdivresetdone_m;
wire ch5_txprogdivresetdone_m;
wire ch6_txprogdivresetdone_m;
wire ch7_txprogdivresetdone_m;

wire ch8_txprogdivresetdone_m;
wire ch9_txprogdivresetdone_m;
wire ch10_txprogdivresetdone_m;
wire ch11_txprogdivresetdone_m;

wire ch12_txprogdivresetdone_m;
wire ch13_txprogdivresetdone_m;
wire ch14_txprogdivresetdone_m;
wire ch15_txprogdivresetdone_m;

wire  rxmarginreqack_m;
wire [3:0] rxmarginrescmd_m;
wire [1:0] rxmarginreslanenum_m;
wire [7:0] rxmarginrespayld_m;
wire  rxmarginresreq_m;
wire  m0_axis_tready_m;
wire  m1_axis_tready_m;
wire  m2_axis_tready_m;
wire  trigackin0_m;
wire  trigout0_m;
wire  ubinterrupt_m;
wire  ubtxuart_m;
wire rxmarginclk_m;
wire q1_rxmarginclk_m;
wire q2_rxmarginclk_m;
wire q3_rxmarginclk_m;
wire  ch0_mstrxreset_m;
wire  ch0_msttxreset_m;
wire  ch1_mstrxreset_m;
wire  ch1_msttxreset_m;
wire  ch2_mstrxreset_m;
wire  ch2_msttxreset_m;
wire  ch3_mstrxreset_m;
wire  ch3_msttxreset_m;

wire  ch0_mstrxresetdone_m;
wire  ch0_msttxresetdone_m;
wire  ch1_mstrxresetdone_m;
wire  ch1_msttxresetdone_m;
wire  ch2_mstrxresetdone_m;
wire  ch2_msttxresetdone_m;
wire  ch3_mstrxresetdone_m;
wire  ch3_msttxresetdone_m;
wire  pcielinkreachtarget_m;
wire [5:0] pcieltssm_m;
wire  rcalenb_m;
wire  refclk0_clktestsig_m;
wire  refclk1_clktestsig_m;
wire  refclk0_gtrefclkpd_m;
wire  refclk1_gtrefclkpd_m;
wire [3:0] rxmarginreqcmd_m;
wire [1:0] rxmarginreqlanenum_m;
wire [7:0] rxmarginreqpayld_m;
wire  rxmarginreqreq_m;
wire  rxmarginresack_m;
wire [31:0] m0_axis_tdata_m;
wire  m0_axis_tlast_m;
wire  m0_axis_tvalid_m;
wire [31:0] m1_axis_tdata_m;
wire  m1_axis_tlast_m;
wire  m1_axis_tvalid_m;
wire [31:0] m2_axis_tdata_m;
wire  m2_axis_tlast_m;
wire  m2_axis_tvalid_m;
wire  trigackout0_m;
wire  trigin0_m;
wire  ubenable_m;
wire [11:0] ubintr_m;
wire  ubiolmbrst_m;
wire  ubmbrst_m;
wire  ubrxuart_m;
wire refclk0_gtrefclkpdint;

// XPIPE_quad1 Ports
