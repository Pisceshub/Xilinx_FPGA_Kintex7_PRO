`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10144)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9JR+2FTwzOkJ1yLmnse46t3GbkqvKGdMPXCsVU97ufEdNV6W4u47IL58
Jnz8MyoPlqMjtlqhzRXXLit4FW7q1CEeRroKbHBJmfNijs1tjBaOT7URGEqz/N/ORUCJc7b6YDID
flYJi5KZgm+BbtWEB22qHAKg3jeiS3/tmCorTq18iJQU/qRGzgipSfaj81WlLCxy11Gh6P/xg2fd
kMsc6DUZGYAkFl5QMO/k5QdpclmuhozoUuCHALxyfaiA+wTkbX9OgvP7UVlIUlaRSDcNqphtmpUC
j6CIKQblqxhY4jV4pqayCg275DTel/IONGioEd2qw+/ScUjo4Oek+4sM6w76lNRNyEtAAmx7VIjV
wVxgtUmMK+SU5ICtSe1t/04lS+LHCAf2o1H/xsrcLyvzsC2HQrE3np3IEYKSPH+68nBLRzKCYu41
HYqDP2mi+h71TQryIHXHVW3byJwwfRkBtYf075K5dbuJhlQpDFRdgwvEemiNfhRGZDmuMEaulvNS
Szp5zINVsWpNeAvW8R3pAGyrCr2/HvVg+jQ/A38VJ5bLMvpHi6plIqdtcn6ehfwPGhO2+IpbASK0
G8HQoZum7eWDrCD6qN9LSFry5DFSZhbjDhyosOuUxi+DY/HfLRpsq40eQZrqRHYAP7ZoAg1Abr2v
3i3x/AZ45t//RW3viI0lwqwqSOSQ3JLvJiIjMiZZWb1Kuh3crNOCQFOPTAQodCpUMXn76BHyUbwb
0zMLkzd410b7ELSXR3AbH+AZ59yTcDGAPFzYVNTZHGPuqMRTFC7EAWsKwQNNi/E9F4F113zSRRy/
KFfEiMT5+Y4d3moBKJVwoQb+cwWj/b+M0r4x6SQ6GlrIh7uIhg/Y4I83jnQtwUlmM7FOjvkK2oR5
bTOIi0EFovO+O+mR9eLf3mAqoOmBJpfn/d6Ut7k0dB2QHa2I5omv9WO+NwmgRhGsRxG8mBI4vAdQ
dGaupK23soOA5SKmsuA4idg058OXYrE1Zy25zDt2ZnW1cdob5H+pUQmjl41xMqDOXYIqhkfdvxD2
CZDaA20GFkuvMKhJEAkcNa0Td/yXyxbUY3yhizzIntTU02HitZi3Ch4rtgxIbOtVLTpTIDihqDsI
uZqgU+vq2ebdBwGSz4/ZOlqBC6qlhjO8Q2qvIHE8SUDVO15mg8Vus5QCr3FZbJ39kEeqBpsjbOu6
9+9FedS1U70PB/dobq0JsUDTPMM+dSa1rY/MDVhwHY+YoqvD86hpiQVEi7TtPyEtTkf1pDzwamPM
82KYPJWdtb0uFi4gjaU1A4tEi97RrCXVDim9Eie6lwiUljCllR+tvqGJdAGzLb/lOo8siJc/sSKM
6ywZybfkZX616H2wGPRI/+SKLLXwkS0FRdUYj7jC/3wBO5eQEOXZM4eihEjzaSQ+5oiAycvb5c6y
2MTfUhSHTxKJQT+zMQntvAOj8UxZK6Nx4y0anuw1u9IvWtHdb3JKzNlPCZvfx+gjGN+UJFk6oNKT
rahU2qecghGRW/GH9yOax89qeZLq4WWn7LRDZzUF4GR4scYWMAzxQ+ftiYx4iV7rTJ/MoLaZPnQl
98OLNQR4AdgB28m4J2qSgdseultKapBv49CYPkwOnMOlXnLwTMgZW3Qa7/a19MdmD2/7ow7D8kXz
J6GGj+vv4OqgyWsudvS6H8a0QD/Q9gr1nO2g3sPBesx1iFc63RwCPi76IRHfh1w+8c2JteCCjiG4
QaoSj0hce3w00OEef0TPKHm4iK+i1AnmAtpDoMJzMDWgh/GWqsmfv53mEy1UAgDSWC36qpy6AC+1
EtfEZ6KP4nZ7OFAfBBS4FZrMnlYG/SjyaF7r31ZM7akNbJHuFhF69MOslzUDmIvybHr2ZcvH7u06
dvItXujGN/r4f+vuLTuc3a+LbclFk7GMGuP5qocPMA6PbrMYbL1RAVIR2uXKbmhsG2T25ooWJv+P
IY+aF0eY/xpwwakKEKhjVInRebLu9kgCbUncFmgObtsf3aUq35iAGmX+0WYB6MXzFqTkwldgj/Cc
87MnIMAfkf5p2uMrGvTkwdYTJME4YsedaFeJKKNsGF5OEcWgPWyrEGJ8b7vtiYfv94Qb7WWagtvU
Ww9zTCLnwtg8ENObMl3jtjOPoVl6El+utx4r9iSeOcU6k24nCX9nWVwdQdAFkYXjZa7k2ArUkubk
xx1C+6LdE1lbhAk1KSWb/ns8buq0rZkQErUR+npl2IZj3XWhyXR1C7iGCYz2JtDkJzYRFSqEU0a6
A6NXDQqfRtZPsru7HY5lk8YZiDM55vtGH3D8N6f4MkZAwvfV0DhE8+SWmLjsgFdqypegMluuGlYD
l2X3eJQtskGj49Po10/0pzU8ge5qix2KCwjWwbccIHiik0ZjA7t3fZZvaGQh7KMIYiQwcMxl7qje
2hMRYSIG+NyIe+yohqZua2HewzNyZsBGxChq59FvP50UNPLRXznOOLNlKBC89EiK0cO3HUApqU5U
n4PHtzrd61932SWEWh0+M0oAfYTgat64j14qUFlBXsMpMC5/b539z/BgbXUMNHmwBMyLvEg5GW2Q
skAQ7zQYsn2oi6ACZOQCzPWFNGw64JvZ2jOMD1iOwqCzXkn0CERANv7mx7gDxXgkLETgq2E+zgiJ
ju++W+2wkXlrnky31P+9iM+tXcU03ZdgCEdT29V/ZDFWWAs1Sr9HoVolBlsoB+W76yxfF7ZTLfn+
4N+DjrjyKmpt1MzfJ85YkKxVDIKGD7YLcG/K9SHgWN1ZU3pSVxtMf4irXQWKuI82cp403Di+ooT/
MVMi6KYKxxfTPoW0DUgJ7u7uV6LCq6iZprGv7ZWHW7ISVUO+s4G5x+nwLUUKCXMgR3lrr9HkU74j
mmOeJqSROL3vgAetjCJGOAS94QXB/r+Mu7JcycVDSTv+YR28Nat7j9yOMtx3ppPjYPilKYbVvZH2
ZXrgfOCix8+kBRXr0LzOYHxHBegYztjDnmZfU2Q2DMJn/XiURI8KYoWfjn1auPpnzEkAYM+0lvMv
9MXNlfJvKFIkdEz1g90Bn/XXuo0xG0oSlNH8JnpH99yuW6jk0jLrYPXjeCB+3bChmNY6tQpR2HA0
QcOWDkvqk+Mpju8H33JWxIFIbE7mhMYyJYSPIHsFrjOAZhBjkEqpx6oqukcnAuUzGlV9YLLPXrdm
sayyBXt2iLsRTpV8QcTqBfajlZ1MSW7tY+wGOjnqPxmNCu8XahkGH8D+KJumTFmSzpsp/FQLkJis
U0TeA5q8As3UcSKhWknIso58a0qzHoLqbL8PqVbv29HtL+gTBlfYVojIqftBlBb4jeLoIX+cqNlZ
fs1Mjbss8t+OskS6elgfWxQhmoBUOUMuYmlGTgibDkzpaEXNOIoGxnuRN+RNaQ7sy72/yOHC9hoC
6woKsaP536xxMsaaHJfLDJU4peag1wemypC0NXAJWEJ0VbHTxJrdL415nSV9iw/7whQl5b7h/WZY
hGGO3E5rIDe9bfQFjBn9eP8gpMfWrRbzj+uzphAuPK6XAXP1IW3a7saGhJb95PVJDCh7uZkUi+7P
dDTYn7aa/d502IqDvzjpjkV2uNGFqjc0/6n8+UucF9hqHLAIiIRLoHg+NP6bQUO/5qsEyDHKQYz6
2t/gApboQR2FaauDAQm9zoJwdp+5v2p9D8IGPrnDFcl1xPSTYKoRZiR84lBMtSc+Hz14cghCnE3U
MDy5rZlqk703mOTV83WEGBqqb46ZaqTjCWHYoGJiyQL6iByfrJKIiqcQVggld5QJr9goDBAz72VP
jt6uox9hP5fUkSyRgJpRRoxSzNzDcxgMgokw6pIhfgrUOTtberYZ9FUgXSur74oSd66SW1EJGAxC
Bf4LZnFZee/jJ+TK4gRyKKfjJ6f7Q29+yZBF78DDm/TjRqaatU76gIGnpH+HAaTNMryCghNDbNSc
YMlRa8amYWquA2mQ3s6yDFDBZCGRjyQTw/8w27ONLJjXrhJT72DoFO6zJnqo/+lQW24Vpk4dkemI
s5+mz/2LdRjKcXV2HftP31luEs2nRmT7+sRcSOLFODX2wzB3niJeV4E9bLjNMmICzb2LOEMBd7Xi
AQEQaE9vipdrhpsBtI/H+v63hQwp8O3UcVc3/MkFNPX+paXJZzMdoN3vWkyeGlrkuZm/iFddH69b
N7wEjqLR0jrI17RJcDkQj5vwSUu1pLQ2zv5yl7WnZYJvmL6OlB957TtnJnhOQsNtbBZsQbsp+t42
qkUlRzaI4iH2I3zm2LnVeFSVUFKoI3i00ZNXBpUZDho4UGumx6smxGDWavCVZ8LXBNanjLvBZwuQ
k5FsF12DmxuJgbflSW3cdpVX/MaTpDa+9kIXaSTDPSnZufd7CL5+j6+S8t5mFVEr/e6+flhmuwIh
EkA7bj91kaUOIzqdblr/H0VpOpiYh70QZpiDOuSaGCVCs5Gq3v5YC2NHfXqSio8NYI28NZpYvbi9
rLdVJ03qD7wZQW0A9INTpJ4Aj6sGEV1YN+UFdJZMFbcFAa8Yf4H5/MAETMlJLrzOLVTT+ixJvWzJ
Nrtl550iQRRLOxsIhn9pQbzSLp0aHD2EQ7BcTl3JtCV5KOtFOhnBmWXy6C5Pr3X+bkvDDp47HbSy
xtASTmAYnCa2uRP4lLTlQMVsEUJDEXQzetOxIpp9K9GKh/gSctKP4W4IiaL6VJ2qCvkWLQ/LbZl2
4/gPf1VHKsKoFcoQRjh2kVtqJ97rx4j0TtI8bkp8pzUhKs+Xaskaqd7sOPnzruOK77sPH+lmXBgn
jA71tPBYFa9HZVchmqHZcei5DMZLYVyNBxfPF1uUzZl/TEaVvAseYQJMLITvaBbSxc8G8zPtfhYx
6nXgK9gQkOOEAUPLHe2E0kYXWXNiI/B3LdxBMA8AJJfYuUK9br1xsbWA76o41aSvsq+9j6YtJrfs
j5OztAHJ+6t2UUT3ucSq7zC9Q+yJ9PJkk14S5ChPL/JX+d+40LXd2uH4W4/FEy5qupazpyKJpy6R
cb4M43BoV96LUuRorPdIPdlbEHg+LwAnAamsoidtCH4EPTRso7dffoEMYKjkBamdAqttaeNjZ+6V
CBTLrENeWI6I4UJAcGtjbE2KfFl4Z2H2LhkKL4QlKzlC43K+p/D94nuZ11f+JWBak/WO56EtKFNm
m28QBFLuigzlvnVBrgs9cmSc3FdpOcO1cFHBI8xApZAVlOKpqX7Ux0+SO8lRN9sPpOBG71fpWgNr
4f2uAQ1bUHf5kjbLlg+HZD8odsw9iNcugeHrrxSFQqKbL0oGeFyGpz1hDkBAKfJ2VkORCKSN4KNc
ZY1L1reGq0vAwhZVBhskitPC0+5qz63hXdG2qMPyQod34FvWT5piANQQoCexMsGYKgv35KDhYM+w
5qGFg9HiaccK+K2Rp1RmYBPU7py8REaVRZnOvW8XslHVeyflSFjN8PIXB13W9VN5ashSw18Vgbz+
9KnRL2wzKoiTCkKXiOepm6V9ybi6q9PuO9B7KVxWXHl5JaYUUF+CEKb8TMXBsr8rR/Eia8RC7chT
IbwVC0vhazV54mW+E6/5+QTD2zYgNuQYpy0LZeD3NnYCgcBgV4fLesYYYx7nvWyCakf9jJMzDDKC
R8UZEQ1+vLk+Y2j6AcSItxR3XmKJzYEQKDexv1/C6tr8TuqN0H0d9W6xu8ZXr75lPKFKcxKsD/Ap
7NWG3usVAa69QscjdQGKY4jlZQyEXPQPCRA4yYGFkloQ9KKl2+DPJWRCvgp7qiZrC7NHhFw9SEF1
d1LHvqy4u1CLZy7zFWWjl12GME2krE3IO+KC7AXWXIbuILVXE2OHzLrAtDqhgeI/bxCRwQILuWzx
qaBWsd0Ivqt1FJyYhvARcDHefB+cEqBa/FDukDEIxPtXvTdEDj29BGspGOiEP1QVVaqXQO+XGQwD
1Hw+FaNQwDBrwLMjRcCXjAdC8R5yKwYkJq6lMHtfba90/EDQ4biuxfFMgmR1uhZWgdVK4fCG4QpJ
eSNbYqpAKRe6DUJIkF8k0ME+DmyYVBlht+MuRk7AHhQ1OqRw+gZ6Q90ho3YoQPnohX4NUYF8rDtv
KRl8aHJpkCe+Z2GgvpH6p1Yd/bJTnwryXuK2pB22iBK0CMesshqEU4VxvxeKtuDZDlDD34W6ir7i
JH/M04wBkIHbdkCybZ85XfGeXv60MwhSiuxMPAWF6hgFiMa/APy+Ys2+6M/AHXWoqMuhhGKIykId
yiyBHpYGqhXqnmBu2NTyBlBmI6NqX1kXNAVsPpaXSEIbAPC+3t/pLUpNTAuc031yuBYDvAqUHcZV
Z8ce9nRfQQSs1/59uXFosx3fD2Jc8Hf/pbTH9sWmrDmbNMxdhcLO7aRZmRFaqcNhea4yrYxLkGoJ
ZdTv6B5MtCvA6QLATNBOA3nlI6+rqyLVEwTpwwTadtrTtM68Vqepomln9xh8i1iI1bdZOMjJqSbA
QXH38IE3TVA0is1bj6POSat2kvHCaPdKTpm9FyhSp0e0KubHXXag81ko7TDrDdJeFS6NYnz75NNf
utEzJhp9sFdsePyCuUi6ljGJfL7uQP2ZxMhpIA88s4YNrQUqJ4EvSGiZlqWRp0OSCC1cQYP6ZOW3
/olhvDB+dTPu9/k/N3/SWDCutdMbr44edFYAiU1L4tcFijuGECCrr7jGuWn9S5X1MEIEdVj4KLBT
Wqfnbm8t2gbsEEHW0QCRj5nZBuJpw7ymO9TjtMFcyj9Lj1A2IJO8KAc1IAaHb6KaAYSheaQhk5Jf
WoBC0ewMy+SwRiehjRjRUoCozlyZbHK5woNYFk3GRLLyus9ry5J1jDq0B8XgUrvGalyY07nCaxJd
RgkhB2LEYJ9Qr9rbr+KlCPY1RPQFZrzBJKWI06rB/0PjiAvBwCZyseOC7m8RaYQehhjFbrMIJzTz
kesqVxVDEuZGamCdmMSNl0bqEh/0+L3lu7Q1SXO1uqkOy6ZfM9R1c0MNiiqXr0c/LgBHoKkbPCKw
WL+3Yk4rD/SaSs47iRvsBXQaLtozGlRbyZ6OEtRbmFA2ajX/g9s7RLfX+Rj8PoeFvxoju1EfgD76
pGI6N7q0PptycgLYw84R8oOhE5HT4l6tFHdu301BjR/ms+FJlnfBV3zO4Qg9Aqmq2DZZnykNJ2zI
PTkUpeCauS1grUu1cso+ao4LilViupTbAw60szl8OJOcGvyB1zxjl3MUcnulxxnnEkqxdudcI5YH
GlvDnnpazT8bOmwpOuA32fXuLGr0Vy2cWB+rKSM4eV2BGU/LGPin7STR3dOid3n/Ynbbva5e9BVy
/jN7rDiQHN/4J+M/oB6WbwmhInOCJ5AhdJE+wwmprQu4kGqtXF8+SpoKi62hnIPNa5Cal5N9C8zb
XC+ytiBzDRTe9lV7/M9afUzSk3sA3cJ53m0kWH72enpQkhcz25xjnkrm0/3+Tt4UDK41ZB/SAxwq
HrPupyqd0sIU18cHVnRxPW3firi9CXsFNImB4BoLX5r3VVtIhC8KYirY09+ZLmHgwVsEDsVrB/GG
ZV2lBG2pewsJfq1j82Hfz7Wn9cvInFg35c0Rm4a2SRgxvM3yASd4vOqfdrc62vAgIn0jXUF/I/3/
fbnYXq8o5EWhX+c6pbOfwLFs93tllgA9wZfC32SePZ6NGVVngGiJShe79T3y10qJm2TzBGVwZPoA
lC4J/EZQRpd5p3TBk6HFl7vGQUYzw+5HKE7HgdUB5NvNVPbfKXFDqcEaZX6UVVa14DOZDGIyACeF
wQ2rn5fcvgEsR7BE8jyORjE1mOg4+L7q9phyCfUBhHRGqNZwl17AxKScCMeyLbhlqfWXrI3RnN+P
hBnsvnCRYgbGeB0K+/haQ6zs8rwaT2QzuDhBahtbDHhwlSMv533RMHcu2ymuJjYyYN/sYxHMgRv/
WVi9DaHjRA8A+talqtM9uwZzTxmic37NuxigNQ2+iwEnWOWXGfAoe9CoXrSxiNwOJcdsoeGOB2/4
9xnjtWJ4tJKYdshqUxPY/Ni+2xu6dvRKMOcqcCh5gmI2CxqmcYHtz961YZ4J0Fcg2eAuSkn/HP/z
mhPOqrNBbgC2SMnwD784BjawMqPUFF49CtltnkXoLUSves2QDFCM/YI1IuC0uv0x3pTOsIIeBVj3
dzMeAJEELMDpjTgzaTmmONCnbyFNOOwQK5IF+D6S70DubO/l5PFwwbVGtSiKh2/Hy+/NyIqN3qK+
Tpy+NC2ravSQ2KM/rgSy+fAQAVizBQO5i1zyuUIad/sC+pFi5Xsytn0Eb9glLHOkCaHzo3FI8VR3
YdYJ+7tdIIfhDyMnKujydOL3DwezCGpF0qMSg7oz/McocETjYZj+3m38Vl3YQT9/u7APIbdxfBBj
XC7Q4k6F8pDmwKl0oYmlW2Tw54/qCkCvzeDEkoAyTUYLdc5C8mO3eiSHk519MGU+ZIHEh0041TY0
qplZv6c7p6dQz2XRbmz7uk52oS/uVogSfzgCKtgJWlIInjswu+cTaQCstk66mbFuYxSC0E7EGiXX
MOpRUyF1W8NbuuBRV8wzo5YSIBhm7P8COOLQp+O5PxddAteC1o4xegO+fq8r+6d/cOA29vcQFXgZ
VT64KQNvAhz9soH22gaZHtKpQrqtsNnHocF6hx478q/8wnHwu79Kl4HN3ETe/K1KD6FzhaLkCShF
E62+WTYjdc5veOx4+z90pPaQsGkm90xGnFftAJhQAKC9p+xtHiZqODJVn84K3IqO5yWHOuz+k1/L
Nok7NKCEBeBvF0cIqwkQqoCkyD9RHH7kDUm8429OPrJktbxrqyWoC8OrPe/5al7QlIRZMGdxMm/R
t3+4LxQHZJIFWgUvAgIhrGwAFfNpwx76WR3i1ud4A3OvMiJORM7ZIulV0HNFL5hLIdO+IIXwYBNJ
3OHmkXrvKZnLrUAO8DxghhU03eyCDz/JfDE7r32o3Dp0q9PWADgD92NpBrEf+JmvgfsyY8eO959N
4bO0qK6LN3fFXTnaw5L6agLgRnfkEfSNR/5XQWkACBOsTcpI1C4nsqOtp4EqN2qU0VfNLiHWIJ9x
PZ5R1RtvXu0NmRV2SE4eyfHghgMDoOco9JBkd/HqYGGUw1EC7j4I1jH6gSAFNB9ZH38sB1JdZPTL
lLpQ5y9z6rkYM+x1M3QXLeNLAs/eZssnpiWxwBU89EUo8+hL8PTJOeyCUDiBTqDrc9wegCzQvZap
/o7xFnMhFa1pmDA0pMEEzKGBkoEb2fjNNPc6mEYM1BHkTqxpKdJA2X//SBAjeC48o02wFwBVBgy5
G/6Eipf6S44PG6EacS3Yj5Xibkuq8RPQTF9eoyHrA6VtfhO0Jmx39ieT3RThEKewD0OZXeiBHXtU
eKmA4sAouMNIofD7RwxoGclFMWCa6xLkrGE5TfeOB4Ptu4brqF+2o2GUnh3q5rwgyf8K5DU5xUz9
mZsK7HU74vlnVeNxipbVzFbu7T6wnlDTAOz7wL6GzJUvtCPahC9On+2Hy2LhrzEULbTByeMKtJMj
u99delFOYhR1+II9ZCEbc7FT+RHJMqzYmJppBKC7hMmOGy0rJNKnWZYg+J5RXWrMGKQ3LnluHqdm
pe7c16eCz2WTdC5ACuGDTEJfZGbZW90jMUr2hN83TIrCFuCxndAF13MMXOMWonWHkNypBns8BP4d
6+OKAu7d6U5AzodWQuP/2S1+yOnuDM3/lhDa4pk40spmFXTzxKzQt+nhYX9J+zQWcGNtbR/Lpve4
r5Lcny58UD12XF0A2LEImejr9gE3fH1yP1NnsGy9PfgiSJgeK+5K5kRjxg7dEA48MAT9mYPZk/Yt
scuy09TsC6xALOwVhJkHHfV/9/ZV82sEqmTOUdlOqSjDwx3oXcRgW9V+bNaitUM+ltv48Dmb7vgF
YZbdU9Aj5jGoN5A0sKDzGgJ3TZsaH1xkp6r4tUb09568kkJ0VbOxT+pGlUZbjEZ2BQ88xhOZxnrl
x1MxHiVwxg8wsnFBx5IAgpkQKskPuo8Lo4/rW2ztRVURPhJSRFStgKT4ViwbUangMNoqCK1CoYss
dElcyD+eBrlpADs7rZMprLJpvc2yP5oXlQt7MkniW1hhwzHIiviRRRrnvHDzdeM5kZZUaK44IlxU
06PAN6InR6t5/Nns1MBxX0jM3je9Z4luhbUZnQvUla2DMe9y1aAVzYlb+UuRJvD/1B03oU+dsaVX
VFgxXH5xWpWL3nRIwOyKHxwONERlrQM0nhVLd4eVd597PFQ6GBmE56A0iGcWMue2TFk26LDntHJs
jRmIKSlIwkZ0pAurC7cbwc8pj5rgIKDphRJzEpQDC4+iWm8++zTKqibAXqjUoX5lozW3aty8WEgh
qFetuPiLLN5NEIuSWgPx9k6UfUpvjg2Cy4HhyUtCTYNJnD1zQ437t0GznKh0lhpI4LU+R/nbYrPX
1OcQEXAgzUajvqWLXj4YGkL1loHAZR//spUJu7tqV9XVfJdIPZKA/edG0d3Yul10mILPVCshnEQ4
zqp0tdIQAAIVZMDlpHwEls5/CLTvDLYG9pRFQQpaq1OciF3BGOTPhmeygud+hg20n7aHeMvgdAOf
FrXH4oy4j+KzfHBeFrbQzJOZE9ed2NTV3keAfiR5Lgo0hRHBnrmsjJxP9og5vv18YAW2KuwgpoQT
3pD+tNR37Zd00o0YAqhF04RKCHFU50YMjFzbfTkQq8rsZERttxliWGBEa2N5yV85Q34eEb0So15o
SwUZbialt50IYpMyC71Vww/ulRzG4R+HlIoV0dBTIi9UUJhAHMLDsnVhF+hm8iKigyidykuhORsY
a0usifJWqKfn86TIGY8nNAywqEaghoBywZrbOGOXRyKTQC5jmZeK2NXGvbpC8FmGJqXEWxpy+dCb
1xDwt9JmUUiarKERYlRYNQh0iNrOTwVUke+ohfJAvbrZX+xHDeP3HtZOToAQn0mTdzS1tb4+IFAn
4fVFJuL3sEm2ckHih/lv3l1LjCHwIq4PkVN33qxEWv/eM8OW90WxLQ6QeNCe3saNuFCSdWj+hUJ7
A7YnK15Ji3mYWikT1AuyggMparfhTEqAmIRxybZYbopXZnRoKrldFOrZ03mQNGLqXMOXRCC1SaUF
pAxNwNt4daxW3bFZzWk0BmbDYh67S+6bbJcyPpTUN9IM3cM9PIZkmBWc85N0lwKe5T/0VpLT+jt8
GRL+lco39R21UmAWw2mvS5nRqzgbw/Pt92IarVvfipK01uOpeaZsxK6LhpGWxIFSZkbSccswwTTK
cf+NvsJRiMGZM3uhIAw+HLUXCWFz8+yoDgmVcNQoKosVThlYIRomVs+J6qn9uEibpk1lMipbIkhZ
TsXiSmr975g+HMnJCWJ6vk26MU3nlMK8Yvp9HvBJNiojaXVgbredYe8gI6n3UrG1AuU/KTEreIEn
/6omCln0alAg09Uh02FLj5+B34G+SCilbR4Gr8GSicCgdhTW3J6WeXgRIR7vHQUW4Ju+ksxwrap8
MCraYzebYZ9vzZviaxnH6JZ4H7CIT3Nyo5YTAWKWnkEdmXNMi1dbmmQz9Mi7DoQc5yL3U4p1yJgD
i9imCzwdin91Xf3bal8iBRXN/IBYDtXxsrh6EU216DCllBdQLSi84aMCpcQZoAnvRzsmYPE10w3E
2lXF0ayJ+ek3ibFxsb76GuSLcl7wuKanN6vSN3/UaNbAo36hgY4VpmgZaiXGFSkG6GXLjVKUKWrd
Bp0p/5rRUX8XsidT3aDQICp9peFr1tYPjDdNgCkbWa23zOVzf4n96Uo9nRckVoyKEQ6FJcAvfQBI
ukk/WV6zJRvDzFpXgC6dKs9fnKTJJkr408zbH41li8W+ry3s4CfhVMdR+m/MJue4YPdmLgZojR1X
h19TemyFy8bytJ8h+Vk1pArw/BkHnBM1mI1Dq5Dphr6rGXMSOof9J/BjRfQmLbEJRoVOh9977mqY
+yGYOqx+XauTlpnZcFEeOuoL7aSzLrEPYLqayV5mjpaQz14AUEF200jDJhVbhLTQQVu6az7DieeD
Ush3n0Vudo1200GfRMpoPdcWRb06iOjp1hYyOojINeMTUNOL0p6qD3g93qgn4LHiSZ1oFrZAkho6
2wMab/S6VmNQnbJtdKC3MoB0gEBNxini5INOqn9nQBasx88bwuQFoYAQTE3htaPJ4sma7+cz1rdQ
hQO9JiRkwvrX8FsEspT+SApT6QxMuQdyRPByh655HO+Cs0Scj+bgelDTnOn+y//RPjbdRN3zEE6R
VioPTdhXuBfDKJwnAt6diPkNp5xGy8YB3tKwakW5el8ruhbPfGATiD5vE+MCfcGoR1cJZQTdLxhy
au9W9LuEr7cZIPL5Y/nCW27OjiGOTL1s3NrFNJ5vS1fhsMZQ+E1UHS3O/AmW0rnmMDQ/uLbv8F4y
JlIHifcoePcPs/TH5uMvoKld8y1udTOczxXMGJL+iSpE+S+pvSvDn3h8Q6T0dFmdkL26rSGBU9Tx
udjFgWm6EKiMfQ8DXplgMzKklbesc7C3AoBBpK0l/kCAzIEPRGKzZpyCCcADFz5VmexowA161nQ+
WtD4bLjFtbzJkNLBwhYmrVZiX+bQKz/G/DqjMuCpyF+TgYXDtDyXNbFWZCQCfu0Cf/TSONASr7Df
kP58QFFld04oYjLcF0Zl+ciZNzLYFGrrMbgW/FOjsI34Kck38ETIJVxRh+cowqN/9i4qmwYkpnNl
Kno0RwaR+ox24RyTJaUxkbwWk4W6h23CCInEREo9yyuSUhD+eLCjximScUx18rHxCf118EG9l6A0
MVsKUgd7ot2jiIr7+iaYJZYQUXhwqT0tffl+DbQtAr+9XGxjN99H+taMRjzndp/xiMztSd0ONc+f
1/6WCShMVGNjCwsxSugKsAjtAs/utDC7Fz+l7sTNy2skVh64bY8Kl8iiG1XAs232319gn9m7hdC6
nj6oRtGuOsgpt7xcvlj0L8w4swDRI2cKks3h5BG5KJgSnsfRqtx34vRbS2AWN5DjgRuw4h1SFg4S
7+5YyPVDbQbl28uxrGE832IxUttnlBBLieiCmsuHCeqpY/xMrTt9XUVXgbRpQaBFod9v8odsGlin
vR3EdB2pGDZHC1klfN+1ih2RdNVyFcQ9H/LMIDr2nB4CTjjajH9yGBTs73DlxAZjxcqlz0trnnmj
TGsLcZ3ESoj/uSpezI/brxVdhpdFEo8d4mBX19Nir6HD/xd7W7rhTQ2Eypdhxv57x5YFJREQ7xOR
0Hp06mJy5thTOHemY7gDFfTypMlxTBLizOQepHRRk8Pfj/XvbSVRapSKIstc1+WG1bAXlum/h9pE
a9VIfAGzgZgM7PwyXyOSXU4OPif5fNyLH9cemk1Wf4kwCfI8uc/DX8RDAnkdi05TN0ihlo2wefon
tKRwdxAiCYz6fKMhQawmH+qqFaNK7YLENygtNUDvtveARZ2hp7/KohIoW57fbqz/q+t+2stAny8u
+i3okE3no0NqjYhA628ENylaTF5de+o87Z+YLd6hQhYvaOL0ohMRYkGlabwrJ4KmUDiLD1EESw==
`pragma protect end_protected
