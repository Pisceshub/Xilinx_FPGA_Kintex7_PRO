`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 236256)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qFdQXdrBXCEFYEODs1Ipl3tqV+sPb7w4kumP5iXLb+GW0BqEsbHb+HDQ
GQ3aAQ+Gy4AmebE3mo1FGTeiDXcw6pvETTaKnt7zAgRyQtEJyTBauCOi+YCBxzRB8DyjhQrGFtNG
2uLZI9/AMCvrlgGL2pSUBLFGLRJOUW1uWeWWl9e5VTI2hQdNw5uLeVvWtvDbCKDiy+S3hkkMxC52
5OTgC7XgQd0vlhx+jXzaImh7ZNB95U5nUVNR/lvX47YRCYiddYJGXQnPrK5/VFA5nwfJ4aLipx2l
5W/iW7pBkMNdJIWO2ODrP2x9HqgkLoAwnok4ypOSbaVRhTE7N+tFooV9ni+5ShE28fFXdv2Wp4IS
dzRrrHs9Zmd9ionCFKvvBtrX5QmwnYafpLmA0NHLDdaXUy50RzO6+/BDEIqtdTrg0OY39Dv6wwsJ
X84I8mk58uwO11Pkyw+yJ1zXO5NE8drOYss+ZMHZVCaFwEOO6jB/XcrmhNR2OxzXgE3kO58lo7am
ufjRmoISZ0vpP2RUm8/BP6f0/dbRe8tVhKOWvT+pMhbQ0lpNw27jI59TgpTJrXP27KpGmFVigZ9C
XZKLaKzEnWUqp15DSQaRe7tQBpBUWPrpSU9icPpdXovzpMzq+UPv6eKvvNeRhqxHhRrn+C0ciAHT
elEcslOD7+VV9B8yVEHrSuor30YG9hpDH3Vr9FGVbp6X3xlCQNbDkb2dJ/0Yoe9AHmmByN+ii6qL
6doLcMOoDh1FHaJzWsG0BNfWWjiDTNLz5ud1l4D61ZrRcru08AW6vpVpFmrSH1ufGzIpzInzVWsw
e/9qwa7K2bK/GJewOlFIELgg4F2I4nJCJzCsVt3zANmvT+W3C/3vdpd+Wuwf+ESLE9MC5ndGxePi
6sos3qzV3WsoSlZIMWaEePrHIwjVOX6VeS4CAjqJvbEQ79p/X4FTkj867EcL0cH0QTvANo2r4ia1
NtvWIHwYqslXiHJrS9q+uREXV0g3ySff1nLACnHJhTfCrQAGeuaXG5JyIDmqwpiIqamZroiYWye1
RuQrFQUS+7D1h5wzOjXlq8+tY42bbDBdWDP16x6GrhxukBXCTHUEZTbAuxJxmFREfxMLdcs2tbNR
XAGIwk13yMncSuBAvVsFz6/+4BP+tIsav1d2iBgu8GQadcM5F+jHKEOFZdnXAY4XTJ5zhPdS+50O
dK76ZR7rKWkCSdvso7l6I2fEZ8vjHK7NV0x39KXcyhsXWSGRZ1G17kIpKXdFj/JmN+pXuUfEJcYd
+v7HwIIASN3cGWX/PETro3RuTO5Md1WUF49Yxo769S+uz5B6KBZ/RTTGwe8xt7eEVCAPBkZvx535
KH8bgydvgGDn4P7nNOa7ixaQhctan2vO+GVCpLrnjqVTuYcbnjkUMn9MW3lf+wS3KRpljEX/aW49
XZjuSnypwLpLvnC29P3jYpLOVpRL/aiVlW0OHY7eTyfMWUTvljdrWX7v4uJwzMvTzAPFil0474q+
Nh9zm/peGA2GSReAt3SOyWKPRRS6IZnVAzAcNBCrWkN3EVAtSBt0YAYd5DLgxNe/2yKXfyQ0Zd8z
LQDWhRqommGyAPy+jNlqh0XBm7ld/WsjGwjbd2GpP7n3F9GdhYn1eFA+EmPWYbzcLcGZet7WmXdT
CtwAWDTUjT05LUb9YVQEZ2ZaiUcmibEietFQMOH0oAUJT8ZRVdkdJrw1564FixBPpeDecn/ASlkr
Kp2inAXqMtvg6bCTFbSKlLJXG0oiKMX8KXRIXxE9xdUqNNryGGnswn4ukyuhH3r/3OimBOIbBUu6
TtGTXZPvAUQc79jwi4428qjrfe6r2XtFCgPMmddLLWLQX1HuTSiTZmDe1fkzUDF306pqo8shVJKN
+TbtTiQJWbItM/Fq1BiNRsEkHGT8mSsG5JNDLeXMJppqY/geHASX5bMbk9wf38uAPoFFkp3zeu9p
39kJTyo0N4uwoxHkkWz0ek7G3vLvcNHEw3silKgF7dfwm1+evzWq4BsVi3B+wrnebh9XCZnF9hU1
EbkYnoCNwLTA/9UAPJM+tgSe7H7ew8LW7hu1pXYNHAbZQxf1xJh40O6vHQNboyfEI2i+LWvilIva
u5sracdOHUACNhBqn1fdRpcTC8eo4w2nk46HreiGKbcqZ81kB4gDpF6CSp1wh0Phs28/6cRReIpH
5/pEtwxbs8Oh/+X2TNPIKSEV5pJTGu1rYn2OYlijdxVIqPHAaotgjGPzo8lIhwizIevWZbFhUVPy
6cBfaT3Za9mVJrSgMRZQw6BLIqX4UL2wAWHlRyMLcvj/5wN4X0gLD/aUGMounIbwmnrEhCoLHTRy
hyHgr5gic9ZdXi8UmmQo268g9BxJwThUqFftyDJ1DznyGIyNBz/0cuXl0bnVMIGZ/vtrhiVh6XzV
3SbEVIGqrh4kiFvWtYNwsQ0hQiRILv9MKkNPQ/bMcQo+vjeaSrbdxNwBatFDI/zPP5bNsbhBFbDH
Z5k2qUXfZzDwzPEBBBvXUcwIdG6Mny69KS6MK8DhGltGzywXuHG84hFQa31H9KfROlciTqkARkfj
ZW72sHzRN8q7vGGexNoH6sZtb/3vxYWgjLuyEOPAfT0INCgK1Befllj1kWcTBroirZG/8if8n282
Al3IH1rXAnynvrqAmzy3p4WhWRKpRFxHzGKT4/AgQU9gyVRnCpJDY6Lw4Pc9lKtKFbzb6Hnw53C6
N0Qoquyy6r8MOPbKppXuDVXkqsKXOg8vv2snYJozmjTWwM0v3GK9jjIOWtaeYWkeCH81TtIUadPV
HLY0E7DE4KlQ9J+DwpLsL8MjaZG/oOWtS2xt9WiKLP1lB1l7AwQr5UTUI5ULyVvg3QeWuN1L69Uz
Z8uNySTwBld2Y83mfj6RzCMhhKpptLM2j00vaR108yu3hXn9ml3EoOM/E1OGq2ojoVhdd7+Ldc1j
iawH8rsGH7fJakxErTANNc85tTtmERTwuzkzbrliDQfzla/7lGcwOXbjmoiJN31G29vcg3sGIw4l
Awk11j+WZqpP4nOoubSVa803C/In124BUxoOamia0OnzsV8HLkG0dnUzA2B9a8lH0nYZbIS7k4WS
Cu8PMTaGEOaX6yOdDM3dnhORAaIuKG9JtzZTzgDTNPxoLlM0yHJ7pZtZkDzr8UV3FzZxzBtTdUKN
tfvofivGL/yO2h+YtU8LZMVI5NkJ+tS2aIT67JJeeuIxgRmGD99jA6BuEenPnuXMKpXCQD0WMbZz
KXIM0tyCA6z0s+c+NtmzDr3r4DkX8CvUTkXjmyn+v+22XftqGlpb/FJaVoQtTW1AMLAWU+Nb27fc
Xq/Bi+yI9sYsEWT20qndHZhQtcUZcSmCqU2Huldis2jbyv+1xvOVZK0K/XjWV3lWDqeCWMtnQAEU
iiKYvb1o6fOIt0K6tafLmS0Sz413RB5zHLKc43OWhZ6oeDjs1TArK+/+L+F58U8LV6jGwmHUlByw
6RRok0IrIzBEuIbdQvsaKKQAZo5myhQauUlPEXZFvuWdWkoDyey071LgFSuN8SxMWqYyMfEnxDOt
e7iU7lyd4vdypUnmVL8rSkD5Qe2q6RnIb29ndXExzkBWWDSW5TGbfIZK25ttU09Qe0lC7x445lZv
vLqC7SBjG6DY1RlrZ4j0y10dvNVr1LaMRHPRdgP1/ho/qOm6Jqcf0/kKoMK7FW9dBbwXHNWumG4a
DXO1W5VIywCIkNCbfNjvKWsXJiLL5mzWmXSIdFtJlXZREUXn9y5rIV06vkeqBCNe5K3zf5RU/i9K
EFdQ2nsqK7JGwf6/semG56XEZCNd/lcxVnmkxot5im9LaIfa2ddF1SKXkHzP3Mp1kj/jlVvBNB9W
NFBDVrIdnuC99aCJDux99bYnDU8+HtSOWFv/5GeOweCHElgc7fb0G+/7WMgjn4MXDrfPN5Hk7IS7
Qco6DIO9s1iGbFaM3c0Yo5f4I2PBcC7JHAlAYyaUwefhWZruO6fK/28rBLxJOijDXX1Q5MZ74PAz
5u0X4DkozfvMxDpLo3sbG7by8T7Zf11i/mkGdfTC7CajaU46kGhhyOxaMhp/D5k0INXcos0uRUQl
EDcnaRCUsxekmDak69TxhUq7ktL6Nqn/6TxfcxwXyvtsxB2ugFIjN8aB7E+eRh0W+U6nYo/cyREB
+A2LHvc6xcFEDyk/DmvriREXAY5KKVeMYKTvEOXz+IwJJBdMjp4iD4Q3q+nsN7kg4ATMV8sVYrLB
wPvg9fnyDFFSOfkZJPggDrHi4CBX/mBGHFewkFrKev7imCNmzfZOhkDZnpwWVuLJlhYWY251nSnJ
0MuOtct3zpB1mYdDLGUW8m0rExOQt/leE3e1MIx5VpfSbfPCyXz4kg6PHubsB/0cDuZ1jLinNP+g
nj+HTftbgpc/Fkw/PiO71x8fTUDZ5Z1qTSHI9heQKH7Gy2SLmqfp+YV2YOurI3oT/ZvZYluyUJ2p
O3AmSLN21AgsElExTMgLIKcRKnStXbX5azPVqD74Ligg0PlimkhDn3582kArl9p1UsLEWXXiRImF
AE+Bs8D81BCqGwTR/s2W94qzAZY8Ayo4MET6LW1gfKEoePTW6uyhMHYrZqobMxlnn2ZdtxlP+oXU
MbEz9/Ha3Qm1QPwvskjxlImbYmFFVYICAjffAMPf2H/MV3tw5jZx1Oqfnmindtr9p/xWRfQmyoOh
MgF/2ERPqD0k6dGyXTnA4CeC3NmpTZFqIsbbGVAwaCS76MaIb2MC6tysN0MS5XZUurTRyvFrcxyX
ID1T7dQr1JhEOMxPcqTA1mpjQJTl6b7tAPNh6oUswZYkQeV6mNzmgcQyvmSTfZqAdkTXOcLgbdVz
iEDfAH/2HQfhHmsqvsQ6IL1HtLjCKVOyRagBsermyIaBzstopfwyqOpRybi8qCo6deh7ELZy49FT
XAycrYKbnipJzngym4D2O3Vfwf9vxSBBodXn6qzYI7Imwa8K+tAUHKNJLcY/5Rwb1mttpUS7+AEc
wpOYgH4woyMH82PdxKPUrcLNsORcXt2IEJ4HxRisT5nMIfqEf0IIdJcGjjmorIfJWXEU4krJH8Jv
B9D2+81K9LmBshXmTKuioAciPkf6FJGBlUpNt5n1tExVoKkvOh6HDXSTrVgPPnDL7CoOomBpMt4L
MZABsGuuqSwZK1jRioxMyYbvpnegqisRdxOmfSFpTc+pF2Qa7W+yrW52L+8miBV7WBUDyTX3wQym
oPMftmBaQXOiZ/GcCH+Z9IvRAGdKUejudo1IycyMBnzusBxK9bjiG5emmkzaS7138BuRoosELMls
P2+clWbhLlw2rpcyHjrgC7DfTYWJAQZ7k8JLjBSAnLMKQ91T3/FkmSz9RoQkg3WKNCSqRxh5wte1
Sg8cPFtcy41t+ig6Uu6Z06RzPFcD9y/+ExDlICf0zRBJy4998ITIFgTSaMetr/0UW7zpkkWwyMum
XSKxOC9ql7wqrrEQpMx1bCsoEqMSxKPTRu5wVKKF9swVVF+MUgczMBywMIlT+7r+cEmCX0pzWJgL
fUwucj18xbig69xK6SsTpbG7Q629/h+lc2ZM3Sk/v9Izufd239IaWG0ev5/x4xo7NeyBhQAcVJ+F
s6G90k+DaBpXT3CxZmZZsD2eR1C7vp1Xxsc3lDRi+9cXOOoihDi+VAk7sXeLCG23LCOhlVGkqn+X
D/MJoxkCi9LRzAepKt4AeI8HdvWMAgfAH9NQe/78JxxHbFdHG0//6Ike03s/HNP1J9IRvxOMhzT+
XWWHCRE89Om6JgMFNJYU/oduM7F+NYs8GibFOQ/AgJWdLGF8xvry3zINoquZ6yNkIGul85YcoDbD
P9PFq/ZM1LRcHr2Kc/jvxnwLLVyIemn/mo24zzF1t2c2xRjH0DDJOeUCQxjd38MScnWMM4D0J42s
/MFiaKxgjRWMq2fbDpnT+yZYWQ6MLzOxYHBC6FTfuNBVl6kP1yiERqPzwnuArBOynjNbuIqJ9sl+
5+PykqGa3663oYK+hBu92bwURIuCtXKWzNUnAcXO90PdMemW0hVmf+3bB4mBAcj2YEc+f6VU1bgE
DXrisX5gxdqR5bUK4dkOBRn+QSA7qYj42SCuoEkZBLIjUyUkmb4BqGt2pUra5hMu5h4ORM4QVF0A
LpT/dV22WhZobCd4cSmON6/ARzL4CDWpJDdycfpEy0NaFnJsd7hbw6xeqXNX3sc15GLF+mgHt43k
ls2x/05lWbdJ3XV/iNXfvDM61w4wRy3ldHZYjsQ7oGLH0Z4VHSe3otQP5b4fs4Z8rbksSi6eq176
E3auThsA6NF/MTMSm667DyuxaS2bpzT3BSZMpHIrLHIAFLX50Ji6eQnHYyAlVM3Jf9pUfQtYtWLJ
tMbQ8WcC1ptyEFN3orYsVEpAo/hVgNwYJSj2LvpEWuYeXPysXroCISyyRNdPgG3DC3uBESeEjqVp
+MmfKrTo0d0ZC+jW+9uOIdcogBRh9VbA5gzPcMAH86tPFYOGdUwZU9yCzRY0g3g68ZwMCDWFleml
TwX+s4gZaDhcztgIsXe8BUz/e1mWIIrp6Zg+OAXJzE/TQcR7ZmkOmK5bruNmbEEXNBgp57E5q2lb
ZT+2kn0TWbH1DSBnZr9wA/RUpgyNATAQIk1UCsmgyQF+XDa1Njv1+jN9VujUi7nvdC/G+075pfIZ
G+WDHTv+6BmSD4urHtv0ObVgq6bNuieCy9YcPKc+3fmOL5ttiSk7CxCONJi0O8CcEFLTq3IJ/8wb
Jm4egKVZik5Z4yEN6V2u3l50TFwdlA86ruENvUftlxLrCKveweIloyJVCHS+wsNnLGR4inIZ97CI
fkb6vN8lYxMFRsq0TmdbLe9LzKUmEDR5F+HteEw4jH7OSFvcYBzYv2l5oasUsqWGkmu56SRFXCHs
9dLyli82BJsiD4ZZJ/Q3967UR1MI+zbToRAlx6xyXoxqOXs1logOXJSsuFIvzEalht6wZXebIrq3
gjvMxN91t1TUSEcy470ebOSJbCd4oQ/xLZxlRpIuAqxdyNV6CIbPRxiKnoTMjaFCw2tHuHlOFyfW
rWFsJNb4dFl3XPm9QdBc1HFDM48NFOHuyZKP3WTr87Y+sgr14rCVjFwz64u6rb3LTpy1oK6RM1hV
dKpwdjMMYfMpTLwGkpEBoLMOdxeldL9DxTyUaCT6aH4CFAHOAys3BaeUnk2XGtbsj76DG1GgIw/2
1ZuyP7DWW+nMvFkRyu3ZKfvOVZKuXCK+M6UtV0JhkksbmMDUAY49IhUi1CmoZ4pZ3+0sGkPT2NOj
Y2rqN35WudWlpyGA/6YDpQsEhcJgDB39CJMMaj5mZh/jJVN4wwjguNL1KBOaj29VwKaiaYQ+DM+C
BFwv1arNvSfyhzRkft2/KyW/AE1+++/cts9YCtq7CEUX9dS0B4af3mmCFu9vGdE6Dy4B179KSeYy
No0DmCqZyiEhjvch62yukoJrum0csapewxdDdgvAyH6U6HiTGV5to3CJhB3DJWeX4ic4YbGbKiCd
3Mt3ZF8+e6w0acp4T3uEDDJJCl2Y4yL1hL/HSgc8I6B1vlhjO45f8ci053eMMPeDDTCAgUe2kyEF
NqGfjs+br1IuuLdRKoXzfMe03Dd578GKoa6vmckvG8B0uhjC1vYZFXmptMh9lfkzVtjcsjo9I7xd
7+ycnDoEvxXOsNF5u6q0Q0LTQfalY9BbSM1yuuieZ+lDjaCgHgLIdd/Wv8uBUjICsywC0Idq4cwO
8SxLbAm8YBu7AaqcmToXz+KZbGtQYcWzp8EWKTvPkzcl6pPWy97yvg1EiZI5jiZUCKYY/+P9M8V+
pAOnzZ0xAHjJteN80+qYbnQ4ah3pa+UvpVUxYztGwme9ywI4x8AmSBQ18qpiwMemhP5yNgCTL260
CS8YicniZ/VSJxXGolVOssqCKuA/8YvNm9bHDR/WDAGTkPz0yQF8g40fYQ0yG1ySonYUtqy1Me73
gA3C7xbURxUp9eOKhsp+nJhO6O6ZW2+NdhmG3eqxVDn0tBeN3FRdz5dobc9tmV/pQPdr8VzFoPGf
GrfxthDPRfrN34W9uclu+duEQBowVGDgVG3ij7gkdVcDfFVwm0poSta6SCnT44hwp3NPj+rp9+7b
vCxCRMuGbZFctX+bD/PttKO4Zpqy0/k2YKOXXkRU/tFJqMb/DeF+qKN2chZh9fOgD24bZIfv/1PC
Vr6kgcTTgvxEPbfwCEPduSVSKUPQJ1lJljMSsUQfX2UbNf6bfuV3flHTSjacRXWWczwvsXtywRGw
ECYbbECtvCJ8YtV0AtsNVvAFjSQzycwqvzA1V8AH/s3W8btdR9oCnW47avQ1Yjhjjwc2EkZMqaUS
Y7nt9qSJDkvtUDI4hmZQ7KhMwdyMYZ2kFpfG9I/9YvVXFhfJN1VXdr0BhHKyNw+W1e/DUybsa85x
YSEE6BmulcV6hr+JGAvXVbmpajtOYEXP3CPHv+STeMdFJkM+UcVzTRDO00AkvPQ43npRUdaHEazp
y3VhXP4+PfPQlpKPC6e8GpquszC7XFcS58OXMK3qCEeDBGJWDWzqAmZSP2GVcaIBiqmbLR5p1WnP
1AgrNcdEo+k2sMawwU13l+NFbPfu2FE2aRh+jmI2SPnFzZLOHuawLB0F9rWEZUzaR4a/jl26bTrR
0xULW9nm2dcw/6cWQvABrC4FDFEdDlbpeh8aawSMBSQkzakAwsd9XpxhuRzgh30Ayvq6oHk4+jxd
ayvMXYGXknv3+G50W344+rnWQe7hwd95w5D//R++3oTLkXXQeaLycmlf2HpA1YyHlIH2KuDJPurj
VzLfqTh1Wbea3Ez7OloPHAod1HNnKLlV6VGFrB7c154/FgMD4OJcIc53viOBTMkZRNXgZVskNC1s
HXknObIVT/9f2tHDS8HIqCYTWibcFgYaGNUArTEkHX78nS2Y8+70Kb9x3tYojhmYae83hrco5YoG
dty23bd0h9F0oZMSX7rUr/sMpOr/aPktjdr85CIXRhRTq17NyAKWTB2SQaNVHuRMrj0HUwIzoEPv
Q3g6FnxDIspYGeTWsVoWN4ivdp9L2s6ZxGCw1gAkFYKQlsgWZssSMfUyixxhKs4SQmNpA6qbKbF0
g8ANIjk/EYA5VO5u2kW1B6PIYGxG13ms2mota6+KyJhzuLQGBrFRIibkNH6iywJQLjQAQiRDv2Gl
y0uDlh8YMrpPX0gJkAznC3kT1nNrUlnH8Mgagi3UXsNS0z6/gpqXrrLLlOBxYFnpj1wkaS9mz4R0
8cVjuvQc58k3d9YbiM37ST5HoiDzunUcdo6iM88QSbEXQyklGkG6qwv98yOM4KtxEZjp5pPdnpW0
p4zFz2uRstBN8mfazVAQmNfhFp0d/ItmYcYxiVP5L/9GwT5icBFc20LgtZHzxx3dnPHjY/Kdc4Qq
KCDs0A5JspZDam+gv9+ARtL6d4QmfL/e1B6xPLpTG3bxj0nFhsq2BDQ8Zk/+Sz+XkxzVzP/2mG79
VmNnxvJ4S/7eq3In+p4ViRRwOE7H9wvbNgHEt8HkP3EfzYK8HN6bwYJYqpEMrVtXHJJF1ksJRcz0
10xtTuOPkZAQ/7A/Jv81/I2QBc6H+tssx3i23PCXESdZNzyBu0K5foBJ+RSQ7KAAHkwjKkfflQ6S
uagQ1GrWuzP67nP6fU7r2sIOLfxVTlM6iDeomB+PRl00FkF+oCj6aXO+g/OO1/oYRQI0e9wPhlRE
YYWSBI1G39EAUaJfZKWNPbhwgHXnla+vxpNHY3yr7rbd9yDhgVh0iWb0OG9wxF4ToL0BkU5dOVzf
6XNjHCGUX7H2mUw3T0a088FKMkXRV5Y/ooMTWRQe/cisxle82wBAPEl8/ftmdDsyUwP566uxCEXz
tQyrhXnzo0oCbTaUdhIt1/LOFedBozlia/+rL7nnSZ8ofIz6l6/+fKCIUGYtuCruYEtB1vQ4W5Zk
MrvH+pqLKpAhh0PYjwNThgi/vp8eT4NnJSH3OovdXqGW6qFYdHxuY4SEGgMGgkBWvEpeW5pafydN
6BOuhf92CNKFt9l50taR2dAiHEkDLeecvfQJ4pHKTv0P6wj8UMWJRzDucyynm1efqWN/od/4SU6L
QRJADCUECV1+953ftBCJOB/5ZqPLT01KCkc55dmuLNNb+0qM4nbbXvIyqqKkFxm/g4Wuhz5yYOYo
VwnBCKng+9ZYBtocgoCVWhI7eFPaeJzKiZk/+CHj14xsCy1fADHdcHpny7ZYY5E+Ie7s/XT63r89
fp7bSaGo5ehYQApCJ7AaZGQpWEEa4yyX35p7tWhFAcHZiQl0zy/8QKGCMBjifyh0sCb1i4ZWjFsL
h9EfM7ScxufbxiamwDCtdN9bMo1l2YHjSlSor7ZfwTdjaO960GrA3dl/2Nl/tyPpbYQuDEyVePY9
l8MNrV2DkyGBDmYwV5oLlWEZnOz04Jt7nmclZqOz8nllrpH+eVvKdnrHEPJWsiH6jKMNt3Btr7+y
oLkN2gU0sGuNJDCVd2uDyW/0Zu9O6PoS1EbVyk9SCEj2eqNdi6GHKSKASIcfKmeIiqA2IUfzEgdo
Y3LBCoSyI+3jzEgdveCt83MZp/7PpALAbMzsdNQsp1HEi914YWDb2s3INlQGc/V6PiFXPDhdGHhY
QF1hE1+ZRkKg7U0FS91H6gtyGu06MqOcsTHXhO0Le+PYUXdZntnN9FuE4FsxyawCwvBkWQZ+gcMY
gxijXKNtcccu35JdlTjbg/1iyg8gq6QkEemh1bPynj8FWUozhBWp4HTkNOWnSh3MCl8kzQKRsD4+
E+Ak6JGQNz4+QE8rLtxnovI3y6uoUvapYCI7j9PLZOIfF1IbrqaGAM7fTHp/NnVGOnY4BPBLQ0Uf
bzhsFY9alO4vtJkzDIlWQdGKzVapV0tk2d5/iAe8DkiRPKMfkFKjLDlGyCOnTVvDZJG9ORkvmO43
TfuSWK/QcY2y4ca4/rTVs3DaepgZvQpuuCMcwm2dI6mAZ32pDWiHG3WUHFfpYj1fiRT032dCFVda
qO8Tx5HvmLk54gux77OlHXBk7u8TUHFP5+qFGfuw4A/RjJzsRZqo9TweZA/M2XYaahaF/4d+01qH
Jr5n0ap/etXJQKowMX8mGpFHiE8SZGCFHRK2KCsx2YMtHKSIlomXtN+WqD9CnKBA8YRL6+zZ6TX2
wkRLFRX0nN28RJ1Z46QFX/y0I7vFB5vdwy8AGoxaAflfEztLEL1NiyQqUX5ZVAW3x28itSSGOVHN
fCES9VWJEXLghm0OCcumeKuON/MmDhA9mvXbPaRpcWGnnLCrMSV/ZpkdIGAGzjVwK2cWWowhTa+F
AdAMTIMV1kD6t9uw5FJCJSEF9yDaiqGrgC1pvcYto5ylkxfAjM8LIjhEq3fiHkiS/IifqPqs+ecy
ihcBsvsRH9DItuF4Tl8/63EkHoRQ+WAfag6lZuxnrfJwYTyZIP3Jy+8CswXc+Y8N7uGzSSQyn7sb
U2Bf3kT/kEGYyBjthCP4b/E3ksDDcASStf9nBKc9MpNtI8eA9W9x2mIR4zrbPy0lJgg4cMYplUMY
wb4ZSrfgeujYsfGxBIFZSL0u6pEs8DGn8JpbfroJP7kbcUOLiw0ELeUN/DHFpyMAbMFptlB/1hIh
0NjrUG8eKiz+puQPwzvoa9QbSnaly02+DSOl8X09It14W0JHB9hiszCyVBOBIjjCBI1MEHALZtk7
6OB8P0J6xUJUtnbUUS6+XExEAbGYArlF6sZWk3RpOiJ7iUzX3E6G+V1MNVRv8cDlIdoWO3vBkTSQ
Qm2MdHvqWdPvtJYE+RVL4OOW/op1oLhE0QWJp6HO+8J4F2OrY+JvuZgamxqC6FhDim+4XWK5vJ6J
R/HD3P47Tao3+AOxK3xnNV2a1KkN/SPvFFw+1MKYhyBI45sOlI5RNsUQ1YCKPlFZRlGmuehdEBNG
0tNhMvxbcJaOSqm6t05WP8UHOq3xpOeMV1UI9OebkhR0yQXWVOzljoz+C8Bgvnkgsfc7WvUlZtLM
cRASQu0AJCCcBzIJ+lKWI5hKys3+3Yah009SRZ6ZHUs2k9MlUJ/HKsjosTKrWYjHryY4bGl07AHY
XvUYQhC2ateekiuvoIo3HiyByxjz0ZjNwfFgSAIYLOuW+kURHSTS6NMz2LpowEdpakXvCCACOUFJ
66nrw3uJyOu2WcnFieE+0aYmYl0ssQpHpWXxJqC55vk7sRVNEAVoxRZsTEZa8BvBbJRtYtrexKuE
h7//peWPm45WGi+9Gdvw4e6a10BCd5uNX6LkMV50tSPtPMQRqG6Un2dyodvDgfIjW5VZOwIZ7v+Q
voIWsFvK88NYyG+965NtGAR/pVlPFXRqIZ+/YjI8oynivkWJyMSeZLEv4gjadxMvQMLi3Kel1dCC
LXFijDB1eVTXYqez5MiE0b24w7oo/PD1j/DL9SHfFKJXx/FO/5sooxdhu1YXn6Jgmq3UWqlOuiF5
XgAMn+2mPg4KowUpQwvhuMOr9J5qMVWdoeV8q1cD7MegMHMYwH8sSpS9WsAz6NY23pJugT0wtzfF
t/DI8Pq1BElw/7BpkM6QRLaO01+220i1xpQJBKILQMKZ+EQ0dNADvBluh9H4g4TGmnfSvrN0o2dQ
wmREyDpHq/ShUS5EZ+bL2vnsbRdCcqW7zc8NW4CBl2E2LmpFOdYTAaqoCiwedzMsXJsQdY9nSzA5
GtYhFGEdKmOQcn5fw5ay7tNsp1xtFJ1Ul299DHYlUjmnIzRwdDi1+B/h0UYZdiUbvVk0baf3jV1j
vz906cN5FE+GNPP7wCd9KGlR9pbwztoXbzjRlq2sRhEk7CveJX8O+TVFagIHbg1+trEJkkkh6fW4
WCmItfLnVR2Erpvz5eS/ryukW/EcwlTODmcnGpYvlIL6LEenn/sZjVay5NbigCfQEDHxb/TWZWNH
eloHTvBrJsdc5ROAFl0LXZEWfYOIikj7Oz4YybJ/DLiTixwnHkotZ18jKxquUGqab5OldduNGhe4
CzDV88yNtw/4CbBVxsYVflpCbWSG9v4WMt6wVuUrwJfceTymuyegxk7MMa32O2QJP5b+QHCJP1p8
H7a5ljjR/qg68kGwUPOQP/jM7cXkWOHzD2K1BxOdgifA7n2mgANwCdvKwx4gRTGUe9w1yn9Wya6Q
knDHesdzxXTXKYuEdUeFwo7+kKsKdji9Or3ESm407uTSZ3ewyJZL3wdOfZ0dwezPVyxeAl4NqdWH
JNekJpxVTK1nNdjpuIFEfseUZDYwbuG5vW/18yQR7IMmI5j5cQ8q6o3NdoxX8ppOmxy9I8/pObbS
gr9IdvQjk7Q+Uecl7wQlpNzn2MLpHy4A1HrYcxwjC7j409YY8kUmiUiDWGi735ZxM20NDSxIfuNz
wU8JeasiEgQtz+yos+F3OwdfqaNoc5In8OJyOtp6rdAg0pSmtIHON0GnmXhrCaZHndjI0fYaUht/
1kRVHeRb+91fGHNmZMAqZm2XAiaK6cohjS1/6WEur01Oe/xNtxDY4VxSFlU3HcuuV0Uma7+MCcH+
Atefdq0EkPes2+5Hm1ec4BsAQosEyyXNcSNJ0rt35rXquEDjQysIH6rTsuHaDKkIJY6XEXlkx0KL
iTjWEV+yyaB49guPQ+oH8qhW5ufnDNx9ODPx3Z/rD64LFfAYgP+qMKOZu7iMmbiWMpYo/m2WAOwl
MXeAVqQzs+xJq3ZOo5GBAKwFx42wG4NczkPRvrlQsRHMY6tTk0g60rJX57SYnwHYfZizEkZ2eiDu
73Hhan1bl0C0rmJB8CzGdzAtOm4c767irAOT8J3f43TRQMyg8Z4B7Iua2wMpK6u1bo2egb6ewE08
7jtFPY5RE6b8E+0VYdr89SxthcueSwGhdUDtDJZvfK1+MDJ4mmEvaARDFqmr9o3EV5N3mqlkU2mj
hBuvDsXnhKDRix7Mf4JTOF2NqYgFExUnoQXTIBeUpsC3CH5ASyHB7DxU1pS4awRMC/96eiWYkTg5
zzm5TXT9xxJRMCM56btGM3qMs00vlhWWn7zdfTGekKt+8TWk18CDL9PNvMJuuylqrGMqLtcUtlxe
p2X8XBwuYAdQtogZoZM8DVniU6QNJucZGaNnrA59WxlPYU7GUt8zfI7oV73IRYg+6wPQ7AodlvJY
l3iuwEg9aV/ckYfp/OLGMQslPNrQcwNz0b+PBsZhOeKL2mOghGPO0JSB+1woWXuJAlmEMEaNrbAy
o0+00IWjrF9JoZwmLCOZn6SGPW5CoylqUIlUDIXv+xPfDWKvuMUmbkzJ7LZLmPxmErdqS753HT04
8/vHm0D8Oo5Na9hPWx9VrQISBeov4L5Pqp7gngPDJ7R+Phy2kwPj12BQDsHOYxLPO5SP0GDpf8gH
dwjr1U/7Pytc49d4xIC0DGvxHcAR5IjGXidF4wDH0GDIQ4WuyFtJufVnDEtzKBMbweGIF0zqxegA
uF1g2Vzf0JPV/EPdttmFrNRUsPc2CzQ/gCp9IRSBbet9xHPkQGw/x3uj7zeUb3YQBUqXl0TxXZ0d
+NMfz6Dw3qZuo9kj8uamE3dqJWB33Bcy6w63RC6WEwkJO2GOg1hRNltagpWcJaGMYf29aZuv99Tk
+TSsbQdc4br5oovBrSiaYrwIS1F61QE1Yeab2Tau/bOOFJ1wOzaTCJRjOZDDaOBZIqEfbkacpNVz
MMnSAQRzFNPk9QyVwq5ArI6s516m8UXW9uU4ODKOAaxtqcS2lqxz91lqXc4rCBG4T6cVUIY1s7Bt
ZEE2TL7y2LVkjWHB1fADZLQLk44/yamgQUxhZYrn83KDOuAN/Ayya/CdDhgb1rXFKl8kTNMYoYkY
rPNst55rACof4h99cytK+Zhyc37eBQHZbJ8FrkcCN8KxDhRwcLEpB4vxhIL8vwsKlxc95pfcUYP5
GQ7pAGLsy9tH6Vibd0yKrNMgK9ChbVGCnC5q5ldvaaNcJ1aAyZEof9xhxBTjrp5HZIKtpqn6DFqF
cSB0TXFbFssADpZ+ccA9UEHlvvL82koyaiKOGGHw5dk/+BLoJVfdBPT9bmgVETiZAr4YhgMRstSP
8z8oLSq3yV+4p55+MTNkJBCoPGbZx1yT5hcQQ8xkmwvdcZZIOcekDsSg+J69+w2g0r5NhBsi3v4J
iLCOVG8GdM+TWOzDdIjD7bfIgt8YhL/v0syvpUR7ZbvyAER3BTZut6BYiFpiL5XNz/chTT17lDrD
cL/6LNo7JhZh/kfioItFzrwDCn5tED3nq1cKbNoXiRkW6hvtTrMi2o7xo4WXEygzZxxphiSArnuM
ELrOIF918pxtbwbOt7TNIKbanuBgp/CkG0HUQtyjpMRIUWTYddFinRFZuKu2pX9/FtBcEqScVRna
nKC/Ez1E7HaWcdJzaIqCHH/RVhcK803U8jwI3axkatyc3eBtY92dXe3VnKBcGFAXkaQKbcO0bJgg
xdoXeCtbsOhbTW/3GNwn1Le7yx/HDqaIcGYV/NE6uMwrapp329lG4pdiQ344Kz9nJknD+pGbWuLh
f0nq9vx0l33/oqzgjonCBsXJduotegvWsg1fT73IR4TLadrkzkp+GdsCNlEKyxkiMILZtng0LfuC
ZWCHSAhSk1PXlv9G0uNkm8g5QL6OWcqyZoHjQfAZbadgEZ//719cywKmAzadef5IDMJzQwgPpOW0
SiDsQ18vaw+kE3qSQgz9WqqMqVVbpCuH8SwTBGkh/ImVfGI5nfTOUkppe5k5D/4gcyleSYbVdKcF
BmkNpaPdq0E6UOovSw2dn0oeSxzAiEJwB7LPoqpJpaIZ9qBBHx63dJ8V8HbD+GJSFyT2VSg2Dpkc
qiXRkRqn8mpY/fdeIxZrOy5qVr8PLiOCwgqG5sPYlT500CxjS0K0ykopEIAx5fZwhDZCwGggxuMH
2sg04dqMAltpHzfTLwJYNg2BCiblxSTBv69BaGcuCmMIh2nX6YW9QStKcj5Oau4Ic3J+2tZT8zbi
FDIhQ+pTvYaP5rwJpobW6O/8iRZiEEqeBk0HI3aXsA2tMCRR4Mng5qbZKyt0CAkGgU9tEnjnMvfj
FqyM6ASUGxCpAkpmDGnLQGXAXESDgUnIi9cnPv7Us08DpfUOIbHZEyA3YcgOsUsEcB02a7ImSs6N
430ofHD6Y1qaT8jb3Gb4LteYDMxcHO7RB2w8EucPeC0douxPyj/lq9eckP8Sy8AeAukWJItJoMIL
Czo6ncj0ojokf4JwGCAPsMtZb+wC6cnF7DGLsuPo1v61R3UUDkl4rAS4LPSuXpEc4tcldOgQVucd
XF4K8PQQ/rNaZfeVebNVs0UM1RMzQvX/HMKi+wn52hlKeYqSs9fB0ccKD8FxJS5y4t1sltG98sXn
MO7BgFhCHioyUZOhfhqfEDn5HfvTGm6g4Iaa37KuCH+in7cxMND3jB9EBqzsIACWp0/fVsGoNXko
VOqT/B3nhgyuBxTDqj6Dq4q3paPpDH9tBFtgdzrT0w5DUA0RO1y3GF8SHVCH8QdBRdmBeZpcs+OA
rNQTmwKE91qt8Qmtjs+ZHh7JJONXEE65t2KhS8erl1YPuYgW2/OsDiQ5d6qUYjsyIIa8XRFVZ5rd
swdMxwj3kR3JHUmWRGwv2OHuL9iJEQzV+TNoLkRiHM0kzWLL/DThIi3f+o+VFzKAX6TCNnDjYyj2
3H+ohA8XqxjHmweZJt3PNx87jvJR0UOk57dkn4FyGPCcunN5UW7OPIkKE7RyuqsV9mj8A1kGmGvo
g2AMlvS9q+Sqvt3wPhoKx3tBOM2NbFTGyNgNQbIAq3mobU974UsULDXtvu0mhoR5hwMNPwBzSlPY
zyqtwwbsaQ5ol2+oWztH8KrVxa6kaxMJSeHuY38tnqKosJrezpRNibo4KazEZD3559b3J7r946Rj
DbXiETI3EGDjLOlQRP6AoMjvYqyO613wOqPcydbAjlqoBApmTymapTl3ky9pldpnB4PA3zS7NI2c
+KK/doNjMz3WiEuHgVMEsG4LyAiKsdBOQyAdFGoVSxqOGgPASbB2rkEOfxorLqVmOOE30qlxoozb
tLkAhFaLnkD2CSlMU4/v0rgvpt9FIg8J2PcZGu/LygLk+US+YtGbrjChcErOXdD05FTii964b/8z
VBt8AIYv63DDlcTJcm+K4Z70AmGQm+fESL13PCqZ90mEAn7NuyPG+PqxXTISyfnXmQflDckyYG9v
+e1LHIIIAlWq2pibXCiCytFNVbeDkLJFn6x8SfBvj1FZ6e36uet8oAO/bocYhc7t2IMit3hrjGV3
5ht/C7KH+J0+DANNwWZsF51ssGvyiQUUwgx/GQZksqUu5Oz1YOKZnn4E7tTV3Hq0bmRoub5dGjg+
9kDU6VYih5XS2U0lXYGAOpdUBjB+LwDKVEDHkdmJEHh8mToKGf49IBDQISGTOC6PIw/Xsd7W2Ln4
SP0HaohzHDz/oXgkmD66jKygirVFWre8YbcqN0CBDek1Run/FCtKcNJNsl+2+FxyixB6NdYwB5bH
qO54pdkwecCjuVWmOJcjohXusYirlJXdzqVXVQqhD5m5bExH+MNJb716i+LA+SRG/YleoFe5Vm6O
M280zev6rQDw8r0KqWErvPxbUhldgZWwaOFMZBBEPAoKexrrRqLOHdAQvZQ+kdljuz67E9MwByrq
5ljbgRkV1f+wzTcbO4UCayvugy/tE40+LhDhbalk7D5ulhIc5TmD3pgIgwHhXTfw47abHERY5JZm
wPn0cqSXNpHig/NUHzHVYI7ZSWFnsnLRpDChODJYhhcgdFQotFvZ5CKze03eDh32CI+wEPSI2J6c
XwzQDqOfg2ur/yX8tObIaDotSxLgne93QokeCFFq9qiuwoyqaLVWTQlhakA/jMPku6hDGmRz10t9
cfenSKm3bqrML5AVuTj1ilZarH8w8QxpeTNXR3jh9Kw2sBXqc7RVBCtYvk0Yr1FODr66OuFsmATq
/i9ekJjtciP6j2kT0Wz3N9qyF+q+rAhT2m+cyCvNevgZeRckn4DtsYXIqxTfFpTO6pXp33+GgPhF
aHPuo2PwVPEU4mHENvoIUiHPlVJPzSrEC6oCzxmw46NxmiO23R7uIK1kWE9x8NkfzPHHflaitfjW
JzE0Wv+SvM90FnUJ5wajizCNCeGTgxwq1cZqms7YF5PUB/fxXf0Bs+cdqGra2y8QoUVU6Hae9vG/
0Y6pBzMSo8i0aEWH3ipp6leK9p2UXzcw9Jfm4XQpR0Whi65QYnRc+LVZjDDfL4XwTtPNJbm1usjc
WgUhPwr+34Wv4TWN1x3UWmMjDjhl/KJsn3DPRCDVtmgbJ3W+8prDm/x4s4q8QQMv1Bw1+TVrgvDJ
BgZQH54kujn1eXcjRuAv5l42uxwg1eVFq9Hvcroo93hdmK/yTcUbtP7jda1eYBq+QIN1SodjFvo9
eV4kvPpzI09O49qgHDOpHVyEolhm3F7rkP8CxxmOr97lB/qwQj2R0ugGxmLAPA1C06vUYjjXmtDc
HqZx23rpQNxPKeHJi2t1/RAXnuWWJ33MhJTkCCE7k9goU6XOO4FKgBgiBo7rBf47aYM2MIDOzHQv
07MZtkaumu0fPUQN/uq37pO/H7mn+wt5Et90bKikik79pjLDTr1dKYwL6tpmr3o9u+KdC5mILRTn
QeQfHVrE3OTRBsHB/k2ppUz4Ar8zeiC8u3+8pQMeDBBD/M19dsQEKoj1xZgvrG5f5V8P1C2pX4en
2T273rPC/R/AH6NhnxmQGj66stsc7rA2fuLKqLRn1Hv//EvU1EhMLW624tRrV3yfZHWePYRcCF4u
sE15e/bIOc7CDqHiWQYTvL1zEKv02Kfe64IZdhYrYAX+XGh08T1Ea6inhfyDZsUdoCWx3O5NQ6VM
9MEV4iWbNLP24NW6paw0nm1XRbO0lVJJzMCvS6v2aFMQZXUYjgbDz8aDAYHu+79gYeHSq4caCpHK
dbMWy+cKypa+rvZ03nfKPyjQl70JvMfPFwq/xHuMdXON8Vy6LUkSOT0ojMXKYiSwFRv+xlL8KAME
sdnHrZ6tsznQPeSi3jWQRwm55vqvh1sSu3JmizIpd5IVikg2HsSL9gtqc0qMPdk9rC+fKlM7pSVq
cAgyN7N4EuXRoyao7p2rzgUAZUcDmVPhoJ6Wll6v7gKDf3iZMg05l4aoTl5Efhg4HA9CKd+1bo8x
C6ejKJiIOY9DWSQd9BsI/oy+YoVfHDXaYBeupTnvHyaQQRErczv5h4MPp50z+rrWYjTKJQ9U5Zg0
VILPsM7MNOARO2R6WSv6Nv4KsLUjYdFN6kWh4iQN8VxkMqQ4oXr94nIg2e7edf2AYk8a1yo8PYD/
rgUGAhLX6ouGSWB7HhpIy8HtnQe+cBkcpwMVCmPg4zY94IATptRbzApUuLJ1v5geJTp8zccvwyqe
e6zEq0vvkgz0sSBRkn9I2H8Dp3CV4l5OVl0jFaYQz7aCLKrfZg+mMrQH677u+jvxONh353xDrtfh
VPZ3IGynoTCzq6d9vz7NQv5bP7w+zP7dovZjC9WRCdzCcbzLcwlMGFk2nwl6b8kkfYPnoYSuoJfa
A4GOoWx0F8xvzWdzqEK0Pj2xeCXm6RFahr1+sN7MD00CxmKBO7stAo+jUM0wCVEcJ3n9fCGgPZ9U
7ejYCS1uVv/3YKVapZUXWzIzn4hsQGYjRF2q2PNMAkhcAX7pOt2I26cQjrW0cBlvWcW7vBnd7iSn
oWBa0tFvtL4LmA0uzV1/4RZFlZVGsjefXkN/TvhxLnkRPwxAORb8SrTb4jJnf89Y1SWDKrTaX09i
t/dqTbKpFl46aKC6EkGvqJvLGMikMYoGzDmS3IOm9e2pq/sSLfQ/s8sBPSgOGKa8PLShkqPjjQol
o2oKoXoSivPvj8mmwM57/5ljvpGAWuZBGe+KW7zPs9bTRXgA6mMlM+U3HZDFbcRjVFhbI80Dw2lH
TQeKqIYP1kgxU/GOdJSl4ll0krV30UnxrNuDZRGYHBRgpjW6XeEWaQl8iumVhj2UHUU8gh317Kli
FIwKJaPtZgkUpUr6rc0T+7BXXq4KlKsew6aRUmHXMSnIFk3cK8e/+3n9xlQKpq6VdZq20B5p2Ejt
UPZ+2QW8SUSaUGvnXGN/5Am3Tkt2BQf45okc3Pdx+vW5YDu0yRRCMlTm3UymrXbwh/tU38YVejBB
X8Y7icJbHg5vkwDaw0Y8JdMibyH2l4PUWO93dKjsw/ftw2SUJeyDBM9gJGGRkSxs+8UJH1NPPmZM
Py95GM37yBnbKnxzLETyMlAByI1uTvSLWZL7FWx+hvGH+F8Gaf0ztARY7Ao+z4hDh98ZWGn9MCY2
vhPrf6SCT+xKdFqJ5cK1yEEBYvXmkRiNeBBuipYsXq9ohj56cWCs0Uz6qFbHmiU4nBiHDmQF4xVc
ch9DW5tyza6aKex5cHrHpiFQsc/+PgwYOK0XwuOQGyYj9VW5w5nYDY1utzfC3L0yMJ5gwbJZFmqR
7k+3eEY7gJtV5wKXkuqqSGacA3X1XSd1TlEXsx3SxvggfYpWaYZDhknoX6Hgn4cYOOi0X68oNmEj
4Q5VKydyfMEWr8vY3xxN3xjZYt5fCKWFO/PeLwTB4iP+Wd498h3523NcjZk1+in+TSEm1vca9Vi3
do3sCiRoQKKFR0Cs6CNrMExPpox3+nwztojQLD8cJWEK+mZPTi3ksGblATKgcuc3ak8W38o7k01p
kz1Plyc7QwUt4TYtmtfCsmgF/Sj3i+xacHBzWDF2a0xwuQ7P5c9dV9qaQ5FmRozM9clKCjvwJtoV
V4DKexhU1gl+9EWrcuvHDyMgnDVCRIr1M7aJGcIBGzIJ2sIs+lCahT3xoeURnzPRkVDhAD/qkCpt
Wcjv1RiB7mrL0x2Oi8/8ynszSzkWRGivVPrcl5AQ+J8sZGDSvEfww1mj28YRq2DotI1S1wYtM12S
SZM8kU/4D4zZ871fXGc0CLz+GFCCWAUi0E/8NqO6DzPtPIH2ATXU14ScZHYrS7j4MajjXi6uABbR
37be/vwt8kFZgKNgceuk3uNqKbYOlWBtesJVdRw46E0M9LaGjhZ/S5RlpvKJq00oNFAuEXqfY+Gu
B4PebvfE+UWLGlnH/y4DSZglc/RCzkr5M0nyItUET8zu9kmPUVzpsnVaxyhlvG8nf6TucUfChEmm
ZF+9TVH4PZOpdaqKSOow8/GBrzjYnb+NDVJqkK1vDXUEa3mvbTWCuf1tblCXin39tfxWhp68xyGB
S+lV24no5/Ic0/1VyOh27WCgBrLrQwjsd2j+10lqnhPCFyt2KTHff1T2Nbxor7Ft+l4VUVSEPIdz
N6KtDlOWNLA/jTKNWjgzwnPfSQvba1lZ27jgdavhE/RIsZixwbiZK1Kp7NM6oYRVg3rs2RcIGVp1
njOYOVTDvl5YciTVk/oQsUDKZM0Iht52lknP2asWtKKW8FxPlbppl/fDPqSd5JM1D8Vy2zRC8nmD
Vk4HEETkwzvoKZU87L2e1D/YiTG3Gc4CoLbvHFofNOHrNlgKZhwnsbu6Wle0BUQ29K79GLTG4MWX
ASrBHoK8X/M9vL9rsjTDrnvt2f2PUajYMt7K6i3ygPlPjTRZH9v3dkUE82xOXjjTn/Ogu2foyLZe
5tsif/W7xYcjdaPyRRkwWQx3TryU1fWrn0sMtyPcJLtfWpKIAGNtFrIy0dZJtUxsQcWuEMI+61Q9
mF0RfbJdxslda9TnCW/Bkmn8HF2QEkEeIAFKDXkkR8+r8Qlxw9y1yHNgre7+aVWZ64uRPZeaJcNh
JL4S6u6uLRWPByNnD1Fb7nEW1Qp/AcDc2pb6z9LAzNmfx8k4brmo6uIg8oCtFTgjuFc0CthXnK4X
wOnskps77Wq7xTx0WQD1ED82GkEz8oWGk76L37jIgqPHJ0W3poxa0OqPe/Y1niQYQlidYZXzphjk
3CMLyOOuTpPAyLYgOaQkfqkb66Is4ICu29md2NkIVd9wk4HIMnJVlU0NFOA8PEfOyGp+ej8OqDN5
AuUlKHVsLf8nSkoMMO0I6szkfqgAdaiyswKKzrNyFDuSsYHdzLTZXOI9tYs2YwCvf3Jw18QWKRTx
uQUe7ZwUdVZKYsCat+ih8MCv9i6TKKDY2EeUPhAt7jVmKQXNGtUvnEcOVgwGhqINERYjCEnTsxk4
hS5Gg9Ucvov6qOjQb0UxuMmv4LGfEy6Z7iDQHqGNsMRuqFDHNoKH7ia5gEQbNSX4Qq+BepjBsdK8
maCuy842SpjvRf7BQMqTBsGMGRm3Zqh1buMOlrSc2lHumpD4zTFzAuE8YaFvWq9VDUDZOxZ15Ed8
NaT+VIB1zLXztb4q/L4OZhOEyP8gpId0ZfDCQg5L4D1hzQKiNpND143Otwuq7TWs8Y4KF94D4r/N
tHwGb8BQJcPGKf8O/dDlsgXUAEtMO8v6qPMaZM9I8kfpuH82BVarbE8WUZ7paHhWJyvxL+8eNeI0
7fNzfSUzENxevfHI6WPGZil9vRIgwdrc52fRoOynaxaREudJiiOCfaVJ4MbEJEIxFJ0Z5wPUnGGy
W8ni3ap2+2vvTFQe5FygPkWiH5P79AnshbTsj5pOEiiDSC574ekCxE/RAowCyuCfiuR6WHLkJRL8
nHHeO0tBcv/aOK7d0dZ1MxMXvfIRjNbu131xKC7aWvmcNaqAcxV5crW/kOQrxfLtyRwiBUNNePy2
a7RIm8xND8+/B5Tk8HNG16VFpgO9V5l+AIoG1O7F9qQzPyJqZ95b12fp7X8OIdLh6a6mpX5DN/m/
o4uU4M8NmqSB/0MUmB1BQIm857bE0PP6HtIBlTNJXvskiEkfTXav+DyS1NxVnq2UDmQRX1ItMUc5
SiGKIYqcaqSDCvV72JtMjoV8ubbxpl1ssYqn9Sl4Bq67sgDvEK6EgtpXwc5kT7vyf4jXhS09tBI3
b5WLwkl7+uPrWDiTLzF5DPs62QGMffO0vZrEMzCKtiJ5APWiBKAuFCirv6oC5RuvHhyBKZHJqK2c
P2KPpiFsOgo8m5g+SgSoCT9qiDYPhYq/sbGqGMJcL4qXUOmjSDnX2Q48tTz1TaxUs7CapRwzz5+5
gWvUcNWvTQzLAT9Pcyj/HCRpv/lfm+VzPOU9Vf6IG0mie/48+ZTttby0h1ASUG3FX+znzmfdPeA1
aZPehUAMPYkGYKiVEv+xtEnLFSJNWzcGEr+Y5WS2apWFojTN29Swuw9MMpxZrOnIEY/Y7gGX35PD
iz3mBhlJaXKU6Yyz5sBVRHQupPfvOmVEXxewzgBL+KmWPit3USWnKViE7r3t9WLA5p/YBupUVMmX
A+McvwgMaT1O4cUnup210JlIha93cA4p2X+ZK1p81RRWXuedFCel1o1yrgzfZtUvDIMwsBzwq1Mj
Wp5BMaM71yyGDed5LPJlyNxY7PqYU9olcAm1C/3sJvmrkZyxuzHhRIfaCsoB50W+y0zwbv5ynJc3
k5EvAq7iwVRfXxCx5WtVTnyGBPGtoVxGALNe5RlMxlSrhholohOlhkqr43Uso7yZ+YweKw2/thkZ
Gwh6PQvREiFJ7CYYOJ5L0mqJPANRHG1PVaW0uQ+3+9LSkkcpwXnMFYrIwds8gvmO2lNaXh8L1TPP
/UcAV/r/tOUZ3WIQHTzS0PD58QagPM05rkTQnfXtlsjiJBEGPSiI8yY17t7g/OGoWP2H23zIoKRb
CbGrM//eejlvArS3XkYhYG2H0n54PtRhML2UV2Ec7pKzoU3o21ZgRHWiDQC6WkJsEa5ASSS5MM6N
LaL0Xd39Zk2O49FLm3M2kUdDfUaj6gRKINNXtw22MafFQQORSl5v48MfyxnzDzolsfL/+Gdj+DIz
kywTqNNNNg7Xr55HxkKSpX3g63f0V9yeIL9y/Hd/qGvVMJASxeOFORiUpmL7eTKit5kpYVMDrYC2
6DGmm7ZLpegx3uOgf8Gtwb+2WkpbcVtMMJGJt3KcHxV6p9Sjgf3agBy6Ukf5KAVlA1hNlmP/xFmt
/b0bnVVsIWNEOCWQjhEHGefyXaupiZhsikEUedO4RBphHZZJOYxIe2Ynfj0AkB7/g7Ia4EyHxok4
o0gXoSaeL8KSmByb42DeOgLP5XmR7wwhX52Bjj8ZV4+mQHWD0stwpgVzfrYk4hzmPNY8QDRxSKlw
zWAbYBLbnF30nS3OgDbTHbbnyuNGIk2Jwel71mYHToQGWxbeCWf0TEjPi4/zP+dhPuXR1dhCnHL7
EWdkRNvXZwnR+TOV1Xo4HyuxcJo1kFM4VkXYdl+wIe/0IIVenGUupa/65Y5aIliwBStRpNIGOtFG
UR83uoNyZ6/B8SuHGmJiTuU/ZIaEyErbo+XJ4FFEQeeQaB+WzT9OEmmnTQv0UmLzQu5TjKlySmNK
ghS6qY3+APBGxz70dZ8uo2Gp3phcHAWuUvBIhQGla/alqvngrxh2p4PVplpO43G/acMdTuyljovx
/fJBNxFU+4jxrPA6X3z3RsJdTCnYZQxhTM63MGFMVe83+v42yHpYWyz+xpLMbc1xU4dCsjHkOJxi
6mwEInyr1fIlnLD9Usw0BBjGxzSujLURw2qzHTDAaB4ukbzqnJ8sqEMDOs/j10JjXniNd9K5ZrGF
rTW5fDWM6gNPdpSk24E8kFfJRYug5Kpg3VJIyz8ydMMHkgEJPvlo4hb0JSvxg5JUWdPOvCz0w0rb
3XlnJb4Y1jquwwTx6pesdI9CzwMvEAB9Bks618xR1I6Vi/VRi/K01zx3txbO/bPbaGPMaqIJtELL
ESZmAkM19ZC9B8Lgzfut40e+84NCrVfm+gmn+3bVh1g33fL2+7xA0rUNbAS/ADmfzRJXIuXEDaVR
uxPXExoCdpIkBlqzR/rNX5TJMpSa+kqkc2cG1/B4nmXi4s4US1gX/ToIeBbPFLTIV45yJV60dk1z
WPRd9X0UEkcm2xhppjRk9/N8j5Oz4x/0drjbUfLjdfSE3m1h23T6Xba3bqrc+gwbybMXXyRIepWt
SsYMAsuTNarmnwFww9q1G7W0YZN6EMvQq3FlntYtVPv0Fr8aklZmuRA5+FIl5K7s1uzyHKD+nZuM
96A2qrqlZnJZo8Qd8QWtsnk3TA57tH9zmNE0nH/ce80eYjRquqMVAOM4xmeswbVEG952LyWHSJ16
hG2BM97tnGkmO6qNq+f2qUJK9UB3jbEiQUO4jfYjbd0zzdI3kfi8Y60dG9QCO+J7wy4EjDGnrxnr
NKgODGy/JPsRec7ke8wVEioh8vZ1SinW6oqiY5zw4O0X+808Zzq5Djh3rFR8rpiM4lp5eoKSSMvF
8Qzum5Z7NCWgYJfqTCls1ZbdpDxiSPJWWarRUHf12cosg3q5TX4kXj7PTXAT6C1jnylkBIkkPFPF
L1J00CmjdOFba+F+SRRauDlefsxPQaonfb/f7oqAzxqLBhW/I32w4tcrVp9pDcWWr873Tp1Ge5hK
yc/G9BUCLeUsdEs6ItCaxb1WNuEl7cHczEgpG627jneOXZAoGdfRPOg8rZGQKINlzm+gQGpTTmzv
r29UNhwjsIiCkfq2cy2HtVr0SDXdzlWvT6NN3kkKsyMpvA2aWRMHdJrmtvD4R7McYYCyEA9ZZEip
0WfHUIC+EqtLF6+9VLRp7zkIYCdV+kUxfZ9p0wfMz6xYbzgLAZHnhvCDhbVFexDCicX+13qp4rOr
dYFS5jOdjUf4cmbzwqk8goolu4OoTUiLbKJGudJgXL91ZrmKEz//CCme5m5MTPM16+Y4TNhAOim+
Jj0Xc565iuFMlTsUu1FxjraIRBZDRRfe5w6+aQl+TVk476bxblV6RYEoHg5s1SB9Sm1bNCGRdyD9
Oa+o8VUGaqPChWO33Kiqcib7GThSma2c1t3NgVtExhEW5ege2L9fVZVQmpUUu0OSeqFuIpLN7C9c
X5mv49v/VHi/7BGqlvOvwwwNeSgCsw+oFjT4szpYvfgsFUyWzLkzMb6m2Lc9zmUAxgfb/furPVsO
cXWI+t6VxzA3Srdwi/t7nGsRbzJdUv+giMrKINicquleox1/ZxA1FOTf9ebODcWrp1b2rTdDgl24
o7C6wC9gIAJ936G87hSwKBDVwxa8oj83Kv/MEIaRWchrNcLQ0c4sWjOgC+td8zfm6Fcvrd1Fk/gZ
5zYdVJ+kPBarTzskmsku6cXvodi/PO4e6xqDDBXme3lKLRVTHGzm96cLfu6Gx9kK+UemCtY5Sjcl
wapqK8TON7syH5/MwErSmdHkfFaLnBfYXrx2F+OgFwBQ20njYD+G7HdavE9vwTuhnNH+s1CyuWCB
G3V7DiSNksmnL2ubEkTJf2f+YXLRn8/QQh+7TG18RGkXtKoDig9+NdY84TYs0LlJAibn2+OAIbs/
IsxsDCkDgmF6Em49oNYi96LK/fqWFkynuDgQ8VK8XFIdfVH9iou+0FeBmnS9PuoutE8nTCDMv1X6
YuvxIvs3iDh+DxW2sIjRhm6hJ9s+o7NVBstMkAwj4gPiA7SaCwsxMHo6OzBq0A06DlQbsTHA5UHu
QSF5qBrOidT2WgnALoST/2k2pDPiLkndf5lTM8YY3zuKbBzFANOnrfXZhOYFKlnXETrYSe1oRPQJ
egkcK9b7MYXfhoCtdK9TG3VP/mwsXKopzSViI+UGzTyQv0KSwIH6kObr6jFLbgUsfDbQkZnuy3m9
tB2uV/hEqjSDlv6w1S8/aNPlBguYab+vBSrySh558gn/sdTOsrskZ1Jtbl0VBTk/dhLxGARK2Pbz
N99QJVhx7OCA7DkofWwTsdwsi3QLSY+lN6NkFEfvz3ICdh3XSSTbanjby7ChnZv28rM0agwEwYrV
ZaQbRt7paEiMekUQDsw4N6zPat1NFQCbR14SuYYpMS5R1pQ8OioePxcahjkkEgx8BmAxzp6FVw2t
EOhsBpHsdb/xKx4LHPdxDiJCpEY9/rA7bQ/l/RsiiipYRIl0Kssu0vkEs1QjWgGMHUMs/l4kVx8L
7FaUUY5KAX6W1VQmQCy9vlxJZYNvP/lHWAvHN5HuqVmGawItSv5cRX6beu1xSe/UayQY1fcta5bt
+bzWxIAnXVAfEXQJIgj5sizwduW0jHv2ivELjaevKuakJ9I6t7dRwsFu/cINJaeienJdFDdie7fy
mDIl+aErGPoaFBGBlPEjIOQNtgUKurRlmIaIjBtGJBhys41+oStZoXZ2FzXOIJ1igMlAwoy14kFy
qhpfdKUtvvZfubxqrSm/bVnyBZl1VSb0l+KvWSTHOp9Q8ujhngg/fiflQZwgt770+Q/e4nXnRJ0u
wAN6DDR71IxUUGk08T2UN2nejZvzbIuIazgmVWYCJDF4Vo9WkZmqK2Za/mfnTW0NWo15E5/9tB98
vIVR9CKZNyOa+siO/ay6dPPPgaBxWgqASH4cf0zDnkdxiNBQTEtgG9Ho29G3iUzHim0qcUzzAtBU
3FQ/Y+CU6kYCwQ3gBWI/q8ht3GfMOshwwVkhvA2Roic/QA6htrtSz+ZBxFU3u/SmELl+lRSTEw3Z
kSFluUWVOIrcHYgivM8bTEVyf+nMatW+UYtrLL5oNpdugXLpYzNuZgdT9ShT722LT1G5WZsFH0BO
949k1zm3sB+8C15OIjSmW/wsauetglh2XZd+nsy8NzJdcYtKdc5WWJ9JcicBg5jKo+xsZdRylpif
6DdQeMomgRrndqeozafqFlChEQDrnK1mSSHi/fEP09IwgpQpPjlOYuAuokzUG1BHrAkRBmopkn7V
J67ht1/bF1BkVSICPqcF6XJKB9cKXhoCKqjQ8oyaDu9wD0h5JN3xf2s1zZAWS3wOJakg2oifaERP
rWXNrSC5xak2JVhkd/ranZxfTuHYvnyjyTo6wUP5v2f3pUwss2t1H9+Mz4gV7P+ALaN8d+auaQHn
xIlw/zPMemGy/eCF6aK4Bkg00gTrWLArWUYPk8drWp5iRuh/alnjjy8Kdg8RmVBsmb5xoAzEVnqF
J81ssMVTD7s66IjW4EZrGZJztr9MEklGLXOl1PxijARN17k+Cft8okYzdxzw7K7hivbSp577lZEJ
1lOJd9tnXMDjMt+ah/ey6SGf2p253uALzFuj3b60FCXwP2RuNiu0YWW465NoOwbaRZpjbHd94azd
ijPlsspAR0nr39YjAEirRJAh3k3hXZ6zrRuARQony5Hie0U8mFImIckROODcsf53FIwqs6C6W13K
pkyeVTIipOtAVNqUdZdMbelmE/QtFK4G2TuipDkW1YGs2kZdngIE/0COcsA9kTZ87giq3N12dNVt
rBKbYzgTe03//3cM5D1cm1Rp41dXEU8/H034Pi4mnZb/1yS5k6FGrkUFCUHUJHfAuu4g9Uq99s23
6cpZkqs1RtCwAZyVBt5YAbvc6agNxuqPoDc1rUVIKSN30ySbXJwRHNsREZ5CaersJU8QMFyH3Mcp
DDtXBkalRwrhwt8/302U2tY8CcdrDPhVI5CmVbnsiYhhDdYJCMFi1NgwQTZauLAp+yTOV2XTqQKi
c/lOAaBvitHYpS/XEJCjwidySt/3UYAH+QulBZlCS5mKgoYI5Axqx9I9kLFtuFPrRwS6Ll7b6JO1
ncacHT5OP3XiCrrCZn83sbWpFrqXokyXsEH8o2aXM8O+qfIYTaxsBgF5tU7/3N/8kMlMr+8jfDcA
fgkB88mytfRmECk/eo1yxgpaocRHjFnXFiUlBMrHxP0dZLNygvpgCWJHK4vKYH35W2b5Ix0rrKaM
EFpSVVkogSzVj2S64xkbYQLb5RvsSyIV+A8PROpNYL+rwFDuMh+J+3eeRAeEMRCtm7scKb68KelL
X2YiNB9m3ie1u5Igcb1YSJU68wEDw/SjM4BweGcVSAF1uHHoKlNA4rsR03a81u0fiqC8G2k/MQYB
SKxeg6gp6XvaVM6ZnJroxzbCzEm9Orzv+uI87LYBcGfMfkx0+jvZ1BPpY8F/VrmeJ16iKb8/f5nj
N65jaiK6MQkp/LwTshF/ik2c263pB4Uup08em0CDYL8BvjN8q29robxvJBu9pSjkSiyvbMq/PSRr
u5snUP4vsuRvXffl0zscoMAxezbiGrU7tzf5qmOic9AQwH9rglrx14g1qQVgvCIJDCQz5E47ocdJ
BUb//GEiI5HDAcli+kGmsuPI6lhltY4WZG2mfmomHJHBMJEW4XOlbv+IKNruLZhmXXBpajT+lvmU
bP9u9thgPkOwWf/NskXJeIH1KeJkpE3gDXCmHFl26cCDY54JUEGISNc7qzxhf4wADb7moITdGlIl
5sKVobCERxhVYPbUW2zEhfUFrFY6XSUcenDn1o/NmZhVMFCjKS67By0dmSufLOHVYnCeNNy0CD8y
kzlWLnEHvmMFSKjXVVbVGl+IKVBmpummXT0ZZtdeslE7SND14FRqwOLQW+4SdoWwcPYjmXqgyZNS
OKW+bbndx2ButWHTCXAzZ5CakMXH6lI5sDVWDo1hX+52VOvN1uj05gXmuxLNfHnv8frP4S/kuGc2
wOo/8vhUQv8UIJX4l5EXguE1IW4E+9XxGAfFjlevsctVmC+VZZDlvdnX+Kk/DBMNJ34FhkMgG9GK
ZlexUoGvNLl5Z+lam4uZcD2UJ4K82q8cGwRSv+Xh4Rf9nggB2OeLirsmuUTIg9NvqTQVWti0AHdT
v/1vjI1Mk7HITNrNqKjnJefozAr/CmOp4EypteZd9KlWUS7Tu1Y2j/xqWzHclxJL6zsduNHARxqE
m3h18PPUrwKeeL0pthr05XBk4U3y0Ftw62S1EHeeYblxSbqYTKIL4kUc8BJkjzKscqcEVXKOVlLM
PbdcwNHjRSo53TKgwCLiPaSo9XAmQ1jmoGWar8Amvh+KaqOJbSLFGqCHT9bxjAJGjMg/e0Q1+qHG
rCGaHv4dm6FY/vudonQAwexMumQcRTICGqNrzJq6Xynt3/c9ZaBKAfSQ2aTddO5RLMfgPHkyaa51
rxSl2vJGtarBjntRQrTvmHbyQD/cnk1k29BFiITP0PjaarRdtSz47QruVjK3JsNdwbO7vlZKI1u2
XWgl4XBdIfMvyneNcX1IcJLQ8ExHC4mfD/7aQ41YY93QRdYk8y7WGXh6s8yrsgthPcY65e8pHdtr
6q++Q3FNrkoWhqLqdYNDsrBk0ZuNoI1Ti0TPidUyWxk7im8cAndwhiykHwZdr1NzP0bncrub8w16
trxIReJctcNDtuVU+bW8+/pWGZ3+lMWxPk7EyZGctqKN5Cw6XMDgbsKN1G4pJn2f8HDtcfWgxeU6
kF+bLA698hmS2eoxl5ojZ8zrf4FFB4WVlz/oWqBzHEh2hoEIGe3v7C/qUeHzIc2EWu0qo65iiW7e
iD1Uvmx9YiUIexuVfbGxxKSlD3F0d2+T0BkY1QBv9I+SPNZBThFCEdHjv0bx7vQdLxXHpadDBHoE
Eg1aueSFVnBf4R8PfX9kvItzB3st3MfG41xI0rpoizFyBs76Fo9tQ3WHTx1WFnOixmnodRseSi6e
09fPLmOd1aMBaJxK4Jz65gP42YYt872HppcPxl+/o4CuK0JBdTqIvI0a7Iefn2W15Kaoae4Byiv/
9NuQrtKr43kg+Iixa2xtYg1Ns6zq9KAJBsM3dwXQDJDglYDg8veZa4zQb6hwm29kIt1vG0X1zss1
zgZVpoxlog5BDzlcnldcNL/L4Bx2K5EMPZf9/ZbD0TQISidPyFXT85/9PVU+pMY6ds6lBrapKPbq
jNYcXor4GjVWriHK/0Q9jWOmX19NSYK2jGdkDb4fxJScwYUlync0jHT8m1Y51uW89JQ2EYRBtMcl
fbb+kDBLu6Q6HulhtoY8H5o0pX4C9YmwE37gpd0E+G4WbK0Y2/wzgEkQA32Me5gRIVbsnb7fjzgm
PjZTBYIB22hL8ty3YP2bwT0paYzak78VLpBdJBxB0V50BzlYUEBG7/mIUew2wlBPaHnJkiWP+iKk
q9NPXlCCKbV/RofqUOuTYPZ8VsN3uCzbJ1PQoSPfzSaY1vUmW0TkJrTZk/V0iWIHNtfHtUjEvC4b
wCYY3uQZk5c/qa2Em6lDt8k7C9RQH68d5OavjjFV9KhTlWy/4MTkKn5qL2iT/wEBKVdtNkyRvwHh
nuTKAaUUopvyLzgOg00xpBB9LCSU+kNx2XvBq9Gk2wJcq9FnFsQeDgQIU8p+CAs9JHbk0yRHGLbj
tuNaAwBH0coTIGtMA1fiEZr4JT1oveqmrz0ODMvFc7+kvE4TdAenop3lTF+glWv5RdXy3JUexOAs
LLQdKCFKWbWnmWkCaV9eFrUODOtjndoeP/ToWK7wDxcOhNhZUnWob7463iOeEiraz7Te8wGMe5D5
AeypvUMwQF84FKxo6DglRz7mVCPc+0OPE7y6imS2l7qZ7FfDZ/2c+cP/5ZPFejFZuKrQOvS6Oysr
q4yCtwIaalpjqPNoIssXqjuIebgCa4G6AFdcomEaqm97eR8PnbsZQOlfVEFZ0ux39/K9sFV42iW2
04eVHdrtHuAxglDvh6A5PRelzij28gVHla2/cxgdCBcdbRDbQmsrZgrmSIsEry4xQntIPX+HG15m
T//ohJAXtFYzt9HZgxzlREG0/TraJdv3OVltO0lZDi17sXN5vlGoVhELuWw7PFQc7SCzYIV9kct7
s4qelz4Txa4AYSiJQqaf+NZ4/gFnFc/cAIEsgRFE8yGgiWoFCJhTTxY25WsdbbPWK9Edg7+13pfV
d64LNNx9ECf4b5liF/4SXwCc8rF/W+nvmCsfewt4NpTaiFd8aY9xIlY9t+Q7oSkykwQ/QNU9SKBR
wook8K2iqoifvtMcWivPMqmXE2WrRtqrTGJE+ioxYvhY/o/taZpBxcuCyXWzbXNjfwoF5pfSheXG
hOoHz3LDf/mGxY8r5tnXJ3JgMEuHYC6oOctsNitJZuNva9bjid/9iA0lcgu2eXghNQqjKRMWRonB
uP5POAahp+iUF2dfjq8Ogt2fa5yWamTYCcQUne7a/7GXcu32UNHqJpVlpK6GuTOmOFaEBd8YroBt
NrJRGkja6Cxn5tcM89fms3v6kVTxoWhMGk4i2MMNEsOVjpbGm0TabEuBSdjYaNPtShgp5Ux3kl4D
LETrGGN0oY4zAPu01a1n8BGqDt8Vur4rcKB+MYGWuFG9LTYmMXo26qemqczjNuO4XNsVN1EIy87B
EHS2OH2Wh4xyQgK4HU/VU6NjR1JQiVnUf8JmKWnhKEjkzv4RG8sOcrgN+GGlNT/SDyv+PpC0yUyM
PPyc9NwKuvgHWJgygzQfRNnHsGjLq6Tkwxh2rP3lGsztKuV6aQ0iJ/2gDNzPGUWZXiqMPO6Qb8Gc
73dECE5rY/7MNXlfOCT/NzY5zqGlWhsOcQmuKgtSSE4bGwLYW7kRHyOyx8XPePMF6HpZMTu2sEqh
joh5yU9LcEQfVkli7TNSSUyQhp3Un+ewq/hmc8TfgnoNkLfdXnNasjXwir5mQhTHnDHtZeZR2zlV
8/K1SJOatVRlMLC+SkNYGK2Uxp7ljteYQVsARToXx97LnnmPZOAIjZNV0i9i1xGeVD5jUaAnasEv
jHNL8f9/jIM6m5xo4vkQthEmfczaJ3VljSDKC1Is8uCkj8ql7gi81vz7alF4P9KOHgS9MbfC9+2U
y9g/pLoLZJIPvU9FZrTfP3hPLQExxz5pHpM/cSdH8kr+FkrproO1Gix4w0mg02gjaA/Dg0XqWS8s
q65AqrCkfihSamj8qw88UFA1zi7gRCKtLVjKeyg+lwvNNWmYIXlCFh3XQ2IPpmO4tNTwlEf1fGxl
Jx3GoKEYg8Q28ROOhjkwpRjqEla0/uRmUBby4YjClDVAWbY7XworTUvxBLj9lOwCSpyugNqfvt0D
gdmfaivMz4EN5A/E8qYZtFvPRb/CQESULnN+4HA/2cqE4Ejpty6BAdlYERaFvuyDPGU23YJ0fsdB
rFeQh0rp69/9FINPdNJYm0wei/Zl+gozpIPMuxUnqbDkwZV55xjgrHZkRD932P2EeUas5JPNordz
I9piphlK1T7g4h/6vW+SIO5+Ls3Ge4uH4F1DnfX981+FX8xDgaDkmYZpd2Cbh36PZuX5Fuyw1oDU
+UhDwmOCIpNSvkNxLeCf621jcDROdcqmwsdoSPuqBCbVnfiBUj784CKhd8/dggIYddhm1fYJ5vF6
OjiHHPhszew9t3+BOL29XAeIryub5fy16GzjyaT/jK1L48SuZlkdspWZUQIwR9uuTHs+aeWHwSjy
j/rt2i7/mm+m/c061B1C33fB35+lnwMy5OYKRygDxGXGyCrf9/zO4kl2pghEMgDgZmaeSR1iiPEc
ETL+Kqb6J0lQ5pCD0HpK8iFM0+A/NfAaPQvuisMPp6yJFlZ8kDg2SumTc6cVsSt2iDCNiLmS7Rpn
Us22Z/822YKYBhkaHkaMu1TwKNaXnnzButesrQDs6bWGNjQFk44LJH8eytiIkeOyJILyeedaT6t9
DndJxcyfG6dedCQ4zGgQqrYXbajkMEj0HjfCS2A6ke9YBurcs7Jj9C9wm0rvxUqF0mUNNVkoAY82
4k1fwfukds0T3UWNE0vZ3fxN+QD9joR3trVViPe5wq+6ynL0vWlQKwI3NV9Fsh/rofoY/15h+plD
N4xXAhOUjDsjXk7pqPypxSSCcKMwxN1jwU/EurVhDFbwoasm5j4n5cWXISo7BrFPSq3P3pTjV4Fp
L5ZoOtCf63qaaPU7wOio8K2OMUgX8GuDSZF1UlyF0P6VReUWB9ZVZJKFM80EZrv5CwOuSrAKEVva
qaSRfj0W/kNHusDJZKLAguDIsYHWKGXCc4ihFWY+ED3N3PWyGVldQGbCbWrBFS1uBRbQ8YTcK494
r63DRH0GTxHqhgOm3ggn5ZsWSgngPpCVPWx3HGJtTCWeyIZ2OBUc5Ech/sj0JmYvuG0RXVh0ilZj
dR9kLnqYUwgmAtAY6CyvpdkEvqrKbw/+O3CgVhiwxbl+ve7aLUKXRCMz7ftkyu7bfJBSmJqJ8uOY
JQHiUCc0PqhHZ8SQiGCjSUnYvrtDWeBsZKeT4lu4y3iiW1y9pkDGegnnn52tp7VvfbAQXqjtHvcx
dyTi3n1rmLvYrWLSZIMSnZ+STukutF/oh5w2zSayQRdrJLRqxXKN7eI09Z6KXAg/rY7CoiiCiJ0H
VbERRPOrIQRfa3duYXBGB+OXXZYqh1eNA4D5vdn3w8mJZduwBz7maC3x1bOuDzWPTt4JjiYaTb4k
xCHzavoXexglnLzoDRlXwUfxQN8LYmeL+V7vFd3kttrRik1E04Cz1MinXQcW5Mepk71xOFGXqcDD
SHR3aKYr4IUI22TT7uqp0jz1X0+9XqYZU/X5pJk2F0kxNYggewi6ogva31EIbV4DDGU3h7nn1GCs
kuX3F08J08Lkbk4rc44mMTtF65Yya1bAEk/4JHiOJQw3FXWHaoUaSJFkt/nYOFqtzR9INeEIonK4
SptH1aT28Rir+epe/newcwpfOGorncaFnEQY9tLOv6ID+/i2vGnD8WEh/TcN2eT0luln7SlymNMr
hiM3kt5URhjvt/5eLeFPpwPD4cXyyVER01+77oVRbB6sPrH/3NWqzi84GhHo6SG0JhyWvg5eJKBy
qHC/JBEbca2vJsAmoPf5cv87XMQEa1xwK+gMU8i2LFh0aHkVvWhkVxPskHex+3QdwkEsPw6EkpCB
1KblNjXeE+Zfid2kkTRZ9U5PF1+V6wVAoSe8wC05ruTO1XcgLQZ0qGXiF93lKOJjSxp9K5/8YBN5
xpBQbFNYt+B5IE3/+shnHyO4E3pPxo0tJOQZLB6Fxuzcq7kL1S8g08k2/GQyyiqTtJfWxCiyPmyW
cITyHNHRkho79mj3+u95XUqlGlpd6cu58v9qfF5BtDtKd34KEsZECEivMI2AZMkE1F3DEtgnA9hG
xeNWFM0GKC1mwGKe0uhGwqCtSMcZUejmQpGhDp//RunRyz3HVTWqPEKXxMd34pPGiS9OdHVYcqSu
X/nosESszqr/VIcPkly0f+j0DBpoo0kbFMTdaqsMxKRXSpYV8y9/Q6LrjBUtfWnZcVA/eIb1RcQ/
u11QM9VKhwpxzgbKb1heR1RsyDEhRuP8cLrt/WrAMtBxjlkFz1AMMu81eXWbGiwJgS+Ssujh1ICE
S0IbM/F/R8KmUmovkIVr0Dekh2e9686H9z9p1jD5Qv7LIJ9y/eMB7+NawdXw+kG8uJGwO6zqPBYI
X+g8lNJatGU/1nvkJkp6kP8HBgAqziQq5IWG/DBbfKte1Ov610qa81GdUkqAo+b564zFVlLk8DL1
sywlXLs0Jd+0OT5ByJQ0OiTlPB09kF9GIeLzYce1XN+Jt8Fuf85TGpLDNMYrGteoXFu9ogUvQjuj
c9Ao5PGFWx8hNzef6VB4j8/9Y0LR2khfV28/+XUB5PH6Hwpv1UtEXAWImGargS+UL1IgyuPuv0+C
GaakrH5No3Xs/zjBQLlZyKEArf8fqIge3WBFByOFSv9lK/+BcKSI+E0nHzCrnBMK6XRLb3gX6tR1
v840G/qUlstXJGRpsCLfIizWPnTXS/PxxNmk0dagodsDJYvNEDZgcT4JoiwDhG32y1DVXZJyVmp8
de3qjs9Pon5ksc8+er1kh1wBVtm7VQpeNO7IwZrovKGKachgETjGtygRI9onYD+iDXVHzaY5ghiu
RD/imxjMoAOpE+0IlD4XSAelX37EgeTFktWxI2z/lT1Q328O0re29H043EcJDR/RrJv1EtkUsO7F
kMuKMTAnYlkyhKfEUXZMNCR+/uiSw3qQHXV3fV1yjvnWWTAvbgIKFfobI79cqenythjKf7t7EHVn
8ightUsP62pIZtH2t+0VtGCdtZUewe5iKeEmXqrcBCU43lRCUF9XyJam3BRYat2OsjC2Q/op4rlN
za755p6k5/EKRQYZpmWhQ2PV6UsHSgNvRJ6EZy3hCF3pJf6eGJy5xc1GmTf6YLMxGcYBblQvDbJb
vXLrNuAPvBwzFNoHgCoEmhODULFmYAPtXamsMmKwjtVgMBSECXKGIoQIlIHR7DR08lw9r/SKPt6X
pD/S1YhX4R/aYSKFbTSOfGikqBq36rGTBAIdENVyOIermVaJrxWlS8oP1cTKHdrU+UPDlUYnUNu5
xigsN0D/tqtnL9CaU7Hvw0ns4bjxbl2uvPpDpLZR2S3gORiL/cOdHhcG+mQ1zsZCDo/Vb0QbE3yo
TD+6ZBUukzPSlgR7aiivPMGm+LByHQuZgOb+0p6kcQ1rfeXZ+FVwvcGfe/DJA3Q84yNBRsyp0MpG
ujgKKmIKxuOhFxSmt3vQRSY+ieXJJnkb1Af1eq2n+Aw4a1yJfjZ7GUldsFuN/rzCwVjI31sJQ2z3
yjBJ+6FCbKNgBGT5sk/WGniyzGyA5jzSB+gIPvyLY47dIfaTF2H1xxnYOQzBO7tavkGNG59ZFmPs
0Gp3YMqJERLiENYj7WOcuV1Bz4KOxu+E98gUeFU3353XgijLYH9BtGUaCJ8/SnNRoP+Ql8mQnCYR
LpBRwRsiUBzD2/t1uDHk4PTqTgGT5bYfbcLERNPnQSD+K2Jn2S2VRL1avYyAE43Ap7G5cz5YLrYC
wBasCBBV8EUALGZB+G4uVnYDWfRhUaTtsEz6zbRUy67PNBeKuDi8myxoTvlqhNlGt7jpGwDgPKce
jixnJIMdxpPXiQWBoAGAF2woZ0aojqscvIE+SBZOD+yy62BNccJhm13Oyn8SmkAOHH1HgQb3w2lw
M57yVTPdXX9Amsw1iJyrYbw9pb1LC8Yigu+1AUcghWYiFAweXckcuNLzAtp9syQEHgaaSkdy59TG
CsFA5NJB6KB3fdIbwf1Jk0oMnvdR83wGXQg/VirM5VgxvfpA7g1XQOdDYSQ3gjdIGo8OWyN1WMWq
SCVEJ6Wc41Fwp/aGYCxLA0OlfTutT/npz9wAELXZumxgAtY4mFDOr1UNdxOwYpMUDB6EJE/lEIee
ezlURfOEyf9Lk/ANYmsoetbo1StD9/el6nIQDZ5QEvUy+5bg4XLEsv4BViVlob4OqvLW09U+ECyA
mIlg9V9OEc0Lu9uRylLIvgg4cx0Hj5x49ULo9YP+R2k3r9RyFkDn1QAWJ9od7M01RR2slExP49T7
0H3G/u2gGgum01ssD+tugGALvhrg0/TRVC/H8sIt0tzf5LSu3j6ucKdA272G1uwY1TjLzCbKO9NJ
Fbs5461EoBdx5sH9duoAWRTHjBrzvWQKvP1SjdAaYduAGT0NVXbDs14y+OAmC2kJjxf/WBYEw6aL
w68rToJndNLuWE6BQMqH2ep4IrLj9SU4Wxl+Ozk31UGBokzDnKm/zM9ZWZJPerqNopbBw6nIDAsZ
/ivnzjK2PsLJ+mOesvCTNeO9BOjoEmOt2BH6vEprRqbJn9qaXKg9O8SCI0Gu9IXShH+/53Kubq0c
C4vRIGj2Fxq0qSq4YjIwaPVVA9hv+bxJlKZrdWhyc+jr5A3aluJ21LUcFFSHc74hyMV+5KQxhhaf
HpDzRb0J4hLyOmVwmZbjUnzxl9anUhJ0w0PIkugIh5lXdtjNmsDcOo/A0yaZJMbgwVPZGXuxSSd0
9LxwzNvwL2K0dnwfjr2dBAD80QrDiISVhaV0wyHRq0grHR041v4MSip22W5oaKT0ZVttYFckODMZ
Ega8AqubKpmuEOHWgJZ1lDuKC0TUdbm+f0jOaenjkEGdnh0kl/ZY+bpFdLmjH51Eal9aTMpdMS5e
zvEhIbVNeMGn7OfMPDwXzTsDdWBiN5senlOYvHkgoMXsTxCG7q48GYnBjJS1h/Wfo5s++tSz6Z3k
Op1MMkM7ZNy87KBAnk0rjOeIgdb+91Fom2MJjdhsWxaA4TvybkspvDl42iehXrfspAcFDee4wlXJ
weI4/oaYu6KVFA0lNdOLMCvqVshrxlLfEVsGC+wR8cdR09zvmtZ+jSyBMUktEnkbdx9g7VoQah/+
ABlFU4x7M1SufjEvp2ntzl4f07I1lBnJO769JrAN40NKGZefI2C19iS/Nh6ZWYmc+QON6XDMHvWN
t0V5wpg/Qfl92W1wH/mhyT2Vuuda51+WaXEE5uuIQ/xcmJfvSzB9Wp7tVp5bIArXvrssHdI8KaAn
BfwCwMz8RfZWCMctKy5ln+lrI1LDj068tH1fc2OEgZP58esVTe3A/PznyLmWII8bG5XEeaMhaymk
aMITwmHYtjXzxYwiEBB/UFYMRsRzQy4NAglx1t3Rgokb6il5f+bpPLO0OCncb8Gb9EOnZY4FFkm6
KpFczYfcVGUsawnGzEA0OBM1559bY/LR6mVNYJmMSGZesnzGm/O/fNg4Kej/Y5XPkPYuLmPp6hTX
rxeaMtiMol3pl0IT7wxkKprtoKQIiIiIr1S0GP/s42QFZtMDLfVxAeXd/qzIfF1vd+jNad2BfNQ5
BIwBGu/OCRipzUlQXSKTlCroqh4LM1BHUcG6IU11tDZZwV0ReFHg6SemYKrApk+jh6Ze0tAGLBNi
Mm1Wvbr1dXGLYXHkeD2bUtPTzIAnLpUMDfAXPeICeWMH2kYMoaKAV/Qv6VcZkR+NaKrHGDzwfYPy
M+Kra6lheBi5QYK+AFFQN5EuNkJ11clmUuXFFpOSaeJmTVgkHX8A+UlKr+gCbjd44sG8jpReJwlw
eZjs+DoBymipAPZ/8mneu2x6fySqIdbo6jd9C0BH7SbiLreqD0ktLZCyMtFvHo2ZxCXdMasTgL88
6Wd4PwlOtFMwRtQJdH8iM6HZ6B4MRN/YkZ4/PCf54m0jtQG7Pl5idGoBuilqtNZn0q0IifHXYyH4
vKA12QW0H7xuradp9kBPbfTsY77pSq8a9xemWce5xrXKeoAsXPmNJFMGoZzYo1k3ox+6Gx/1LOZF
l+HGGG9/hJzl0UMgVGYhP2GYn9FLDFahgrs6Oav+Cteq9JdEsl5HNFir2VMapgmYyDw48/r+FTUO
qqXBCmkXBrdhllpPL+No6RLHQCXDHRKcXftPrO4iXpxJ5rnHCN/8Zhen84XdrouLEX3s0qyt0UXc
6juhfQ0jqA9WQXSufi1l8K61bSGvRyPsq9vBipUXlBOjuLBnseuLusg8hwwuNHLoA+HlwYiaHbVk
CEw+bRX1WFUsX4Q607MyUxPzlonZ1k29JT6pg6b5VySVlCusboKTRNihMe0tPdH6AvoHJq5CO8wE
1o1PkP+l4Wq0lXhfUcHzRmFYmmvIJf+0yoBngMTK92PeJTtCJHrDoLfR/rrQ6hB/7k/2g8S8MrsF
gfFAO4tEoV8Sr9e05NOtQsWMYC6CgafJJfF/uMc9SPVTHjjp7muqmRp1BKGoohc6dQMb32K5RyVA
m+n0mp5if0WqlloiNfeWchC4Z3kO79gN5hDrdDE/P6Nj6Hqh8y9TGizbX3L40Zj3Jq9qj62EmWq/
o4QdZqUIK5iGoisw2dTdhbwnpp4HBzYgTbN8lYDF+MUgydY07QOcVqpEwJ2rJyrKQGs3UhZvyKwC
NGMMb7dfu0jDd5Ocq4HbmqIZuCVh4ogmb7tniDz9hWkSvLR+c1SL0lf0q7l3C+wW09ImcAkA1780
ri5C0/PC5zeVFa7b4soOwelHzd97eEPVHkS5DPnxGXQiYH/XrEQAQCemjt+ZqoJi5J/VUyEzhZ66
GSdjj9jqFmSxEluxX/ezhGsofTu2nJ+MUWddJIGJl6PHGLsMvMEQoP/LzND+693iqg+oOh8ZDrj4
4KAWIx/rBqpIKNK7qkxJ2gbvi+GJJzIbFDq3gM8XkdReqPsl9TmjplKSL73e/LIe0jSdfVBiOC7a
oszgMgb9G3aPwyt+JgqmybPVsbUJWL96mA77OoAcuOhMRtEmyDKrEVxp3mUW5dPGXNrneoN7uMFl
23zdrU8Bv2lFtZDmfic6kwBti0uUAaUsjVmvyWIqfUop6hfIJt+NgW1EqFNZieklssiLfgWASHNU
Trc9azXlKSeLe0u9nbGOx595+u1lqR4CbzEUhZYfNEZujRh7H4SmO6/CqeDw0mDxgE/y/GIs5LFu
p1wZ/VgTEAnjfU9tQv4+ovqZaZMUhs+d1G3simTi16SuJtX7I3coeGOUEC+wErf1rTUa8Z5NT36O
3KKO4Sugn/gHEkjDmtZuY9AeYBX3VsJ9KgsJ4JCsqyDK/jseQ5uzcjsCDgQgsIygYJ6L/t+c1j/i
VlWC61Na9zjnOg7eEDp1NS+AMD0MjS7oV0uRChEqXXzmxMqDPe46QwiproBMly6ZAiiHvQjr4n6W
JM9nAnjE05C2jJajSSQagZHPbHnlcxC5w7kpGtrJW4F2wacWSHs9hpt+9D9N4FrFiQcsFahnV07S
+Fe4MUEjlFMN7TTq19n+zXO7L2b2jc8s6wd9O4bOdT5sxGOwhaNiCx3D2bIwCpZ9TjbnoLcYVrjL
ckI/iQzK7VzWTihh+qv/fGVn1Rcqp6k+/LCZP2O3hlxXMJhZsA68ZWCbwK/S7g81hPnQ9BmnMb9F
mrUHqjTlkl8oGmbPlBpZXA1hkixMSrj/9tTiuz0Fl6KwiUdm7ejZt4gMbiExYy1OSVV+Qz66coZi
kOw2ZAUK+CvMFltHPoNd/islNtqEyiFZH804t38xd8Ebi26kO+nJH3vm2hsZR556thWyGOE6dd7B
oJLtBYoM0tpH3U1tkls1Oc6VDbiwNqNMZ/QSo/C6Hj4Of+fmwpCne7MUyKWcTbgpiJYEDA2SEr0y
MtEa1FI97NQkP1TEMsF0pwA3InC/3pou5gp829riJZMeHWR4TILocadcSdUfHHakBSP8uJIXCRvg
UMj2UH5VQWi4WwqCRW5NKs1agGtpY/vqAYfEnUZt9Kk9KPSaGs/SZ1yDPYR9ZpdbR7NRYFtUrBG3
BN6bGrC9Ak4hAkLdcUx71wkzr7BbIoxggkrKOrBD4CtsWfTQmVRV9UwNXhRItspfQNqaJuHIiQav
I2QetG4LGSVQ37pd/RiEkn1zsUXQJGVyX3QZWxWjZNv42P/tZoL4YkfYUNnHihuL7oiTCCZDDGAi
f49Xu4KLUz6kMf5ywvNzeOm9PUz1sQQAQmlfJWkVFhlye/B7YRkJ2jmLGUQAwIFkvAXvJpLTYXxB
fxNvhRL9J7iGYpqe0LQxVxjCBxDvbM64R3E8gQJ699WQBGn4ZWs50o60xYobkJwqoWYAwdAKzhUJ
5Dgf9T4ygs0YxWqTXCOFMQec+67gak7Rbj0T7OepzVw3CkmdP4qrpE91Zd/+aVoHnU2uCDquPOmt
ZkYJIV+Jl0BBily3T0D7+q2yMJTHn2d1C/kxgEE3kvbEVhdqU+Jgikl0tcD2ws5yfEUkDapo2Yy/
rlYWW+pSFxL117ccoZ9I8wIXX9pJcF5NWUZTHFSr3CVhs/DpR2M82Y6/oG/NCY/IvWQwmvkcaqok
e2BsuBXMZP2/l52z9e9D6PLEwnO5HqIYFAFdXPaK2YuCbwAsRK2Q65426llxwLvkEbE6YrZLTuhY
OqeM58Puy43OxkXS9vHg5rj/g5T07ZFktB1gihcOSfiXaRfcm0ojNCV7ZMkkfIeflcpeRjv3fhLW
mRoJ2P7eVzNAg4PYwDjfDbm1mQn1ReUTT8fENLc+tZAESHT9s5ctFRdLwRF1GyFEHwx+gLWlHP8K
NLnizs19X5eE03lClZrqfxmGuvZXTPkwDQJ5aidv9Z6NVvz8eb0G2l2aSq5HN/edpi2oBWMY5DTg
a+zRcwuEpDjlBDBRVpQ9ejYf9DXquprBn98gS8c/QghvOfzU6RzeDloVU52GurVBu2RUgZss+h1H
tHWinXJtphxHc4kl1/xHPXivhfeIWBK7bHQVjullWiiM4KExnMgZs+vq6I3Nr1Man2srmDYToDp7
XgwD45ZqeseCpCBsrip6wLm6ZftRFxQEoW2cNzaCgpE7lbJP4ptQJtK9TspiMAzPAYsXwV/iwEAz
NCM299MGaY/k4PodKdToCQE3p86eTsR41swyFGnruVIpgAdSXqzo+2+NBNYA71Why3GeMqC6WdQO
aTkw0i6uH6qUVc/hkibKws66hbDkn/rl49D8fyHh+dqqjUCcvARYbNiDCNxm1nNuYVRpOVPq2rYk
CeGAZvQixdKmzYEgB9Hkja/M9w+tNb6x9MrFXyyIczq3Ksx1TAqobpXlxWTAa7GVGTHMALV/RFPq
fzFiP8mTn0nIX5XpgKSWj+FJVkKDNEzlpiLj6XqcA4LECUGY4pS18JuQxpJ0eRWsTDp9gXnIM7wP
mJdoqG3kAm/kTP4itbw4E1thfMBMf+aCI7adFMxa/8f0f4bLum/P0fkqdSHnZdCLWMxcOVFmXPMC
ruguyi5aTRH1pkZtTd/M6X45+DitLYX18d2dUSy63+dufxa02nJDejGVEKYrzCFBN6CJcUJScsCi
9YhJ4v9HsOUzU2/XhCjC8bSRwuvsEy1dLB2kuYTNXV4r+3H0tQImkevKanL3bHTCYOV/fPAkAn+D
Tqxmj+K/upoB2FbmFSqa2LPKIRwA9regLgW0pDqRHAHkFAj75mbNTfNJyXov6R9Hh8Lubp5Yw+rF
xJYbPD67FtbFXUGQowTP8tIWjg3F/NHoeG7w6RccDzUjGhOiu03e7Zc4uk/tC3+E8AEwWtExtkYP
W0L1VyULK7PAfhuCaiagAypkxfEAiZwlRmQJLDZsiX0awQLFe+s/IHKPiTX3QZXpTltL1zn/Q4V+
epz8VWoSzCohkRFQdL+sUzrl/RcIHZI3u3gXdTtZCB/TwRcqUZBfeHACwaCX3LcO08dEyXDIh2pB
UvStW+B5e/6MbaeEqecrdH9VCRLKKWh5ApU76elnUNrA7x+o8h/Hww3nTsYW64fKwuZYcnSoUwwJ
MqBfmqi1FThtI6fiTtydeXGzTkUNUThX/KTW6Sx1+g+wzSTCSYxbvqjgPxFt84hfDhcj/q1t8QOT
kGUNtbztB57qMJlQbi74WBhCCWbLbnxJJfPw9e4G80+8Vdevu5G3Rg/G0yyQ8FalRgQJ0I81cebV
p9Am55dUCRg7cchWq2Oy96vfplIuIQKUi1Br7lWB/SAcBxMVtI4wvSLUeXc2exJxEIXDLVxJGwWK
wHXPxSV98FQxn5QEUOhC+DsSbJm3qjlb2L0/2MEf4KUfjy/g7g0eLEqr1BxsfIo5M8BCAlwa0t+J
fy2cnsoR/GiwfG8blsGxB29YlXaGRWlJ/aUIBLBI2sZ+XPeiOest6a7ChGlTiZWuYHoTTuxgGhMR
S14YvVjxX0lFBxHt8cOy8jxbetD6XfI+FrXexqaqa/Q3a8MlYFYc1d5Sy0VCQ774Rcq+TJlUi9kS
i0uygQuDDkp9MItkL+fbKCXKJ1wRUjjIZaJHLa9P/FxDBm2gFvMGg7IKk/CXbeFHvIHL27Rfba9R
aufTY0l2KxGn/PQyZQY0KYKHR4T1TXlLZBpgaTi89KryOvQQzQ7lopF4MlWCPpMnLeHIAKQDWPpD
wB+IaiE3CExHApc4FL5GSq7o2dNIdvdz2bfMMx6w7fmCiQ1jQtyXZ8nDhqSg7EF/M9cBn7sQpzWD
ItPcvzzt2G5472dQZ6xUoHg3Hq9n3WSzCLq4yEuKPOMXIfLIwaMEgWU64jHnJL+9jKY97tmceV2w
KE+KSzXagYo4cJQgV0QFgYP3NFqecdPslBA7nGoX44gSsAEcphzBTmUV3jfPeUSkgfl7MedGmbPB
1lDddSjG5vNVfxDyc7XgkBmRsP/E5zi2qOITD5dEzL5UjvCbFwxNcLc7plEp7MgbxSowB4HuwlAU
ft2MJAKEk9quxTyCIroAmk2oJheNvE8Rph+FkC+piL8+xputfH3PB6l5tHwTAdUy/k4a4/g8qLSM
KKkmRatu48w0rgOgS0GNVNs6zpPjKXx/tpJQFCJkEytuIYXO7XVLEmmbFABikVLN84pNqs67NB6I
eZOjc/MBRP0dA0U20xjDoBHuv89QXmF5T4rzft5iwHEhXOmwkduL+EJqnxuR1ahosLKU+wtREdtQ
vwb6Rq5GBs5yj6FhGUFtjrKGDG34WklDsDzTBN1ce7ktuo1jlNmUL17CVrtwUPi7lFdo4Bi/Apr+
9+Z7dSGKHbWLGm3cyfOlJ/0jVvO2lZFqMJjt1Z80X0wJoVbvR0lF8Kvu7MTfGNxDpJ2fbJEhr9UN
biSf5Wrx46SeZJEljAu5t+VDNRnWHqP2DiXjxeaNtfr5PzdlJkgQC+8e1ubaNeeDvg7hIm0wBula
KQD/PXOHbUzGuEVPgu5DkjiskC04vfe8+H1TTf/rmLxJisRKlDq7mI4l+q5dFK2yvNj3Jga/eCXD
ED93ior8CLxgGw8tl0yVGQcHytPyjTzsdGZpEj3pVfHd/xfh0EKY/I7/8S0fYwcK94RrfidXyQX7
kSti9eM8exRdhv6We6sMwFoIXgoiCB1fkqDAVZrH3fBhT2GhFxJhjHJ4ew2CDYVRs5a+7NYtMqks
GwNdNJnX5iID51pFnxlblHsM/cihX7xElLFX495hxdKc+JYB9jlSL3XjVanXWcNRkk2AgubRoAAh
XSdiJKth+TvpGYOy2hP35C0LqIr+NPYvQyx03RUSwqHFwEIcjxXPgkmyctaj2E4Yi3dZD0sgc0k6
hPcFr0fQqcpxQUOq1pLThtUFOf5XO8XRma8NAgkanbTma/BKpsJeoezPRv+kc0zMUWka9VEi8Dhm
h9CdThFH6WrMo1qaBUXont9zdC7QCmwH5BlUSChoE4tkkGdzElBYNZbq1rujqT9Lyced5pkCoSOx
AjBmOewA66qC/x7bFonxgqzae70mhvyLNcEoZxpT67UxOVFIx/sLUULS8bGY8J7MPFURHVAPZWBo
Z+2eHc8yr3MQsZW8pXJgJmQpWWQ2fqDKgBYLnbzgslQMvA+UXzg2hMKp8XJnNL/120UODEsdyEFx
d9uSvUJdSgWqZ0UipAmRs57ATYi9bdUFxQvdaPaTpo4kC5D1Af1Mm2wQC7koOSE//OEcQr3FMMac
3EPM1XygOdmeZZQ9jYyLkAIZb12Fr0gXPXH7KqgFvR/IoaXoYNtaFWn94kCNd1J37wTEYH1MQDej
jM6VJhcee9SLENsXO1WrpC4EqiR9COpaL/OefQIqZwQTuccWpzcpYQswogxmVvY8QZ1ur7mySus2
eF3IlXKjYUjBB8SCY4S6jgB0Vtgv86Fd6xS7mS7csmALNnl4FgV8caj+ddVyzbfD9Tpf46MVPr/3
uV7ysCzb/icRuu9leNfw4KAGZABjlAgCE/y4sl8asoiw6tjrRDwge4wjfY76c3Pd1KyEB1mr7Z8w
HDDekReudwBOAaj91jZVjaYfmdYl+TZybj/IwotH7RlMO+Gb8Eehp2eKq2hYsC/lESLCbGyVgIJ8
OiOREf6cde4PKPDbAFT9pR7kWNE3De+Y4DplCBPnI42Zg1qX2AJ/1mGDORNqu4cki9YBuZxwV625
yzPoi1MBoeUts77cjQu2KcHq4iKmQO7SJ8xZJltHelGRqF9O717SHmb1ziiPeamBw2feOqOLXiwx
D9znRlMHXO6PAklSMzm3W2jA/UD0toXANxtVgtfznOSepLc0HAKgPRnuoOIHqh8qFWzwadh5+vKE
nNqrrXNZCbNEYP2ymGV4F9KfHL4s+ZJwzDvs50JIHT8iepujcguVUEqgzOeW5wh56+AwiRYnfW50
51WXJxeL25mXz2deI6QQAgP+eD/VYHa0Cj93JBRVH59LZ2mxsC7qSI55m87AZCigVDLuNCUHYyEz
eMre8LTHlD3lWf0P3Yzua7RiaKaimLmulXdf5B/PAygOmI0EqRt8bckGttBKOnGdxIW+hPy6j3VY
dggIR5NjaH+B4JVoNHuM8YCX9AqYz32+fsWpzADypLeYu4RQd9IFIb6uasp/fgWYbu2sBJsIXc9K
y1FEZZf2+KxhhF9f5KVzVTXU+IeRkh/Wj+oKf91ZmYUKwg3MHCX+p0h+DHgOvGqxQZ0mwAEPDjs8
yZovZ30uxEGrG/fnEqPF9TWNkn6BSFj/Eig5Qx5zzXTxMRq0BzHStpIfXasonp/wBZiIRBz00V/Y
ERIWzZrZ/tEdNJodKXdAtdCIiwrz75L+frfVYpg1ZLY9uP+nQXPD4ALoKD/bwAFWGM6mGb5DQOfk
NB3kn9/TwVtpnnRX0j36kSm+onXrLDnWuvxoXOuEpFDfYM3l+zGLbTrQabmZFQw3be9rW9EYtcMs
P79yBWz2QbAEU+kk2BiWflzgk7bjLlN9CiNlay/D8gtgDx5GpEICZ89AdKvpmW7dytIsd+i/+nWE
ArnfzCtUzPeps/zheTxShCRbLtUsf7j1MPsQF3FtIDTczyaQWxH02LpIKnEIc6o2pj+iurDxjCMu
DGkiBW6TgTTWVTiy56Q7GnNTSYO3T8gdaoRuAi2/tSbpuTnIynQk0vvdRRR5tFFgoYs4gdJffxVS
Eyq+dyOw+aYkYuxR6b8SfTNJ6+nvci1Rx6o79B4X0Q3ddWQkKxfOUc6PPxbmlgADe+bYhrHqvyRl
dyyV6kKVsz9Z+AehNEi31p/UqYDQ1Jpwf+JynRoJjITcB9OmaNsRJ6qGYbu1sEA3c3DlphXU02O1
xenjRIzxKaKyODFOyTgHUMZu2A34Jjc+F1KzhsJdGrWVYoQk4U3xfZVjgKTzlzbltGPVgW2QzO+1
IqTkhTHRwx2Uh6zt6QIZvyC2mwaP4V2U8ygtYXd1RtA9UlPTuFjjALylNs+UdQMhmvn1CEVOnhJe
hqzaIghQEMyMmLVjMvLkhDWGb6PcDIZgvMp0s+kIquHcyUlyTUFbFkOvp+pDB9niBQWK6t2BVCKl
x2Uk9DVuCpIWOK4PYRDWo9EBwLE2C5AknqwGJZkQACrR1VDnjPZHQwSuBjjJ9/5vpgjymcs9BHPw
1gCjqKf/kVe2I2F2/kYSMcI+XGblVQH1o7Mx44UALn6kiy56oHvuJbOQNSbw2ZKBFmQJIGcHxli4
hmikR/mIRC3MqxcykdQSVOoIs+A1n2kQ5eG77jZ9u9Wp+mfG/sUkVicY4UTcq2yMhnkjZn2pgeeF
ijG34ynYOvA87QGwtcRf8WtEQdtfxArW7zcL5amooXj90of7Za8QrOLis+HbHYgIclDV2TfnmZUA
GRay8w96vILB5+TVplfUhwjlp+vX9Pc5v6AnGVpZIuWUEapUPOhyGGSjz+R8MIKNV4zpy/MDTWEk
KBOEA6MOFivOahf2+vxCiiJlUauTDR94gylArixJ2ZSAKPo58FfmtMd1a+DhyBuK77zB+YbU0W//
0WsA4zZ3kJ9SjZFujMu7DvZTZzbH0w4kaYygcwIEXe4/TDfzt+dD7Urd2WzpLHLVU6PJm5rvHvBK
CDzjDdkZW3gTa4ToPv+aCTN+s/OOJDBrH1GKGlqwQ526MWMxxIYizyqwbbIa3FCYxtUlFSm1GCV3
e95adrnFNSkfym1s4kbl2iaflTKH4ezVm5yhGUdWzR0a70uKOY+44KD/Qb6HrP17fba1j9nUE/Wx
MHX/IAQsWqw5pCgnIIZhCFYa5E+uhIeUhpxu0B2bbajsE8Ezcl3M7uXby7s+WuqqHMiz4V2Eolvr
3KdcQg0B57KasHVLLbG+0SFt6XjQ9KqXbgPIGpovqPHIYP7UczEPHBZi6NSHWJsDvmKCyHAVcTVd
Jr8REh5ZJ2Uc0HMxpM2V4kOicUSKMf/g+7O0Ny4Dh/j3B9qC5jNCfUt6GbO8qaPkBWci3cfGxXpq
jVxHnQV/wXHfAf6pIL3Ums/o+6mJBWiLcGC9S4VB8x0N5KplmzMVpdvshyw7Z8ubPsP637y2k2WL
iLpBI0wr7XATs2hLo6+vL1OJFkVO/gnSqtemiOFoFlPBMhTq7jp0599f8i/TPQ63M7srTBpC09ie
rgQDR2wNPqWQDL4IjYBv/yuGm+Nu5/vI230fMUtLsDv3eFriKdw9zJnphuUduysa3mEOMjrXnKnS
hgmc8SWYV4faSPhsOC74EI8LI/UNV2rsCxJIHOputYFX1CMbf+rxYs4rIE1Qf+J9BVbJnR+CZPXl
5xN/y0Zt45rgtuRaVKtaX3rPoI9cx7tnvS5dQGZDxxG4KvMBEdiQ4LcEbiEVO+N9CSzcox7IsesE
qPo7C6K32j/4WvshDCBODSDnnFHi/ZznbL4L6ordW7uBmloMsO+ZOt7JN7+l2nZ/aNcjRIcY70sN
o0TX3ksPFgYyHd26oxlTAHvpePLja8N83CMYRx4V3cADp3dS4UzOVtVEHXnKNApqdYnq7JTD5K68
Cfjq5h1RnF8KIDQYCcrEvw7fdnEDkP1qVOVlppIOUjQFtKSMdT7LPkwaZYHgZGM5K2NLEPldR5wK
EubTLRZKBhbAdHG/6To9ho93VoMp6ldeDbG49p18DGki5dSNdGrKQcEy+1GLiHlLw0c2KstKHMJF
6wrp2Z9Eh70XEOxWXGLOZa7NqopgwY3YLyk+OxoW/lQ0c97yQIpxl6HftKaa2u9XAtciNXJIAtjV
abbF7Kan81pE3KYIxWc+KmjeW4BaAGryyuwK14JY+wPlPimwD9bThGj4Zu2gjxPsKbieLwAcq0cH
GCXkJVjad8lbNJsIFFEmLRIh1Ez5+z20nzZMDwllrl22lwsqaUelC4JkQA/xSHPdxGphtSuAfR9M
xbZTYywmpfh+ML7qAvu4Gbl5bZciDxH6sF2/cppooj7THKiQbHYb9ewKqtu11UtCnTwGkhEfLubi
IgiSsOXbilTqQ1pXbnBQQ50SD2h5k1WO79qz/sJRdRmc4GbbquuW8WlMgR/qqfvUlKcFBFoLbdt4
9Af7x3nT8jO8knDG3LtdCym9LSdgoxLhYrEN2w3cYLADsvd3Fxtv13Rifr73+ED6txCndkU0UqvF
Qa9tAaplYsBNdPiAqQL2o9X5PzemaaeHcasidIESqt5X0t/ygTvjpEF5R9GkZjSNm0zPVMRkDX+G
RnVlHkqnJtTQ0nQNXo1zel8x/YW9i0G+FdUEykvXdYHz8hjGSA44BY7bSwLGI46mHyvJ64khYj5w
Og78ve4QBIr8MNipYuon8pzO/Cj1vtikpi4zVm8PluXTh32qDUfSI8+wrcX9/heHAlnEDnH0D8K6
2C4wj4hnUkAEl2hrcqBrZltkrjHdMwfQ+tOl5lg+MUWMs27ojd+BM2AJdNPHWqLj8DEr2r0DryxO
DykWKG156FL69oxj7Fl3QUcJRCB5Xn7qpvnPDEPvXPZNoJ7l1q6aJfepj+UR8BDIQXH3vAgThAcU
xM1wuVntxGc0VlykVCqtF+gG8tW6y+iVkHpDA8B6G3pVofy4fUNdSW+mBpMiTjq0c/ecDnNXrQdY
pE4QUe4xgqjo/smuBucHUPeUGFqBCfrdlUkosYxwEvDYw2xecL0VTPdAuwP9yeVHK7hq/oNqU5ML
n/QJsMmZdcePAt5XvbG42WHVY//kvaGn0mYG3FZq/Qt8LBkCOyCxx6hG2Li7AT7rE/6K/DbclvmI
848xlNUhfFbJMAZg3fnlg1Cq3I24Ox8NA4JXFNaT83Jm1NBp6cFSGxHayc/tY9/Rvvcqw1O6prKH
QRV35iIYsVqGti+4XWhsT9vFswlwEL/QhF2c1Q9msNnLEFyg6wX2ARcwhlO7KUKQvh1uU5YpmQEj
It0xqMvKeToWbHil9nEiz1/l8nv7vheqw2CI4L4OGKhULdHa/7F1UE9RDEpDKLgz2IbZhMMGCBI3
BGNWzEXX7ahD+9RC/Cm1r6GD0uO6NabKzdgxR3nxrC4wwQrUqJCATvKiZaci4PC5RdoE11weh5uI
imoArk8B0pD5DX/Zto+x0GZ0J8FM4qs0ZNGtwr7luA6isVWjqVMF7jOTZFK1m0EsLmSFO+fpQcNx
nDFDV3ZK90aZEWS33wHIE2xJAtQ2acp7fptYtcZMqvyMYdh3q1w5UktMbRUZ6BHD1Lkdktjtw720
xkSBSO6QqOpwZgVYM/11cDom9L9PNxAQDQ7lZdGaUP9KqAIUEzeF54bD3k0VQTtVRnefyQCVR5BM
sLEqCeUCAc5t6ZCS+ecb2GmIIyDW+I2Dpog+AoPf++61EjTf8A6qvYZALk4EM4PDbYc4+aJjsV97
Ea1NQmuDvAhmc2hUKwpDa4WLAJvEh8Qve22XeLvWZWnDkglp3ZLV7ngSv3OoLpEkL/8EJObfskY+
uvb7xSjiAXJWWxucy03oEFiveN5X1gQR+7gtIYqYUJKNZEXJqUbOxKfoPAaNfCsLSmd2o+zHco2x
Yef9DogoPcmfZdiIkUm7JvimB7bLIM4KXfQdr5DyIIBJqKfSqzwns3colOa2sq3XHCrBtcSJiQNr
4Wr0HJoz1JCvMvs9qBcb88fJW5a19s+VK6F5tX9xMk+NAkp8c70+zOw5VObQ2eDk87jee8fpN8Pq
4bUrODFBmnNxeMsTv4+vSNpgcR0w9WH9KdXJptFukt4v2nrurZyIb1hwpqTPLv/A2JxAs2eO3EDk
ogkBhp7nOgHotcVE+TpUBytg1gOauwWfoWOpgVhepDSfrd/g6H8zPiYMkNg7exDa31EmQt/XWI4Y
7XeKJ5PbIJ4i5QHOJFrFUrFTWhA7+9lqJiwtKAXORNb1FWv3bY54S+CfGMySmqZVpVs1nwQTLBWk
CB9xDGsRLw0k3mxyvimExJQxKC2OouknQ6OCxkQJCE1ZcT8xaWEaigAfNE5gH7vuFWBcQNfWAstx
oQuakn/wxoIVWZa30r1jkUxyh0R/JC3wKSkkwlvCzMaCx7XYNkZEkVljqjTw2/nY2QX4WCsURAMo
0omgzCjEmyDrTbk+eg0FmnFA9iv6iR9AwEOMvvolq0A4i7wvINzReXa7ocpPckECyD+JiSEHOuKl
glnbUKmz7u6uSBmztun4BNaGfamUrtar5Wg7OdGYI2BGK9yvGR6El9Xb0Wm7lkpxVFx/q8ImUYAu
7LZCUrvTJfSWSk5C8VObAerdO7E/M8tAZIfApX7jG1B/E05Mamp7ew6Z8O1MQIDy9aqleoQAXapT
wBqXER6ZBygMMA2Xw6c0MDG8qrN+Qa9R8z9UvNG//c+AZuIpx1IY6rPhLDUId42OCK/2L0Uk3+2D
rGEaFqf5nGCMreKFMCBbasJxedh1QarFeiWJTM8FLkxTeIfS1NXMa/Lq/I0sdsepB6OO0Th3WwEy
amYqVb6hUXHTIpET0u22af8RUNncRPWT96zd+cwpyal5ZiRMINNb7lwDz3lsyflECY2OKtCD1FeZ
X23RvsNr+0X/oBewDyI5MFEr5vtv73rygrLe8/sSxiJcfZOO9QbVzTaNzThTDyyHjA9UlNc2E/o1
TIr0LqglJrZoXtXTvbvP80C86maMfJMJauyhpDS8LqTyB/zu6VZIL/4A6Sc2ZAsSCubDiHOlJ9j8
gLng7d6wcl32/Pdi+Q+xbW1yDsokjTvCrnR7ioua6zTbSk/kAYdHt0nhH8Ebi3l9PbdMV4MuZ08W
m3MsjbMvp1yeP/9P6m5wLVV3HdhJtiv05hHwrwv3jOaUw7ERz+nQ36LjhaPoLJ6r4RlzQ9rxJu+P
28H+MUL/j1C3cgZke1asVLt5kG+EiCSiNQftdNzQD1MQo2qd3JIcnNJ1feU7KldjLDV3EfYRqvyI
xtl+esC0ZtddjSdDCa+wEiJnWh4gDMIJ/6LfyR+VuM4cUfRJlpj6IN+daW0iTUz+t+CewX4ENEGu
Ge9xvIBr6SKmY0rtGQbO5HM8SvmHqkypTUsPl7XjGJI+2REuVZMBrIELWtaiEqeVdPggxATqbpQJ
x5kRadBjhARg1Y8ilMWtQ47ns08H+FKB875BDSavFeccFM0Z7vt9vQanmrKMY1nFmzD0snm6EHR8
D5zNQDJK8tHQzWMtpX6ytv02YHSwRY34lN9xsO+QH+8olLJHZHQLQUqCYHyTy0CG3tqBLD5GP+Up
1eXyT64h6b/U1aHWJenx+1pzdarJJeXPkV8fbTfA1riYwtc5YTGX1vU0l9m2pP51J1gTy4lIkFcd
XNgKNfn6HJ9JQVj08ZAT24z1ly5p8K9/bmmoX8CfgosD/z+JZ/59j/XNgPrTg3zIfz3l8RxwBIHp
Cpi+ebx+WbFqww74KwqVPr36mlcdUqesv1pvZvgFhasR6bFYVNv6bZA4H113+tRHuiUhrUtSvABL
OiWGNaiIlQol991TFjkAikP3SgQeirx9fzSao9F1rrf6DAhbFnuaag7CcWXcDQziQ/9ieyuA6pAp
WIB+BQ6XL9hycgffcpNCa3N8NG+iPyOBQdjGQyucEysczzTQYVu9BiH376KfQH7djEVS1DoanP2y
dUg6vKZVx8QM6V74jK0JKx5lGsXNyPJWKpxozIwLHwBLobPiIxwT4gdHhWbHT0TV1a5swchGn0y0
g6XDLkbRewHj0ljx7VCJz9itLL5ZD+4noPnDHUOMBTYhsNVoTunXETS6gG/L/dHcNqUGbQh80Cf+
Z3VwKYfhbZoL74aLNpd7scpAwa3YCckSTKolpn7zUgGzmgaMfUFAd89MRKkimTm4nl61PLRlMBht
1J7ZT/zT753vPd3T7E97Us5fle40+9weZCqrRxqS1tf1UHelmwMel2jYhbS8rOAgTNCAGd+zi4Rc
GlUZQSxcmJ8JoJ2f53lQCvr7M7GjoE31PpM4ddI3Pc58RsCnvBmb20r22d6CEDBbOOF8my1h99nw
fudlKmmaD7pikJ9HDgNCEVhKIA993vsyZi9+WGeAfklNb+nEDp8rCiS1FxzcCtjdUhuxsQVoCx0x
obGp/vPbw0wumYfVNOJks7dwwEZcTUkMlu1XgRAjg8eS/8EHmw/JevY6x6GZks+RhT4ZCm1zfkw9
wtzOXgGdUbb69pbJ7QdgSWv/fGT/9VwtJyPyhpemUW9uZbxm0roRgGhwjkCHvbbPDZMQ6qJx6ZlC
nC1xSwvA5t6EtyRIsGrsZfp48d2uXNLC6VpoB60/g4JKaVFD/o5UBH2lktsTvEUDgYqFQB5m/1Wj
Gm2tLW1vkrmg2rlwRPDN8meIPlAMauvIYXbGc2iz1oCS9Q5RvB/E2f0D70LjymDa6qO7glxBTJuc
f8YVoVnSpUPzzn1ZAMTaf4QVycp89eq5eHj2Ca4E/bv95gGBmGz4F2JgpiGU6Ym3v+JUKjbSeOde
UpRrYO15/e07Id+RSal+oPVQ2QiyOehdFjP/YY09wZ1SdaYSsJejC7RbkqlRHbRoT2T/IwfBaQyx
XODwcjoP9aG4MctZIKYEVAwNTQgnPv9iCS9VENLP7Nar/k/EtvyzjlG5gGAadcTmYTmqtOVCj/GO
o4m3WB4g/btaVg8w3NtqB1LhL0SOSrHKHN8z93s0vSe+0V1TeYohtXK2iO//6s0HMnl5+FsAHAFI
xAIZoAvz1bP9vqF+C9oCHTFqVMR1l/PfV8JvzxvlZ3EiY5Qkc65oVtVrs7VDe/67xBL2y56PhUGf
tmOPmuAfznqytQ0FnDMNNET7KEBQ2h0WIR27r9BeA5pClTcHLl/uXONpqp+dYxaP2un6G6NmvCTO
rDxzOk2Nz57SAFL5o3u4B04IDq/hJC/lNkQ7rnxfE7Gv8kH8+T7ADbmIZ7Yq99VtW5eRRf0r4qH8
IhlLDaFYk6aENJ7Ax1uL5TsgawFOLiRtLqs3O45/6CQ57SCWw1GxxSHF8aWnCJPcDyVVhScbwpNx
KviDqEDmV+jkKD30i6s9AkNoLSwoC0klHTchbUqYM3k5QDH1r2TFUY2i2u1VCMZtiYdYpMBnOwir
7KQU3Ysk+Y6S6ucnopiXzsQUkSl02kX/qHclNe8X//A6g9143/p3SQ9js5BDz3BmJRhEfVGk48BD
J/PAt5LvRHmmLWkeygiDbqv+1bC1vumDQARzhZtRNSYcYnXxPmuztu0M8ZLTWU6GWVHVpdmOmo+9
ErW21gsfjMwBwUZMBgLc8CvGIvgJNzyAgaKwqf8ifRkKGnGMLxw/GRjcCP0xgGlGbY1ZWTQc27Cx
XJ7cwTU/okWlEMi82uKvBScersfpZNL0b7I4WVbibFpr4MMCBCXGMx4p9/Ec9kTucv6KSXS3ObH4
KfQ64GpFtT1XtTksiKmvxdKq/qcN2TEvztDOpwNExN+4uq3j73S0O3U7RtV4mulTa5NkeLXZmF7b
3HY/2MKsV6eS3USYkZKFeDLc0gVlyKT1ZffeoYuRcdR5wBFeYjbFm8CW5byeJjxXgAowHkEPFHmY
5h78YB3S2rawGFMTupnQaw1lggnPA8waPBCC556EgRymmK+RKYprH3x0Iw9kzaXgTOhAeVyf3ZBW
CxgUQQrhN0y1O5ECtrcJONORSfSc/bbE1eEgk7xZn5N7K/5iK+53FbR8cZTkVm4KhBGonkZhUrll
tGdkJ6JFPwGtfvBHZGkp8gOOovbpk1XUswNAuExB+eHCnjTBaDwHhJxqAbDbCk8jywYh3UliP3CH
AgRYMG1N/HGLx68T+pHW/QeC055VmWbZJccHFjxGGad4v5fFvCbqaf3IhNc5YyWw3o/8p8F3nR3d
xPVlngMsGKRwPGTRO5+H6BaHKXrRyCzJRMVDriTtjaTebWMgUgHAVzrF0ZBBPkJsDdRh1AvQjDE1
BD8GyJUDAmZl9nlRm0Zwza/wgsuP21pyA/MA2co6ltDxa0bimLVcMYtVu4AiMHbYDNrz26/xPlv7
xHyWUqAglGa1HnRXKn48jUFmj5MA/fj6jMYift2nPxlwpekQLcQ4rhPA71X33IyHibd3YwvAujGI
KybwgNPjF15ayzdBYbnpNfmGVLPjYGg3UBecb6Qegg2EPIoOm0py3LGgDLnedJswA+f6/qrMaitl
ysZh1oEAWLFqttFB7PcRKHYouUUd1CAEervSXivUdWtKOZ0vts+xyJXBb56pEmoKoBO7QVtKN7Mn
hAKdHkhZN4EjexJKRSPVieYzi7h/VyL7RDS4+fHR/f0HFxQ3e7RBhQ/r5aCAqB/BQVcft6W+IGF3
Pgxjp36bDnSilTM6MaYW8GvfEindreq73eDGx8bsV7ZyKgn4VKCENg3+UuAyUao0E2L+VVdoOeDJ
wLBZNhnKRsT68E1AEL7i9XI7PO7U/suxzQgM7uN1WQEVp+VCx6mUrObLLYkyxKS52vzc4TQoXKZA
AUNkxEbgGQKxQoovxC3ViiNbtdws1mIm94oBBNgkVEdBDDJRJJVU7q5fhSZWUNzvMNoI6y39apsW
3z9iXxvCp7BFunigFP4g6Sfs7naUKRD5IOSR3dVXeohwJsFTafjrgtthzCz5fkGTy8rQriAbbDXM
R6PkFfmfFki2s9V6W2kzP7i53QnQ+Tmjz8x7ZS+UvXdRwAJv1MQe05sazX187Yg/IDdB/hoMiZAW
7slUp58pjKTkFqfTb5moLOYO2o904W4BbGl9uD78J61+EKg0Bupew7ry0c8ZVQ68nNqfmt/Yn0C2
rqJfnrPPMIRjmYb9PqiPoOEQlPTJIQXmDdtpdxjj3F7EAQzSwDqWN5gHidgJT+XLl28mq1kI7Ra7
pbfB7z8dfMWYjxJnHGdD9C35AM3rpBXHv4G+4pfvQml0k0Ji1RUjYBA5OWNfV9h0M+beB3zP5FPc
x0xSzqcFFAsQ936fXJCqfa27p1kHHEqkbt87XuLsvSlbxpM7R2mjhNMaz7J7zcxnyFbIvIREVSYi
d3odDUt1zTAqHDGHuUUSLXWjpy3D/tEN04Yem448LDqjd0b3oNzbWfApMQ+WdUM34nHqj+elE4uJ
7ttvKN0vilBbZA+SrYmerGNNB71GUHUBmiB0lG7ZHEVx4vZpeTNvcAYKlBarGUdaAQKTF4JLFrCW
cDXzNztqPz2n2z0VXhXbOpMniaenWxzz0hzyuh/QEW7Rb1gRVZc8PD6syes0sitYEDDjDa7elZht
E/GT8s0wSRA3OyrG6ZfN+a8cabd3nK/dQpYyF2WyrpmlQqeIZcx60w5Oe+mH6dE5oeg4Nzq6OxPt
cX0hpcOkPHjHMB/EqEPDz/7G2FU7Z/lDo9SSE1Ico2YIMohBZ+3P9MitKkFcvvZQ+l/46fhpIPUy
cpc+Ae27CD3b1cU4G1Ut/8KuoJZC1regohhy8Vk9d6kTXXVeX2bsIMV/1tsoTNRTz2Lu6aoKCGe4
hKfuL2nXgJ9sB99WkM7pBw+ZCplsR2H8z+XRMcKUb2R2bNR2Lpsc8/MenlQNLjWAz/q8lilk9P+t
zmnlEtbLvDIFqQczwuqq4zGvL2tI4meimomkU8Lb3xzDRkaf37SZX6vxpu8S3G5L1PaWqCz4Px0S
6PWjOO3mhd++IcYGaOaUTX92GFukIZbY4bikkCZOL9Ib6F2QIh5gM0NIZuaXVAQHnRh0Xjl/lzd2
Jb7nty/X2dXR0Gqo42j9Mzp7cgZE2oI+Rz2Addv5JoJNyBC8whIFQjMiljXjdFhCZ/zZ59OFVrR3
X9MEezSNOwmb0EyXRzEYyz65vMj6w1+lZvoCSxR9MKbQU37ZXYjHPkI881gIJgpFTMRbMgnFC78X
BJGZDlvd6RjzT+u59/AR9T2HeMauYex7fpUlwnnfyRdSi/uv0eTs7LWLLQYyfVf3aUSiVth2/pF9
8QcBonPbeWbB0Z38+FevmWmTUc0+CRkmMBCb+ai0HnZqCeGlDsI8HTG8UVoutpIx47DhIyxmLgbS
hLZ1f1WWDToaiVkllKoiB3sRuIeIUtZvkxprtTXXE2Bx+8STGQV8g/nYZGXgcg0rRVREUySBcskw
xPkvowwgS4JNVG81mmKmzzOqoYITyQgCmJoqp4lNbQByOo4Uu1b8VZA6DXEljspV2JdccAcRX6cQ
j+waqF27YXkv2HOrooO5hxgzM3SYpAp5TjPQr+v8LGf6G1Y5Dw8iSOM71LOs/U3huNADRKQz+lyI
PLehGZxBhB6GYGssFMFL6uuoH/Lr0IrrJn8WKOLqhpcE+qoxKFY/iB4IOdtv3VYp2Kpzr7cFeXoW
tmVEuypfCogpDcByRAGMvk1WIw99WAk0ppTmHOGVLhx/+SEbGuiS3Y52OtMmQ9ulmC3hLrcOMmKm
GTB+Nx/B9d8TtQNe7GvUY9vDjTNwXeXxMU/FLKKuw3P2GM9UntEYIk8nm79X/CAtRWJopMSOmz+l
NQeBb/qTWPBBNTgX56PBn3OnXpTwuGhjoODuUlnLQyaU/1xTp5wx1dnfqnTMI9Vk0MCcf0F0BQhT
EYwtdKt0gFvgISWCNfQmRAhok3JRdGWnhc+0Kt1vV5VqNwLgzwBtV1JdMhkuyQs3ev0hrud04jgK
n80JFha5Agb9LeTu9/PlD8rdpw65tJjjzs2d/suu4QSmPYiaaOeBVFlTNmu0by15WPX4IX8tdSlo
KyqQBOqOC98ApQnp5Ej3UF1CCMjMTzSMqTErk9B0cw32eMjRwZBRlID1M4CUBqleMQ8emVxyI2zq
/GSs7JqVAndZxxY8XEHZoJs7V50C/k+RwULSyQ5vnQvcNwbqUVSNfgaX8MrUOKFudUEEjFDjYKwA
SFzRIIHgLFpSv6nkQQV/669ol9rOUF0aNYystactgfrjMvdpj6NSjsofNoJ+iK9gO++b6vp74iC3
nqp4q18Rjtzi7lK0eK5pb6bKuI8KYgJoevhmAmYGQ2TOneDidLVvYDRFFvVHCazmIT6SVzBk8pXC
PLW+YL2Pvrof5+7CDH6lLktSCLdlf6WXQkoD1Jq6xO3KXtwlOyBK5LRxDMPsY76k6G2kTBfnTM7Y
hlR6cI16xQBpJMf6eLpHK/EE8xpDKoePU13luacnf58I3RPwrJz1y0vH/5+W47v+W02CSmt6CA2G
Cg4VSLe6ofb5M6Eu4CTna/x+XUULtyw5tDXQ2RUu3DQVh98poyHZZNnGzMli510Kmmmbc36HgBdo
vQBmRmos8p7UvFkQiRPyDYQoLk1XjkFYGsvcNf8IgvBUZuF9Z8c1e4OcBYMNDDMtsGmvcXJM0bcc
OcSTFSKF/9QzyBRRzGU6zu/kLymn09wyrv8SJCRHdTb02ZP+GEaPbaOiB9bj7NHXRrAF7tJ3OEtL
s3H8t3zc4VZ1quvD64teUu7vzTYgcOh5u4mJlgv0X07Xv8WQ6AdsjtA2+86cG2rzAiJeytGOYo+v
xZlGoXgLy9HNsl7YD+m3X3fGMMlSm2bcWqQsGq1NRXHE+Nhb/bshav4bsVgnR8dBx3aALqvGj3Ae
u9WeyjCBe5oHlL5kIqlkO3i+T1n+dBB2AIgYkMKmybrdR8EeWmCFZGhOmTp48Tip0hhMX9HCxSBv
4zQK0CRch1/wJNsO6xD8Tpn5pSiKqqBxUMQkI0kkO1LsKNpnJdL3SyXSbGq2NUtSybG4JdbbgK/f
2XJJruZlcgmTm+BpFbedd0ONiax5GOT6UFxW9lxdP1ekseXUbT0CzIvcUxrI1HsYNKubyfSkeyme
O55zevAxHFCM/wxgkMjSz1gZSNe4fBgbIto73tvZafgWYdEcTd7MwYBt+0peGgsyKZlJXeSbPN2v
lvoHKbGG0xgttmhzhYmTNCOtuslxV0u7G4TJmebsat9L5jENbQYM2OojgdtI3k8JmWVeY876STDR
Kb+poev/iLvAQOYsD2o6KzlHFc7o3NJ0yEJGGPTvTxNt0U0JFEN/wdwuIeUv24A0ibrHx/ZTyXMI
dVLWexO/EKBmw6WRFwydPm+tkG6ViJl7EL9qWX1vR5shGSpv/fOkCVQ72UuW1Nxif4wAQbt5Ph9C
sPw3QdSZQchkyOcUmsg5aajdyMd74Kag4lf8EVH9AMPQ1LfGgqhdH2VMvU1N7iKEhFc2iCJPxdTI
QCkPUNN1D58aGeF/aOtvmgGaI+6l+2q1AQapst+DJDW/+alNMUbdzy8Dg/sGKeCJY6yumJPbFJe0
6IXKc789bRVh+3cGTOBAHAfdRpjrUze1JadyUyB8yrJxrd37DuxS0Bud68RYabahpOvSqQ6MDHJb
OSrfddYNfgr0Uggr/QYYYE/GiqotAX6Zr2zcC6vJtOuf0hZHpb3bV+K96GzSmaNXWiL5AJeWrna8
Ko4ZMmsROymRV2Bw3nh3GYEAUHE4wFoJIFSTIdHsBIP98Icto4StqPYpMAX90hkCvB64uNvk9ySW
ro2WxOEjtiAxSjyHPJWsR484KyLigx8qNqJD0FQFFnKkbxjiotYbuSUtOjYMN431+QHDEsdkm/Id
cYz1KSp0iB4BTxa9FjlMDEdweHARjS4m5RhKlmkEY8+5qta7FrL2TWYGercavjLU77hrqlJfpMLX
K7+4mTF2BnEdoAZnyU7ROoLYjJidFbTXuS+P4bmWwqqdGcQzKj93/Cs0zVMNr+YyoEmuSpjNYfyx
KVRaZJQZvs5hEzNj5sydDcJ6eOlabv6J+eqqEWVGp/r5OvATiHnsb9RdkLyhBS9XAXB121ZP0njr
mht3Vzf7k16Hs0VrGUAFTInoDin4AZij//fm9vgvV/JHpMUAHuqcrHxVmoh4/nVqyGEU4ib8DvF9
tzbtvQ9U04Nap8oxTDUIiztqqreab1viHH++tBLH+TttfNV3ZShlqtzGkkGqRGbNYnfgtlyvPaYE
isVO32KsK5ej7L8LWOUX7ML8qaG6zH3ueYQYaY3LZyYJab9uoxi1TZfS3eeU+WO1XCnOGoiAFFAu
ExiMwWMGpOYWhanhu0ZoHrBYxaqv6ABKtROtkLkS9yDUiUumPOfCOo0qcT2Z4oZ7HF8VepPHWNmb
L0CEUFRQad2a8Zr5YUFnJNeWmZwbTz8do/k6Iano3lrJU6hUXUUfHIg+sjLOMgJ9/yWnYOfO/U2j
PYvzYmWU00Y5L4wCIlM+Hj6qGFwmsziGuj4+7UTf2qykMhM1XkjRwszyQXs+KGF8FhjXj9xp1EKI
lwjPNl/FVCDup91osVvNBzJr9kwGqVKPBUxxxhQKsImh/CyTC3xcluanPPqs97CnOJpVpivrj2tK
F8eGF1O8nwyVVvxe8Z2dSyqgXsYGEdVvq+qwfjkvZFdsAIE1cKpTXZiy8Ks6EKtF99ztFu1nOzCY
jpQta2OQfF8LR35B8ZZydd18jJHbanmF1pcgv+gY+7sZesQeeMMtxDU9zFRFW1+4z2tFgMjase/W
Ufn60g5Dn+oK5YPEe3r6JoYIdV0AY4kJIoVUMSfc55Esv4yNkMa2fp87Xdd56+YpOsFIS8syVFmP
pBIvT8/ts88a27RP+v6IuX0jhCm8l8wMtm0laKMH61OJjZK0j+3ypV208sKNFK51VmCDWRBo+v+l
GcaDxHbMK8BUn545TFOdmi7Qv9PZomMTwL0OuIjREeLMkG0/gRwNkIlSVt8R7pX09MIcbsonz3BH
CayOc24GEVdo4L/IyD7lL2DD7UZ4qX7JDywirucHFkw3bHmtmZfl65bdq8ZzrBVYyRJ1/wtdNlQD
0lETRXDS+S9znREZNm0+5yimOgKv6x47QfZ3jYFk7AiBIpf8iRaCcyyv6C6pT+Zf4ZYGN/2vH9DQ
CdE7mCTdV0kFJTIOtABAfpSb4rxdl0Ee0P2J3h3h5LkxRS+AMH3XGGm9iRRajDIKJu7jGvfgCY6s
gnKnoAFoOAg8XZCgL5sQehpm6FWwYFGIRB4Ky/eQOakd9844TyVM8nJ+Kiwk5S2gaxC74C2OMnW6
B5+QZ6JY+tGBH5XWHDsgcR5rFoMpd0zLyj6aikiIcOMBgCInvX2Th1Q3YLbQDqaW+E8zqQGlE8ZC
PGyPV+ejedc7TbLzC2xvFaEN1kbXmnxPEk9TSCgFfczchHNaXJ3zajIC9TBloO5Kzf6C8M1/kIGr
z8Zt2VF5vbtpGYazu11cd2/8JRiPsSY5VuDGEPm0nrNBBmZbx3VersOb3tM4zZ4eH8Tj4IJsiDYu
mRJcAKIfQrU2Ryezsf2Qhh23KonrDmM/JrBWDzkdXEgdrbbnKo0itntIlvg151ZeXo4cbmizpw4a
+O/EhZYjJsXh2M5nb+ixRdD/yHS5oBwhpUxsw7fg2xxvXRwFv1/M90v9/hf9cJ2HT7ugnOuZbIzW
1GotrFll9pwLEwiRoLewm2uOenHmgFw4FdWHpMH0kSxzrw1a87hQBvAtbmmyFC8VA7xVuuKdpUXv
ff3k/2CKY3aJ07pYsn/KtvhzG8HiALqCTf0AjBAMqcuAyH5U95fhCNSmdtaPCDqlv1EUovpyspk7
xLLLMIfoZJAMdKG4ekD8HEKpM9kfWUNj1Dow134J9WUaqFVEaAUJKHmB8YfdZSG6K0xAsJlDEzoq
U7+rjx11a7IyECaMRIgEjStk+2VWXe1EcWyv8007I7KYNcSpbvKmVVOxagidca7eK2jQ0TGno/tg
ECXvhrbxGDvtKYoNLBrx/OFPNhPSD8n0cDiFQ0q4WJHdL6hnOaqjW4zDMmoMu0mfEseElloeaPdi
ZHs+TEoaPszhbayA5NNrr4V7Jvn3DCCb2v/wZy2GkvBKrtLwthfUPV/mAqJ3TaWUjhp3CBxAbW2x
IVu9N998EUo8y+P8P1FvR+KV8Vau2Cp3cwAuzSDLXAkZjoCnFd3hefrTxBvMojFn4/YZ5YAdaeSr
WL/mgly9jjrfj3dtmVs5l+cojP2fjx6AqvrmXuU3CKzTZrie1GDXiVwkEkzUbHmxObH7yxwCWaOa
e7RY2RuJLp1PcM9+YsE7cypXR9UMfJ8KceY4NNOa8Pw1y4dJCm3QfYKunPJS9THtxqvbK/6kSSl9
0l6+qqDGuvevY7GwzPxwSqjcbo9ze4eU3RCmfaI38YAgj21ScGpa60bpsuH8oj9lOMDfpmvqPeuj
EWYH0Yvq86caNIfjF2lMA6Ff8SQ7yLc5bS081MkiZkEQLIaTUsjR456ozrQ6H9AB29KIh+kg6UVA
0PhSVR4Rt7CIDC83yvh4mms2V8LG/5D6g3adBIzaN0XHydQPxY4AobcJNo127NEPRDIutX0hCwXi
+AkM9Ghwo7QKN453bBs/FqUPuxvlSQnF9RKo/BK7Dq7WkLTRDIRtLxXKEuifdajNOzCjPOEjlfNj
P8zTFRW+dABf/HyumHstW/0owuzyhPiACrf2Zh9OUUOTX37wgMLytOCyQAQZnj4Gteumbo6WHHzy
bEromtPYjo9Zo7jFJ7PbOKEFeKyHODfnG3po/tU6DE0eTKpYsCJKp1LxjpGeC4uF0SMj3XOWfaPw
uzwRWUPD3DoFZiwh2plaXDr6uDNGnG3bjtfAhXgtctjT6FxRAB5E0eF5Aore5CpLnfVyXnUq1AUQ
KpKFSrFhSRw1aJAm3icHCbXv0GPK9C9JuFsuHUroqBV2NlFUY1/Q7yTGaUJoyAX461oQyTh0o02P
SC3qQ9g1IhoJRU8NxsDGZ+Cruj3l3IiLEc/cREYAfamZcIk0IUNNP6l9G2YK0Uy6VHCse0zTYnIW
vbEwNX8bQ/KRiQnWvcZBZgt8cnTOcrckaILuCJU+jluK7jejLy1vDAXt0HIj4o6mXLtfCJfA6PDX
+nEmklHPsCLnvu7qh4FUybsbPBqRwYq1b7bnJEWAvRFBeJEFL6f6SnOM27Erqtb/HVxETbVUBZ9M
zrjdlih+jxRNj0aHQS/yI+8P4ussM0RxZSoZQm5jdQENtiQSFzReEME50zSH09X49lRNdWBv/DFt
JUUfaRZnCGfObDPV0vqQ2b9KgqpYFhuLflwGF8iZ22iutypVDmMqJH7zwNGKHruJNbx3osDA1nkg
qQMxCmJEvAJSgR9YSGgKujuCVPvTme80pgIi0pjLL7Mp+I2X/8ePf3gKZcvPMcNI9/4N5Ws223IS
uFAbN1kWVkpzPmBYHw1qLPFYNDzUCXo4WwAooH5ggGGhbHVS2mPkCGBOO5QF4OPd1IXQkuIimHXi
8W/xg+4jM/ZXOjGU0DWhHnMc15ZupoQp74hvuXyLekP5kqOvbGIhBfbq9KgXOcIPviy8H2eTgFA1
IadTEYEddVZ9Quwe4YR3QUVg9WKIe+JnWbIStZg9n+Rw4UBdYubrwl88rJqzLc3ugyTx1A/sd5+G
nrt6b+RN4HMnE9z4/xmNiXa32XE/p6hFVBOWKVAvYvy1AuuHTZK3LKTFwc+1D/5WZ9aDUbuxFmlf
ajlycJwLUO/7tDbZMUL699RkDuH8lFNTWbJJP1QlDxs/pveuT8jIlDTZrpsZTqsYG8cC7nF0oqoO
diWRz8qRpsiRe0jZMRJn4R9RxR42WVjiW+qFea8g2p3ABAhnRFN9j106fsz5exJtd6Vvq8EMi61y
DtKQxyavC9Sj5LbU5KmHHzNuGxKTF9VoHo2P4NHuN3uDtcgEQv3yoR6DTJUMV83/teK7E+MJi5Dm
SpTw6GejUxSAnXHJOtfjrh4oFi4Bylj8Lt2wq8+gEws8TXJH5eVZj4wXmzNb3AZ0+IyTtnJixdTv
ZHeKT0L3FtZRdffxxjy1wWxxRXd1Y3TDgU3zO/pZ+4XVz1K2MLjtVkrWLLGcAWso3p5baSHfOJk+
dygkURfGLo+8FkT24sB3JDN79/h/JLPl4/+LtHv0MRhMQ5k7cR+6qh1chhnZbUx5kTRVopEDMbzA
CVuCIPtvyIwzOWaHXVN71lgvRvnkBqbRYoD+Tl3VdTjaI996NlWH5zzpDkQMsk/JQHOGBeEscv1E
hlpccCRdB9GZ8iY3uNX1Sh2FEO5xR5qktOrw+nQKoAi6sE1r8c6ZGhRMt6b+m7cHUETBoL9+3Udm
N5zspzdPwC2MQ4PSzRaBCwtm6ZskR2FXoHwmfAIridp8GP2BHd6wPqMLci5v2SZZ9C3w0iZ1wxij
DqvUETWc1RczKynEWbmM4sZ7YDUlVRfDI61GJ/QqlMbX78Ro4khSGA5N/zSWFyX40i6CiSjVHH32
KSyG0oi4czZCwWrdvb34763IaSoh85oWuWuaYj9T5VpCj5Gam8oZZDR3Pv7q5J5bNg/It9dnys8Y
1TBmAfPrJ6Mm0hzuCy95S7LuPMr4tEQSYxxmLvlxC2dFbZ6aooMSknTtf3jBeTN9jKYrluLuMuJ5
F/Yx6NjPynjZKjvasG+c4cNxLSJOw4Q/xVlH0Suvp4KhweYHzV28Bic9UFaVrqJ8cf1NA0oaz9Kz
pFDlNSucgyc6QWIap7xJwJGcCKIeDiK+OaMXkCa1hFaHOpJMjBNYMCP9r3nqEHorIIfP9F8mYkuq
HQT747n0/9f8OJyCC+K/o0pHq4oMmpPvlY9wQ7x/Idd+riTXW7ZL7/W+IIMFrmjZpiO14tFzCXnA
C+dAjAWOEFpE+TElctTFGUv+Y3txUnYu6Q0ORra22/1/4fxVVcYu8hgdRrrqcJO7AwCye7DFnmBE
UUkhDndXmP0PqHrRjcF2n1UrnH9z0tM2BKAzseJ/tlU6pmnNR5WHe1oQvvG8c4rVYG24QwbhbLPt
zEiMHO/u3We0PNvldjJ3bWJh/GrCaEVc6ZGXWYLyy+V0ebG1TXQ3TW0tlzfja1S5gzX62q4xXB04
VC6qgLAVG3PMnwTOsOcbZYAR4YTySLTi36FBt+Gn6qtO2GEgksl3iIxm2sYL1y5+n8841nEPf1Cf
vvG+Gw2/eScfnD7V5Zk+qvFEtt5MGz7H/Q6bLACvpIVpBNndPyGRc/dAxdCFUzz6Nf2WKWFKQ09t
DL5TYguPDryYqmqmmyVbfA+hAHmcMGxS73kCpInxi/IODYmn7o/qhL1JXCefABLfUq80dLTRa4vS
Ch0j2uUf4VE9Vh1gTRkRyNr1Wu//K6LCoqMcrYIbDDMu+QwJ33rk5CN8Aglt23d8wifWNjurzPOu
DZbx+6d5eyIR48PvGg8rUbugDcDOnR4kJl6m4Mpn5u8ynX5/T8q+RzGn83JrSoqrbYA6QOmlLWVn
4nBFqllv+dvsUx7pRhKh1vxz06wChKZsQL0k7zzZf4vbh0Rm+cyqISyCsDmwZBHZOMUOcsH7SWRF
s4WTxf6RfJk+vVkLaEb6/oe6FV9BouJ76E256mdEkpeEo296CUGQmLNi/o1TZJfQxFucqPyZ7hN7
412LPxZiPCZ6pFUkuAWmhGx88OGcgeq8CzU5Tli48AdFtEKEK6dZn/qfAp/36fWt1FSum36vakbE
MZSgl9dTZ5cajwdLtqMXa5bqxRM6ngBE8ZA720m/WYUiB0DN4BHvwkXHpCMYIrTNZNMjJaSh6rGp
US7pYP+Bd8OGd9HbTp8uPIyzJS5iRHL+aAPoBQ+bwwqKyEvG0sfilotvzZsRQ17VRk8+n7PtnX8Y
MpXHkf0jSqogI/J/T/mylfkBgZ0f7jxqww3ob7HcR1xytegI7i6C+d3pqKDKUqDCQXfWMjpsByJu
RfVecsJ39CSnnYhP/Aw3B0JWU13SQ7Z/mQ+oNZMHgYieqxTGtQwl3Q923rMOo785tIp27SP01NWl
zFOTkV0fth1beMFEZgnNc4MKLDv8DlXB0ZTv2DjGDxciGOF7oflvQ5Bg+W2wf8O/F671jgnDnkYZ
LSMSGE4yGhqBtlLiWWOx8IKeyGDZ+4Hvtyqi8AKE6ZmdYeSEtclOiikOK8HzB4IPplf2HqdLjcA9
p8h843WL7CDouDN8rNhOxT61dPaU0cONuxt8RaIqchyAN6p/WdPfR3OeYllI65iBzT2pPSgBggoC
RJSy96dbOvS8iA9JaSfoGKGC3pYMunaz1uRDVHNN867BWhyI2a7p5F1ILfByair/Ek9O6Ton9qFD
5HfinHSAieRxgMJCNPnkyRF1tTR8yhDJ2dcZbzG2BWLAJmBQ3Vf7AnFUoQxgN/+CssN6G/t5O8Ko
1UkdsQhVX8VBxTrfbVJ1BR1RGp6o40Iq0xFcQ08TVPe0EaGEESMkg2sVBXC8gtl17QH1fxzSKVxw
095dn0lR27KV9msHxyxqJIriuk2DEAOxqo51Yc3mWrQo6yjnQ1k8DA3Lmh3Uj1UD3Hra2dKr3IRQ
fM+WaIk8e0LvE7SrFv+lIlaKDsiPdyXcp9iN54Mh9sHcdN1HURizA3lNtKD7PbMVRsYUMx4nsP7Z
hj+OsgpEfSVcMP6sOxvIrIY6YyfgprJQPdddh4cNdEMvoTYWg1h2LNUSmgTovnf4SjsMxtIhDRpQ
UJhU7sogymxodUjKiwRHdLPTxOMPYsl+n8LVRCr7vFQ6OFm/8r3TNMx7u66vgMHWTTinO4pE1iad
2I8kd4H8jRErReINVuHWY0Og7d16d7zsJkh0Qpbp3/fgWan82hkX/lFa84lrOiDBn/IU7ev4sGzY
0HxgydAmL+Fa1gSTagMZKR/lLpCPyrj8GycR+Uyu1QgsmvyYcnWTf9WKs35sa7F9thnNLx07Ooyn
FW93G+kxHam0lwvCDFIlEo8PAd2xVRcQZpl9mLbe0QCaJ35e1PoOMeo+ykZPVZyGOr6c+q0GIvxj
XHPO8O3bJTj1bTHwKmx6tqCP7tBI/uUSaZGjUPxEm1cqgiBGGkxgv2Ck3OF/VcmGAS0hFKNqApgX
xAMtQTqSCkGpkaFlKuzAiDKoc5cyFueVjvdO6xZNfcI5ZCXAlszB9FQQjJZgM6IbSMUicVWAPQ3U
bFX7c8uaJ6UR1qGJd7ojeUzD5j6XjnJemELzDJee3824pT4X4xWPrdZDFQe5SDOXKka1UueOY7dY
hzk7xPkrtkYDt0RprDJHNRv6n63avA9GiGS1IdNciCNO0PeiqMrnKEY0cf6FPGhOYNC58iq2w3XF
rPkvcr89V3DYIdgOOPu7cf+6LunCSOSkJVrb9aklOuSVaGqrTV06ap3rSQMB28IvWNGe1W6ecuPE
ajNSR9zGYeQzdy67cA8qh+WTu5BVv3AuMucjrtz6iD0Xh1HRaeYfO0H+It3Iw0bHb3CY/MJpuNmf
KxON7ZlRCzdPluX8cg0/PEDy0mgFqGHlbvPaV82hJJqUk+zv3+Qd5bBdF4myYKQor88yKZMY2xFW
T518+SHXEbkIHOomhLtWk2OsPP5rwMYjy/ukoa4Zm4QePx1spjL0NpJxEDMVL+B7OKNAgM/3ogkU
nA57fmHP1Y9dd9xh+YdrafAHoo3W1hbskFn6dJuF4tnYk3XojzegEA81MZspmjPl/V/K5lwGVYAq
aH7jEiGdelEZ6snmqCAS13Ym7iuthet7Q2zrtpnGB9LGuM3Viec9CgwHlWwEZuaW10o2nG73IrCY
RWWaDevnGcJ1kDSrT14iYoZUXckKeb4yi1DZ0Qs2JD4uV1XpdYaeI9myRjdfEqHJvhu9dfMugBAx
eg+w6NrIspfh5FjtxqJ+TJDVASORyaIngXUvtNkZMp0JvkjpQQvjuxJfeZvsvqwyRgqS6wA7s9dr
lqRybwl5Klz5HQpMyXVZ5jHCfE6SUgpbs3wJPhuV37h9GulSXSfimnpogbxTMRzVS6AHJ6hMI6/Z
RWe/kxgwrSGaA4+WffvenoJjV+uv7v1S4Q+O1UmG0Yzc2SLuQy12tg81JCmEJvlPQPd1YleMZLer
THTW+tJ343gQeJaYptj6EbCXMgAQg+2mMv687Kme8U7mKR30gsFs6GFg0IRiYkPPSy1Ay8/TpFSP
NPrvqiB3fxC44es3ZLFeQOegtl5qLRcamYEGZPvtSaQH+wIGRNB6kI2EOA2WXTdGvdWeh12RG6D5
XoBeT8+8z+UFybGOoqS0sBPdDgu2ArIFUuXRZZPyOlmxw3Dt/LSo7AXcTx/ooKgy7lQ14KTbxdLm
J7LIfreFHF7IAX4APpmZKqqS1W7jFnt7UaYJTy/r2YB3XMvNze+U6f0qrKK2mA/eQ96UWWMtkTdR
WLdb4b3BRJMpMvN9A9L4w0gR3VoPS7wysI26sxo5aDh4tB0brP0V/eOZHESohgEuC1QX0FcGdsl+
/KOTqnWyhJWfTl4CQnXh0FeRfaRtWgoSrC0mKk4WN0RJbFpTKt0Sq+FETxw3OZHOq1wdqlmuCpmv
zroMf9cjksZm1Vw42HHCaaZT2KTBt+8hagLQ/SjCbxTY11vPgJK1RjH9IUXSJ/Sn7OLvnMfB93FK
OE8LY5rzbBcylUL6gi9oXEXpEnUkPJotVhHf6PeZBpW93/5Nwzx5QADA0S133T4y1S5CbvCoL08A
o3WnsILX7T4pwuelsKbkzXeApXV9ICUcXgaGsT1LTGQpwewNBykUarvYiascAyCxcuXDGo+l59C1
wJNyxuFDdhxJhyqAWdxq3HL879pwDptKG+gMeOyFRq9HPyS+YNsCB94QZZFj63bsvf1zKlXA5nbm
8AnXGxPI0V4YOyM73vfN3A4352NxyQ4ASjARwqfcWpb4O5ZYp/v324Uk+mYo6ZR0BKJQMD7ovgij
V2RkS4iEjpKlP0GVab/PQCDrBSxeNBjYfJxNgjmbFDC5iQmiR9ZKQwQ+mFNRtKC4WBlmjRmQeM95
mvclUvjFmhiJ+N1qMBhAA0YViQPPo2W8q6Nna4Am1Kxp+J71BfT4sA1BszvPUeilI97Mt90xg8a8
ZEMR+V/IacGXgzmM9gUhQr9GLxZjHLQPFZLEmxw6wuvV86mfQrHZEfbF24SrGuEKprGz9pHsbJ8q
K5UGZ5Tut9XBDE2G1ee38kmXq8z2vQG2JtxMObZ0kT8Fj2/wRtIs/VMZ0Pq3LuFWzV7TthWJXtL2
0qDSWPUXD5ZhXP31hMysRB+WkyLp9F29TPRTl3mibtkGhd7CeZujCdm4MvMuiLILIT3wG1FgUehT
WwjxIjwo9ge6K8ycBYRRi7m+wBnyiObsddFyzZkKT7joMnG6ubnjjz2NU/tzp0BW6B6youUlumPH
c4f9lm60YRukjYeaG57oaUI4MccpT0uQ23VM6vBmxElc+APrQ7ojdtWdBh3Y9a7+AH/9W201m0Ar
3uxOQUGhYMeSEVMX4x5R1sgK2cZX6+ZqZJXnFt5lGUO6MrC5dDnmpVDFxdSuWvoj2pJ/rEJ6I4oY
VT7i7pQxvIVE69FVEqbjgD687Gu0e8pJV5Ro/Yv4Wb7i0T22+zt4e1FU6mmAKuXUHyT1WfIljGcr
ExfjlRd8iuI//IyXe7kESSRvdwLLl+cWosROqYlB6nKS2PNTEhhrwC1Lib8JgEjWdbX6K+7IinKu
DSPrM1e4qL9wAsj0bvuDjOBlKIFC5do+b1lfd6T0LEs1ElYpRLeKQ3pZnaIj3G0FH6cBwxs/hj6e
XDIETzIY6txwoGpMJ1RTfLn8ckqmquVXikv6/9upcH+yku+KbQt8yZ7V+8EAnAc97TMcrCd+kusJ
90W9Sziwm/p2YU6xbedlsvs04PF0Kl1xRjk/VDQ8Xi9iF34eFS71scEdpdflJJiECDkHER9FVD3B
KuitO7KWub6f9yMDihy7aoU6YWYhy2vmq9nD9Ex7tWCfqmW4gZFt07Uk/wiV8kt7j2Ck5T/9JyFE
GQ/mmX/A2JFN0uTydzlMPOb306ZZ5SkQDMwtJzPVw3uvpSUNGjBtX5CwzWCOWKvwEpSiEQL4Ko3z
dl+c2b9/4x9AcGa4qycfAJUNPvZvJcemgFX2WMQuZ4DM77kO/70+BG7xDZlByOOgWQDgeL1I7HZ7
tcNDlIAio9whUTLRhQQGoZ6oEAKApM+/PUNSqw19LNrESJeudp3/Qloa8yFC3kdCIIIUCrSSNdGZ
6DtAY8BIbze3XxdDP5K7HZHlR9HrrBKcMFW0YEoILnNFRjpsYeuyzy5ffBFSmmkK9vBLDByDnHat
g5qVO/8X6Q/rFtyvM62jAZrKn62NCapDTvT3RGBzunBXJkuXYt0fqAKbLjHKzLhZrQm1SIHTZ55I
L88tMcS3MpAVheL7IqO070moRFVjB51KMnKzAhG6+o3lTCNPbjNtoPOqmJZIJFqt58WJjPyx6oR9
bQryvZkOPo1HiPYP/uqvK7EUdDpeJe0bsgrXpPVEhXiR8IfFOGqYsk1DQGTGZS/VP1sfWKZ7eWxJ
2GGmNN6u4iesCj2lzjuFT8VfzoT0Mh2dT6LzX3pQD/cuC3OZ9pX9u0Au93sn3lwBSLyvEB7fpRs9
qxXpDlVGDxwPytG+9t/aVB5QBzO5kAmTFnUbABeL+pokeE1vZVSeNAlINDKmClmipdB4wV0Usiiv
VAj243Gs56CGDlGWHdxw5HB/Rp+rSbuUgKLN2POSbNpr7iL9SyZ2bcZB1GOPNrVimr6wvLC2JGwK
Vr1EMjuGAO2m6DpxD7s6AplsJRCFEI3J+KR/tz1mjdTdlAZ93mWU6IVzxCCLskRtyvl2Pfq250dM
R6a5oO8kxLAtNBuDLOWegUyID6sLop2iM3zPU33HCoR+qwrTay/UmDb5sxp3CNKNZIXx/RbkZrPQ
wlkH0mJ0wqZNNhO6PXdmVhl9YWzh4u04vJqogzjfhZ6JEkGfh9OiT5/pOnSS6gfd1JeQ6fUQtgzD
HzTtSy7jqMCQEq40bgKoNbglrJmxTqVnxmHZj2xnwherNB3O15jMjV+W5zojltq31Tzvp3Xegb/N
cQfcCkv9CgqkiaYfNtbLHZOM+ILjjLgbhbVbVGGsYxjI/IkLLGDoQd/tv2+PWYHCh16mdEKpv5HW
ZTJumhw1yh5zqthekxVfldSKn82sxD6t6b/KyA4sTgBmTiuSctJUalsOQ9I+f0/Tja3oPQD6nLDU
r7xUFvWmcl1gL5Sh1oQQPf/SKfUJIHNH4GTpGXMZh3q5J4HZeq/kTiMy6jYnnMZ7gUVMX7hZVdHd
SssFV3+t/kQsOH6XaNJyshtrpTZspCzqerD6xIFZQyep0RhtSJ7QkpWzZ4XMDLykHiyAN/M2jFzV
VS8AGKNPJLcpud4KGKq4cye59vgIXPTMZO1Gjz0YL3fqmQvCTPHY8gEkCZ9wM6IMxRrsOLW/sSYo
8S3xVm1sQNNUSsut44p9qw2EcfL0gKUDyB/T+YdOOnFtszgzy0hEneUQ7X8Mm3FraIVkI0TYxGeL
fHSOUVJiRba6niD+c7uP/jkLPNzc3vL2ULrXd5b6sc7F4vPlOod7zM6HTp+LJF5+Gc9+QldmMjVE
kvZLAqsQPjb6MFsLy8jnP3WToDMzpLCV+drDBR/hzutTxnZH60w1+9ch5iC2Mz7wqy5Mo27GGU8C
6uBgWZUGAOw7fQBqHxtp1RkxOdkH7pY4E5V+oUVTFwTS2T4dK1BDXrfIXH3kZLX3YM44wToSMkT9
JpqZrCsWlnUExg6WccgDgdfL9LMlR2N5P5fUbZ8KmRS+tFbSyEZpPWYj41gNUQF8qoL/XODGB8Lv
GTw2vfrVd4DFh6lkCHf2W/v+x38NcOleXaA1yiavXcgkyhlfUYpbcmDvYaK5SsmoEby7jYEt5uAj
u4rev0zFkrdz+mKINS6qKm3d6dmF9Z6HuwC9HshBn8CsagXrjAjD/VauRHIpAiupgxG1X3p5HWmw
iWHlmQIe9rt5+2z7/GpEEKcGJ0nfaOR1fq1GgTzTERBJpwsGaiLt/6EJmlGYNM1lTwWXCt5u26jh
hvZixUagRvpWXM8mfdBAH5WtvKk7qTBMqddTZ97AKffsEFCz/pneyiilQga93Qe9nH56DTquabsP
V9cdVg5GRnf6GFvkeTFsjO/p3IODmlp2t5fbX9CqRXYJBl5SZGgCFhDHKTWibEbG2pKNt4xnsQV7
FPJk2AZJjEpxA8JzCD5GXrmCsAdX7uLQNur1BCCSyo8q9BW8PM4tZod3g166wYXyFSYEp9yvIdt5
Zkx4/b8Vu2a6eikcjS2E0S8uxV3YwX6VlxnY3hj/ldBZREUBeB3MbzubD720rUE/MCfY1k7N4Iui
o0KpymeHv1w1ChQMmMFtTsvYcbgDivgWm6uxyBmZN390j+quQEbbVYbByNhqVkuNszZJzbDkTRzE
IdUmyzOoqDt8lwKJvqkdPGATuY/TqHo7+yaRtApzD3TG9wEGCZYBrQfDHaE/rg0dEX5mhmpw9jxb
FKBUbF9WvYGB3kt2PvMms5m4bw0mlAaaMZCnIBqlTcW59gidOx7aoW7TpIsG0i2camg+kve2gVap
AyJn5RR+qR2ogErmfskjuoloFpz2zDBiUhHKGpr/wZl3OAuUf2SI8Hf/8DSfCWGyEEbwDyLuKU+W
qGZVNjzOJu0TCPtU1qd4boAjg8e2GIqhldGw2DRLDRN5SxdaBtCIdGAV5WAXHAh0lscKviR834zq
WM/V3TvV9Q7/N2ey8qMdiQrKdpZh8eW3HlCUpB7aKfqfBg73vb3p1cf9ThHxQ4Z4IQ/AQ4J4+ENg
07k3+2e7EKvR5XJ+hkxp8fTXZuobO3PwxeJB8qX8FLlpJFrYCZS74c1aAP1FLSBWua0oAx1XmiXn
O1SoY/9fM3RXq84+67ix9jwZMusraqNvnIPeXnSvBisxgUG3N6gTQPYzB2RKWlTv70saZ20dUJK3
FKgfWSORrgD47ljSuQAZaw6G77NRJNIICYVF2UCty5LzERJPuzHa+/mTCTEzt6GE/3tZRuLJFpi2
mNtXXiOpjKF0Ue9hbBGTA1v/kls+VYa7gO17PoKYI0hqlpamSLmxP+51/pk/DBI07yYlNhAJ8XVS
nMyew2UEehL8TR9wTC7oTBL340b8th0/jzT5zVLy7p2np4ksP/mp2yeXMcboyjx6ABZobiTA4QQe
taxJ4TtYU3PQH71Ju7Uu5+mGGUf8VU/kyW6ukoVXzAvH2unI7N/ZqC6p8AP+d5qhafmK6ji0TF5c
1dQtv/mVhdti5ww6Pvsu9oT8BrgMwnCbZgIYi4cMVeZe35eR6kj1zhD+4lcIF73wbBM8vbM0tc+Z
4CqGYBJEGyvazBATqNvIUQkw311j0yVhf/jQNriB3tW3v0N3LbeqPfHbwGrMCJCDqqOBLaCZX0PE
TO+RrlVM84h3NSxWTicwNLLkH0leA6Z9gQO2+Lw2IB43j6QIlPOVvac5HKRfgD52KmMqLJCPD7+A
xgdtN9a/taCX8wIY1ndA/tt5GyvrR+PTRop/3WxEiqu5OEqRb4htOniGQrayEYP7XCCqKz7GsUOq
fp6+rQsK7/Ug/Yl6zZ6g6RzkKzlcS+eX4RFztSgrQekGRzBahogXbv8WLv3zEvsaNEIeHP+L5fO+
VsU3AJOB8Zq8I2Vm5kFlUQUcMWM+q9vd9sKY4zFranwd5eV7UimAsvO+/tqLMpd4bOSjybOePLNa
8rUmkhFTOMqwMbWlR5WSqhLrX4I2t1kcVfh4d5TsJQJAeMjZiJmbc+yDm05xus2b5lRxaet+liH4
qDy0yMh0tqwmtAK+pgB7dHrjdAA8uCQ6AgxYP77XsIncPu+e0SHGqoa7m5aHD1MTYaER0+EZDoSl
I6ThuYJEIxT8c9K689hrxRYgIzKRAvwrDQmjM3qkscT4eAaw+T6lE+ZkG2UBJDli7SLj4TTZqJRX
rS+t7OwVcRGLIiB0oGQtZ32emdQ7H/vckuxyGDhxIHfh3DcbnSTIMurSyEweg5WFBtQM7KUFeEFE
MynKbQSqOdT/Lgyj8i0QY77mPg7NbZoF2eANPR1MtY5YgWbfM6KQdte5sdqENDtz0uy5lCX8GsIc
dTOEN/IhJM4zGhZzhkto1ruHnJfrrfSkzqIjkrUvem5bUuUb1JuI9Dq49h4Twyxi8FvogXNLAW7o
VfsyliLdgdPU9tO5wWveUt8l6wKdQjdqav2+l7ONe2ZCZWbHxS4+n+pYTNkF89Ts4+6GfZZrSaS1
PUI/vzn/YYbzifoNRrFgarE9BcMuaUt4aoBxg2d77eN0Ma7EsJ3LrnEHCiQXvZqoI/xspY4pUXjZ
0l5G8gP8TLAO4Xh60cuWWU0wCfI5yO6TAdDKwrmhX7ecaagd7VKTOyh4g8S/1xio/cE6O5rm4hCF
iPdqVLGCweHdvN5FbwYxhS1x4jKfcD0oY8O35bIt08nCnLkJ/k9hMAtCh7X03Dkg/Om4fkC2p5qf
S7X4B3TRWk/i5MP6DAjdFJufoVD5m3AYrPRR1wgMMpwZnRj95KYUjKM3/HS902V+NFGLZMFy9dSF
dmFhLue3CI6FWDhjxYeAftFc/0xss15j4Cc9uzPECajrJsWsLMLYzpQq2khRvTtL1LTUKWpoGD8n
a0zKJpTxJHUGb1zPTkgsYr4nHnIGcS8/RTLBKeTWFXqBMukDUXgNqnukjxejkmYWEAd5gxSzEzMa
BsLs/dHxCnui0PH5HR6GHnkir1BuayAvkKJY4Hj8PlWgzSOlP6U5PBbGOO1vgN2z4fW3pqVS8Ewl
dGpwaHjW5Rn7McMk40HywjJz83JUWmczV0+x/MhfiSV1QXO62k6vfWgc6xV6+a0bQhI2p/mfC79B
r1h51Pgkr0t76LSLI95umCOqutECijMU3xosZpOmdVwhbNUFbpBLTQgVITK855eokCsg5nSiK709
YeB+TKMnF+Jbyxg8hNo4YoKCjZNB4iYq8BK/jEFmYolpJaEhO96m3ouy1/hT5307v1RAqDANJRBi
Hu7BQkA5c2lI4HH1bxbeEntuVYTfDmmd+F0rhZTj12L7kKi7n2lU/q+WXKzrcDLB8jQ7lNHwnGb3
QZj+GNKirUhotLmNq4Dx/hmSvykwIcitim4xYO3M3A5RkvQTzhUfXhjEsEHRdBv+8pOry8QXCPTI
o9wTb6+MhoCkw8IfCtnIFcCxP0Ro1g5z5IKK2uxUkr1t2BFFkwIcvIKFBBrBAH/LMQMHDySIltw1
+u3YnCeXJCJQrJiNPEYyuvDSMvxyw8lg2QheL7u1B9Ktp6crVqMjWBzN66DURrO3j9jmN3TWM8tj
30yLcQ3ppRyrw4RJflnw2RlmzQ/+1BX/3Vah+a9HOIDiE2/buA9i6rkbFxWazRq2KbVWauFnpPLX
td/fLShQ1q1kPLxZGV+wGqPAGeNr3OnsY8CPr8egVXlbc2AlYBApm2ZlidMSl5dp4yEFmElu9V//
15IXnbfPDmIB5pySICVE/xxCEDHSPo/Ju+HFfKiuhAr+DsIX/flI7r9jvsVCAfDLlQ2hhA3RGdfo
17lSZXY6W50AQSOxGMxhHxIUr2bhzS0vFtzhnchV24EVAtJCfsbNEHY+lW8S6gIBw2eiFMK+46bs
EOtiVt/58OJb2fHVIlb0rMurf4k9qWg23+bFbMleiKbgSJmd9lbxrbcjOJCd0oPE6Q7SGoKExBHA
rh06llwbWxBtfzRSeyFF1YWVNeR9vEG7nBUZm8lkpfk5q5oWZxd+yWRagT+fJqRb4SJu31sgdBGA
d4+udScmF0XnYA5b+lG26nVlf2Ik3dMST7rpcfDfQmSE5L5U7YjoR0KYTMKbRFgm6HcsqIlUL27g
boGYqXTIUsPjm6iiixPQCEsh9ZLKcmBNum0kXEyeLYm92YBqLswgy84hJ/d6ybE95DatYiqLDePY
oLrBNBHTZ6gwJOOfnH3xnJ2ubGqqlFFhitrsmXjempCz/nkTLQQ/5XFf3FH/ri7KzPRS4j/zQlwi
DE/l3IugDs58H6Qbr9SpVJChgV7w92iXUIKWejqgo3rUlJAaM/fz0DBEIOJ198+IVaHhPHxxgQTe
KD0pnOR0ihtCrKU3738XmhttdojzUB9u31hLvoYlgwoZnr6MViDFDh/3Vp4eWr5OEPbt2ogdEBWu
T8pF+VAyKGsxUMMYjbA9dd/q8hN6wGPZu7LvzQMGmYJSQ8szyU6SIMjW8qJ1smf5eobt1xD9zDBJ
2oW54QK+/mXzVe3JdtDIMn6BNwarV4PkCZ9EWDO1bTe2Vexvjb/IR+Z+rziH7uEjxAOWbhZ29zIe
SRvvoacfqLU1tC5oLWGep6T0O6B1yRGvG1LM84hLPAntrKFM6PCsPLrtkJcAhjkdOWqeCfxqhqYw
M9ptbxpcjpUJd30CITlbEu/bth9T1y7rlk4YAbTNSyp3nEEOETZyLqb00BVQV2yiCaeNiexgo5Ky
sw/vZCvbZnfZt3CT57iJqvrQ0n6pXsu7xdcwKnlG3mmt0lGngD4AbRT/jtlGTqhLSq7KTBPf6QsM
+YeCuFf2AWJX6b3AX6d7RwgViwKmh5itO/HRiXLoTKNQsspw8/icrWCZ3Re8IWo/HY/Q4Yr6TtMp
85rNc2PXZjFHdJD6IYzxIuD2tP7+c2RYvyBEiTLWazsf4KUgri53SF2pqm8QLanirdLwbFjRKJJ1
4r/Pv9ANlYQ32kvaXwUzmr0iYm9Ip1859fbA5LPZTK9pShl/61UeEPjHGvHVMWv0DM7uONZUnRHX
mJSmUYSPE3Jru3fhSJxO/hepVD+qQAZbcg5ADXf7684SEIgfTJaRQBx7No2xmiHb/ZPmQEdvUgf3
xs2oqs03tEhCo2O72EUCVgpznSWp65MZ/k+OSM9ZEuPg/6JkGwSxHgFkYxGBeUqro1Jp1VaxA/pa
kXt5QW4ifoN1aG0qg3LKTS1bxh9kFaL3loy8kqT4vZlLdujbN344CUu4bF6vpaMrHi1ock0taa/e
KymvCjkGVvNHZFkaXw4bWwlv4WPPGpAZNy48rFhhd1N9f1qt8Se1A795Lccsyf/iqdtYXuIgai2C
3i0lyl481xm5FMmw/2iwsGHq/5jJf6dZUr+Y5NU9DHrrFWFlSQHEUwaC9bs5l0P2UugvYkZziE9C
K9oZy//TMGZJ2dK6nznZNOdz4C/c6BJK7PyZNwmxRRUTsDXEMUZJb94HMhozIaMcAmO4p5o0N619
BR0uIveMpvjvXwBhnQiL2pm/ehXX9wsqRwvV1i82GfJ3DHZWOdaL2mQzgQSO5vRc79knxWCTdEX6
s0179/YmcyXFVgbgmr2hC/5W6trM2dLGNuryw/X85IZHp08U/aRxmqap885Q3DGCINYU8Ea4iFHy
dIhdxQBpaMO3uhnhAdo8tMTgsWtHNVhSAMHGrQUpKzvP0tkCdYFHpzafWyQOHLCUGa4Vx6O234+9
IrzvDToFjfLoFNfuqIr6VPyDts29Lhkw9W41Vu3XxUjCRESeTXB7IdTJ5b1PZRDk75Z+8g3zWRQi
RV4Qa8hKr1jFUCglvvyZp1/dbFCOYHTz/utYSSPDSFLAE3Mja1T2Z2010op6GBCODnPdLJ/y05zG
x4ODpu93F/e7Bhf5akoq2Od8DZUTwDhIULLNAn4BMNcOT7nAq4HCg2EMZUg9DI4w50qQ4wjlKeEG
C16I1ZTG9vhk8xN9wko00Q3UVUfDWZ5aRlqSDWeMtxoYV109TvWDpzihySW0G3QBk4H8JtQqv3Sc
efRS0F4CdnYDD1zEDKStct7P4W8G+QJxbepoSVJY65QVxTct9JWT3PYQGtPtO/viJOOAvkMWZtAY
5+c9rogM8jiEyXN+enc48VAulBvn4o7O2Kjbxd1KMI7Q7NOGDKuqaw/yOWux42WjphBMEOWochdA
XwE5sUy/rd+OKYPVum17IRqIeYTUpXlXidVIWseGI0dLT4zLRhym6zpmN3Ru2wgLZQy6UzfOmdrp
7p8VW7WsP1yCsjqJFCtsRhSk3t5kxAhMG6qk4926H0brX4aP+cgBr7SdrEthcIy8CuQcn5HQTgfl
gVrNQUWkcl8+TLdoDL1Ukj6HzOf+157CMFeIpe+1Nlm3YVNJ0n30VUv61QlAWcCcb2KZQuRMxjiT
rEnOc809NgHSd/EBn6uhn9BOUMOicwal4wRoTdAKr+U72JJ0AkHXIEJx1DsQNOFdP8BEX4G/3LOP
bDgJbW+DINGDcxeUeQTl36mzALJyCqMexJoBMrji4tcLdHGOJeGmKA2aUnD/ACVf3dzv/sWkekn5
Mk5t+OFd/pWl/ZoOtzi1PAmb7cQIUjQWmD6+JCTXkyOv70AHutKgmsVd8kI4iI2FfTMlYs0GiCr1
c5Wst+WenENfSMAEvQCqT6/wcy0mcswmOmUhXP+nLPQp/ZYnljjhOQl9RMIojyoszle7B7Rpd5n6
tsqsNq43yER1TbQ8daR9vNlLlwUyNOu0H2RvtZTzpJyFNZjHTFABm7Fvn1iijmpbTAAjsxJm3sR3
Z4Lw5jjLFUKg/hibIbM+FsvepE6ZchDqqvwtREt6S4qzIRbjvGsREMMpZon/16N6Gu3+DKdpSbEp
TuRHYUf4UMdhkDy1RgWg92L/0FH9mP+M/mKeFnkJgf/SQngXWzGenMclfYgzA71wUfR8e/t7/QIh
xg7b4y3GDcUsWq5crDPkyzjYRwxC20JD3Ou9kS0wFffNn4nAG2wLHPIUGpGx6s9CZ3AaWSPjA6t5
hWJhCOi3wimhX/6VCYM79+0sej3pjB+kDGZdcUN5Wh77FMLqifggY5kBb0rFAyCEUiKu1Rnk73Jx
sv4wFFvbZkIYvk+N2R7w1+N7iUf0DEDQ8tDcbI3C5nY4LMAE8uYtEL3Hsq1Y2xyA5gLQ01L83Ggv
pfFqU4d2NuytLcbt21RBHkbaeRXaQl9X2kkUyRRbyBfn1W2mQ2Sv8vfYEWWYAxtJR0S017/d8qS6
zJXKLEOHV2ecyTKt50U8iTjJWri0DVdgJRu+wT9qJOvMXc1vyZqFmTCnPn2iMWWeA/lEwHPvm5gC
Z2g0vOsDsMAEEoQCbLEGg+Uoaf624wW6d6hF3BZzKuwXuf6T6qoOS2RVqks0SZ/t1zWJJzunv+Hd
zsWz0P48btjijp+b5seZtfEIjmNRZVnnI66Nwq4SagDHmPikY3LgPe5GiVoWMqD0zR2RuPM1ztZI
Fpa4c49+b2LekzSsLbFZ2i/9k3bYBGf/eDWZPVlb+uZjWgfUenoGN8wVLs3K8gA4AO25umss/PmH
b2Y50TGhZJfIoQfWzX7/rPVbDwwq18QQC/paokNlraENMboXk3G0pV0ln54Za49GeS7ZhvDUT2yQ
HnTN7DFkY7M8RsIbIsdKDxF6yyHLw4Wdbf/r2NvVLf9SqDyoGQiAhbFKbjknI1TpbQQ1ZzdhQECK
LIrutc6H5q9a7i267y5I6wHLnlsKFVUxHOt8PvjckbMxkeEz1jQ0hFDuWBU+erzXXY517EXfe26V
1m+FHC39EaYvBm1+oIjowoYQGZu4o89WX4+Ly0yUeTPWezUOvIVP+GHHzcZfbSxjMgvVSQeb/wm8
a+LwSk343iZkl2ssVMp9RfIqKIIClsvv02wPMCYgvGC5YwalBlDp49tBlHMKNsNp9CF9/Y3/DSbo
m/arrn9rVfpXzSppH0qZZyT4VA9VT1QK9/e9qlXY4hHjx4GEVwBoqRYirzgc1NRdPun/LXhmDNkA
K334LY+iSoMNjXCF/SCtN95U+LnIIv8Snt/T71veliWUz59n3YIwEsf90YUR0HW/MxEcPYYNmWk/
ec314oNEQOpUWtZsBAefyyz+Ft5y329K6dKwdX4t0048mDhmd8gWd2LtAqsraEhf5TgVxUrS4gCo
kfNtHfq0mYKAyHxoR/sFTaMJH0Syx528THDdd7ljkZ3K/Vx1RvbUKGuGc/jG3Bbvci37UlDYIB5+
JoBfrMqOo/0uj9Bh8GlRBApBRVUw8XeltqKRPvQ/MBzGFlVk/pTCMC8ktsfVcpeotPSSEEEog4Hf
QrFrhHzWw2dIxlG+1MDrtyPX68IsaguX5bFOZ4sIQgSSImiW+MrqzGbw9DWMQfusffqPw4UkHh2+
r6QSbWu0c64T/YHGBmRewOm6xPXO51M5Ah+Y/ofHqdFiO/WZD97EsFhmFtSofNjn6CXyFCzwsS5M
wwGDG+EprFzXw4U/trrG0aky4QQWQl19UVdo0oKx+eyx1G894L/14/GXjtWgZqYj5pHEubWMZfyc
gnJcK0OBqCMTl2OWtog/k+2Fo/uwFYNHazutZtqhfKXGwZXTZT9g0fEiL/1q4fAW+vNO7PXBu6/c
oxNDdCWDhWkqx5Zt/pZs5UYFUuJfysF6Gx4VOwyvudurXBM6snyr4yFx9gs5dipTlrv6xpa090Bs
Q4TYusPUdWtZVzQHvB+MCStoqobit31obtNf/dfvOb4o/6A1bbbitgOgNwQteAXMoi6ggXKAh+GN
w18pKoWwSqGgEQkfR+iVhbrGFKSqKMd16ZLBv112MhCcsMM0m7Uutav5XkybW0ZikFHmoG7coELy
TwIJqXYJu3ezqulXmhD1YQe6esexWVviDvwHEs/yrE/poPNeVTb//xcD4nHCPx6yLt7Yt2MQD1Jk
dlqTXml4KwTta9XW+r/FC4WQntOWZVJ1z1EW2JtUEiFlOQsTqPNj5R+3pOt3gtShVSSB3EYjv22H
FtgdgQ/RK8dwR0JKM6CVGg9s5I/g14YFvYUJQJxOeSvFcT0P60X5rb2JcIPToEKv2XN1cRxPuFn5
dmz29hUlzP7bTnnnsKF4UrQthu1p/arsYnXXc9Z51cxQwGlfw2/wywwxJpttVekzpEcxZBLnjJSi
BkBbVyKYK1b+cYFBDJMb1TMYv87kq4vzchK9Eqt7XxRkNd1Rjx0dUouEb28RdBqngM2LecpQqUEX
pU4dQGkFfTlL9QbDIvCQ3Dy7VXgz3O0EgtF2MJxJ1TkTZBwm1gNW/U1ZVY/ASwopP8ZdcsDuTaLl
SBIN9+cXUad5TXfobGe9QvAXIA2MzMWy1mE9FxCvNIvzhP0WW5PhA9gA/WB3kVlHuWWldEt27lzB
Mz0Lv8IbkEMTZ+E3y0awMj+NkW7umLFr1OXA/PIUCblS8/Oj7zta0sV35EMN4D7Rt5QrhMSWSJ73
AnJl8MifzAx6kvbkaBwdvz2CX0bAxZjQuffkUzVHxsLcoc5qamb9EfPz9ljf4MXgsPqc2SuXucCV
rOwFc/kh1LvbDApYsPpWTJIC8YTc4k92VecXkMq6jAasHnR5ijtOP1iRCV0PAL2bCvHkP6RMGitd
o2T4s+a8wRA6XYQEs8Nf7InLNq4VE/kaLzbBUFetGsUC9p+uZy5vaaspyazCAASJTj9g2epcYHYv
yUq8FeybVVE1YeSkUXf6+WHFfM1ujyrMH+ykbNlNKXV+twGwg5FMfWq6ZiHC7EzmPcSXAI/Zjkw1
PN3XSa8GItZoOnMltEBcbFvRviGpIVSNlTfM/nNG2zPGlFG3L103LAgVYWHM5DJzx4GVC5pMkkq5
oNP3yfwQmMPhp+jJ7DnqQ+e1xQLYeSxiK2TpcN2kFLataqU08Un5i1xRtZxElh7LXyJjC65Fj/DL
QUvE9CzGZDFOGoIQZBvyoXhGXegx1XXh2nvcsiLFCjHlGGMLHBziW6Wh8OG1DXZwcRWWY9UN95Ww
GZhaCZyEoJ3gPEDTXuEgiPL3BbINA02HTqhIIEv2f1RNfOim6v4cOp48CoSYr79iarkQeh9EmYoQ
RN+/XnoiQ8nE7kX7jAIiakCX5UUImoGIqIvydDHCXvUaGKoOXkylAJtl51RffAAgfqht17gBQxRr
6SqxJ+LukHKy1TJjlKpBSu4vtXJKTv9vlZxmhnNAIqg1CpvXZrQSuL4cwq7yLxF++Sh/w7Sn2YY6
lgnnzs0w6X9Ymb383duieT/MSNCZ/jShE6OT+dCzpHuLpTg5ZGeWCIfyPW5E2K6w3Z5w+ogFA6Rm
f2rVUvSXczatxVChdTq9kkQzLskeO0WfHgk/mzioTWBdIFmISxE53EUwEv9wMJ2+nsurs0ap5LM0
84vZzs+xcBx2jAwlpkEXZVriSYPzppp48Bkyoi9LZVTyAw0MfSzI2KBO/tmkUkJD/mtN9svRBirn
irZPiCzRvZbOjWW4eRmZ3oX5FLlXAgj2FvHvdOdvU0qvLM+EvF4S4nqstPnyccXJtS+cojdppAw/
r7AMoe+VGxB2fBwoxqlR1qDR3SBjmYaLxup6BU/hu2gEoAAU4E58wMLv3JOmIaPHxbf9HsYFkHJt
wINgfAzaTfA8mFuoVJrGNGFwRcMXRgHbms86HgoxaB/gpdNAUuHWuflexWJmsHjXkv1XIbYsePGr
yHAHwrkBs2yQO7SYq/cl/p7v6GSUx3MExYbXQkNUSGGA/ObCD+mAk5mt0xfrpzWcg1UtgL3XTZmH
/gstQSSgbEU++NkHEv8JgKMlA3LvaOYyuKFBCpSB4vR+dqplLSrHRK6flVKCi2n5/IE1JjdQJ1UK
f2om93YGblDh5dhcHTlz2iWKfBIzkdY1YzZraFER5BfF0k6937EVNrYb4so6Zo4zSe3jkbk1L5fD
GKLNmn8cUD7ny6PwoHRRZBqDt7AKEhcciiVyKfNzniU1DBEPtmXWKm5AOqSIaKC8OrRB/oo6gXO2
D7jDleMyQ/dqDx4eIGve7O+7W2lEcjsYczrgOCOMUXoukQm0CCnDyP9QtBae6WzcYtWh5zWYWuGp
bSLtyS9GCMoY5Zr+munzE5F0Nz5ivb1azzDRX0xqmc/WbCsC5ewQ1KqCKn5hQ5o15SkcrHj461T8
NLnpNpJoPkQbGkJV+y0yWW30C1S4dDyYxZBFePWhz41if4W6KRnEKlLbk+og6NgINTN53i9ZePOt
W3FXDC3KULHV+TO7cEEb4XkiARYyYRxR8npN45jTJKRSB2JU2B+5o1XkK6OTVHmp7/f+XhW3GpeV
QKL0OIQmflkHmY4vlYPt4UtX0kwiFKEjRcbi9Jf7uCNTGlX8syn9n0/aQCteN6HJCYLkfv3RrzJS
sRoN4OCmoKvjDTdstnOjlBP0SL7mqmGcF7YTKQ3/aEb7sCoASCvFmgYyU165baOa5f6rhKUqlFxm
npC7zfnqZihv+l0kWU9pqBNlEd9a2ECsktl7f2yeb02rT4LkomD6j7Vtq0wAfqTa4wZjTOaDJdXY
SSLkZTy74WEmyLZIrCz8keThLHXpK/K3vvM12wv+EC26inycqyR7U1HfaV9seRC+qK4h4WxX++EF
AqY3sY/zdfWTCixk/Je5StAbH47z23vHz69GCzGpxpr7S9ax7x38f+ESdMFpSFfaWge2PRq6xHiE
egBAt1+LInkYmhP2HTHrbkAIJNiuVa2hMyjAkJBPUQpi6vgEMR8St/cyDFGmBBH1jzWKzPeKpJYQ
tUDvDdX3v7prGwisUkvPCKeaGsHLf/M3MVF6eyuEUcGTufaZrwXdr9gakdu/HEvw4qaO4Rp9T5UP
f3Aff5pbW20qVGvtM+rEw4PXnc1APKeXBknIUd6ZS+F8TCbvONhhmCu1zqdc6pKB9b8AvatKfrT1
Up/alOjrTLr9OYa8osZGC7EepeEhVldCIjzHa7lm94JEpGLnHlC7HR3P2+u/1QI7JuCmxJlIdG4S
NjlEYgG2pjm95tU9xKPPFhXNEV1yUZgMtFOPQ9w9oo2qF6FVySZF1VtFkk1CEtp2vW60IoZT6Z84
qZo3NDqPgyp8zaYcKA8+1adm+MYnhHfBk02X3VvkwcFTxJ6YLAILB/3iKKcx5TEFY4pyU+aOFZzJ
uvVRQS3V/R76hd2b7efxDj3v0Q/+bxbthX+Fc/odTX9qGDPmDertbs76YQeCtQzF/OAVHHiPngT+
b8yYsTwW7wQW3TDSbTBESth3zBDIuDMZBcQe+gCxNc7+mG6UmemOoF1eTdZrXib/5/yyiFYJGIMl
WCWOnxO9zkf96qeRIlZcZCdIzjDzb8WeUl/yCVbj4dF/ta22n2dukbU6HuMo1L+n0objan5Z5Lj3
Y6qs7jfitjOU/jAI1nfTjoy9RfAJWFtTNhDBoW9M8SoZL8jBf5ViOeocCOtMMo/4TnGZK+tRSU9s
73xn+A0fZGpoR7E0gKasHJiaV40Hm5JXygFuxNPGk47U6j8Yt+cqMTF6TFiu2OkkiMfpAz2y6AjW
mHt6W+wx99k90zv6eehjzr1a+fawunMJ+ghv9XejlqNZNMB7ydk8qpf/snY3JwDhoyEqzmcVsVAj
r5CRJoUiHvUULsKxHoWqyQL0G1k08/KaZO/A9+PfwmeTAC9XiQNSroUTwTYzh0d5u7m1dsegruho
tGEHvk6xvVgGT5Qiv/TwCqV/QDkz13WK8qA/JWcUHIFCwZx8DGIHlfc4EV4wnlalIGbdkdQoFV+S
Al+FHYu6Z37jUNPUch7HFDITNA4ncNZVXBTY83pc5MuJd6YUuTJVopZz0dA+xMjcJqtYbCv3I4nM
JjIbkwMIchD9rc8gp3u+ZhvTelcTS/0JatwjcwuBZ/0pNGWwu/xpYfxuGdh6PbMJ6+OBKurzwxUk
EodazkW7dwuBflWJqJZ4k3hlP1EleWKbB+/NHq9e4X4O4tAU0q3XE7ImUo2oRebB2XNDmqwqoC8A
gEGdjLM5d3QzMAvY61/Vm/WrKt82LYOrBffJAxL7ARKfA3rtS6hWC/0abP09oHnpqT4J8c/ty6Sk
jHW8R95LsGO7QsVVJnFXnuGaKAmsqiQxZ492bR5UKfAe/X7JGD+FIjutsLParPLux6AGBloGHoWu
7SruNPaEWB87OaY6OGkgaAqK7v7jpAVgKbLZrjn2zB7127EuFRMwo/EGqn2zJ86cmaWWq8mmgQUy
TlKtH0dzHpAu/D+spv7B5is/2KHC60TyMMW+NYl271nUtpK37iRHFqZ3eSD3hFzKyxM1FQy0XPXx
NCW62bcJeb7MBYPk4n5ZDbPQwwaLxQVHwmy+OQRMB2qB96qLP77Ih4JqaGqURxP4899y/P8+fLQ+
Fo85loC0XAiokxmms/OovJ5vAkc9S6iU30BMOavATUhqQvLlmAaDvWrhz95SLH1mlHisbSD8H/Pu
efMa4nS/8sw+X0N1DeeTV5tnXHNTtl+RXbJyc3Nf4nFkkkmUvjE7z0unkm1kfdRlHw30sXdBbLz1
zQN3ysy/EzVG2PcgvaY9Mguty+ctaPvL9ar5SrTzNLj/dQSpUlwtu1gwBkL8cmRbMEzCgpWm/xrr
5wfi9E+xrlkqSkcfjEX2kHYgQzn/IQmVk31a/Za0QLajHUQ/jjUeu6P+qNZmOFUUbsO9yUnjV+Cr
gJ6+ABBBBgWSvmhxbhk5aPoMGRZPSBTgShscMATcghf7/XjHXYuahe2T89335yGySLDpojgeVMdQ
/czBPrTsaiPDax99M/OGvEdlN4dZd4xd5RKItyoCnsjYzekHb40CL6AP6N8auMxKh2iXKd9MTXbL
RgO8o0F6oF7EKpZAkUjNFy6BWrmgZh2oHRCBJ+dDAz+ces2qk2WYhxqhDT86kWlx671Ezh34iMYF
s20ROVHt+tWjtDEbj9eseo5KpeGKY3CIYLkp2HbENfwY5UrL0ZgM5dH+tz+G+QB5JdAGQZUld7To
jPEDnKdxX6K1hTr5HImlPlGEF4Tzx1HqXXJ64aWcA2PwlgJCMe75BOTciNOaMPkJZqAm6w1/3ydQ
7zDJMl4NdH0Z0vA4dCKPcTlKhqzHsA7dqUU7Ozsbdo5ndwlGts/eAQ5ZXhlDEuvqAAtn2G0uaaEX
hfCsY9u6nQ0cwoV8aVOsq0t4/1pOpasHfX75s+sc7Byzu7BnlvI9N6Rqll6Auoz50uw/SIJZQWvq
6VHKbNZ9CYIFs5AMAwPtWntGsP1E+ifEuhV8zDv253bjbkeuY3z7A5uzAp7/rJQWZNINh6DFZHS2
JqGdVAX65BZRStHZyrh6gDhTBwQBEolFM5YB+27H0g3/EqRpJj0ZLyXMbKwk0X48OAKLfkCo/F1X
VIo0dPgcjK+ZQ7qh1kgjPf6kqqVJ3yyTyf6Pa7ajCwGJG34+++kylOTQ5Pq1wSABPwllMBRfM5UR
C6RGwvX7mqi+hF5XqtzuF9uey9ZT1dNbN3JRmfVv9KHyBG+119ItRmV7CKfzBbOPmdbVFMuRbzv5
eGjP/nyg0/uUc5p4tkMPKjoYHkipqF0FLMWkZHT/aN/CKyikrJfpWimpUUTB/elSB6DpzKI86Sx9
HoN7efE0KzXa/p97iBdfnOEQ1CzNE5LVRrwOEFifIJvhl9YkpafOIOMF5eJbimwSrXB20rzU4LLt
K9E3kMd0H5Nv1ZJUMvbz/UPQFgdaIgtLRIyOMmcYwz58hvscQXcG4EP+voANOFAfOARpaohzWVMw
gZeVOUDtCRRTMG9r0fLnnHWJLNl8Bfhp0zUkLxxjRL56JdUHFUvBo+I5PO3giLD3H/AL9naLEn84
077MNkv4NexuW/mIimbItyJ1ZLNxyJvrKYCsOW86Ur4a1AlD9VKKbPTJOoeJCV7tgNVmy3Yd577z
o5uDeY2flmURoBMJTK6bM2m5007cLt1iGSqaCO5ErgputwKWSVYqtgmk2L5bqvZ5YhTB12vyAL6c
LEpTZjLfmFGkfExuWZsdcP/YM3IUXhKhf0P2wBq74uOKRqPJZQUp+B/4kM/6x3nP+eLana1RewOq
0bbzZCaFh0Vcw3NXiRj1OdKlkZyd6i6n1oj3gZFzwj5/h51LtlN603MucmBobkISku2xZItZjI1U
dqKFJPJrEFWCAhy9kS0O4kfgzhfOaVDg0Zu74PTLRVkvzjERtVNN0gIkv6IIOHjCc3m3iSxWfJO+
tQsetgL9El3PzS4yXKAaPaV1P7dzPomaZCWZaFY4GaaCdnOhsMsVHK1CFpknM5vOExxgo47tbT2I
DBAjGl08bx12USuTAGpQxrwfmRsIcLdZ+0omLXrsVn5L2RlcYUNQjgRbitinmIwJsiO5lJjgKmOS
4/NXUKFCzmv01J2Vci83s2zcHCGfpF9KuF3AybBnsg0sQMfHAuQ+rYvHyF2Z5+1LL95Z3Kf3vo/9
KAJrw+UAjF9QnFVYFyooU/luaJyy5/C+QaDd9pcxjENvKqJlUO+7PSZTWonBVOqyax3W13l/6txv
1CS04oIrAJL/QGIDL0fKEbx1ERZPsx94rOwOE+2HhY1C3pt+yoyJKx2UU55iJ/zK8ghxO4haNXLY
Fx5u9UO9IdOd6R+ZWkrYFqwRuHlur9KtLGPcTx5HF1ztOphaGUcaNbMRkWwW+UBdYtV+qMR/INIT
1NNitQwshvtkeJ7mz4JYWJax1BZCG2Gl69+wkjRLwvZH54NfkdKaPh4N3QW54LcZ5eupUASlO4fe
VJZH+Anwc5a+2lm6Fi8uI+YJAZXtupHyRD2FcScTDDA+LCvvVXYa7MgJRG1CbFErR17zcBgyD5Ci
mb1utm08y0Y7ifXK8tHZhzRIk3f9hVTCD1GFWmLhHWjm0xlK0kpggmbzsmgOoG1vRhsds2ww4SIw
vCceEIZSCTT5PLnLZejC7KLsCWv4foUHBTuCLb9CbGKUEZP13XQp/JvX6gmOFc2NTZcAN/Hkp0PR
pNjmNkjGL8oqXiz3IZpO+ky5RsbAUgTVKetqJP/fZ3pzUxOw3kr91Ry+jjaLVsZCEE3TYnE+F980
lr7JzVuwapqGDbxNI3+0lLoBixxKmkd9hREHExrBQMg6Yk7KdzmMB5tnnkmwY8hxh9dVLROLnMrq
+HxTmRH68YXe1g1b3iOX3a1G2tg66dU+z5pEaPupwrfdxv48OgyoAo/X6d62u0C72a+oJ0bmPefY
e7ygVc3P0Lv76iRBDqNy+OOvkEbnUZWkd6mZju6bZHNqayRA3Cchr+qAVv7H4ZBrcY495a1MdVo1
QXX6OBq43nE4QOZwJC+vX77UIVh5yWfSssOqy13+pxP+vj0rb44kO7TBnv2Vc5uHmsEKMucUsu3c
pCe1Ty99YFNWyZLcn5/ptYnormRbO+revOVRL8KHk18jvQwJz7hXWBguWu3Ur3Y3WroOS90zJG2j
38lfAJmWw6oW8HE0BJsZTQxlsFe+/DoqKOSGCJPKv8o6Jv4zqVJCNv3+U0Dw6kJD3S+7/xtEbQEv
hzo2r7t9MjBjMn6Y0FKUKK6CnMzVu3TeQ+panzTWUrar8Tq2x2Apdqzjv5FGAqHi/lbzwE9CkoIr
9iNso3YWwWcAysclNHHdRWQcFjnLnnN+hq6Kw7/Q3bA7PAnrjjAwE/rTQlYsk2FeG5oHl8Nce16X
PSyPaMI9och4iYt/chBu76XWHKc/IlT17f5Etw7xU7iy5pr39ohv1NlQey/KzBv6biojvhfpYmgY
GDu3bR86vLrEAnWczCGs3ljTIo7Kh5gnzHiOSgg7rhkMa1NSqsNbh+5oy2O6tKEAd04d58j6PWl6
dBgtwk2zWEZAcCcYOwxyo0S3ECzzC1qyewIzI433TRtpTbk6bLjPXPC7p8MgiG6C4FhCVdkT0xnd
1hqKBJtCA1MKDDIvF3ijLpVqESL0SKRQ3Nyb4pV1XPPiLmTGc4ijsLHpf0FaTHIvfVJSG8YFm9hE
VTa2T+g3zvUwidUbWmu1Uvr0zsPxBLYBermr4jronPckrIf490kamMblElzlmMrlowEU1SOD5i2n
B219fO8MSBuNR5OuXJhF/9jF/RsQY3g5s1ktR/kG15naoWkEnnJosmHTM2jdw7mCHmf4BTqYKrax
R9Li4MDENQX+AedECpXw/9kYHrVCvco0DgCMLyDOpbR8iTdr6HBzcjakoCHiXGB0WRrgLPqkn/Sk
Mva9Jhzv86r7X3ShKX8ZtKmxtJ9giQnGaAjO/CwAhGDxi7f17Nq7GYrSA7J1q+qJaHI23Y5Pf8Gi
zbUkzZv7gQKqjdCvVqd9j109cUmwpVlnO538Mt3FDfUnTA2LENM7u13SJvjPtPfzwicGLmVB5tRN
AyK0qYkDp6uphwVcvQcXfj3f37l5dGlsiAw4wwJ7nMQkAf0yG8FCLfIrNFPTUwlFNCRgmeENMYZx
L9ByCCmnlOVw61EJszeF7GySTNopu4ybAPnyepoI3UTF4VCgzdebeO781z49S3nFM9rge3rCX2ni
SpQ7d3VxOoEE4UwogePYaiKAdgUtV7cQAyCjEMRHEa8tmE2SfVVb5O1LBTP15KROqzIBRU/SrbaU
DAPpou/obgUF77BOVkGqgKVjbFRkadtLOdJSRVISbX3mWhtEQpW0wsk1EOkntMHqZsg83L9Ql4KT
i2ilg9wJ/OEo/swBrs9eKMPu+OrfcCRUd0p99sHzXpuPYeYEHmEMgFdxHvTpAxm+s8Zrspq2XbOn
HKVdfoLsAs61A+I1+1ChhmqFuG3xZxiT5F9rFQy6z2AOeDvjy9bBkJ2sARCUj6vvYxBwQI0NVEkF
+wjtjc2qgniWlTidhtawE9kkrjlymNto4S+zcGyXk2SOF1ZPeyyVqjpkwA6liQWSbnxEcqFm+Cqp
GmsMlllmtUQ1EPsyuVxNmwaBnoh5P6W3sa09nbthYvnqsknUkzDWMe/1bJEpDzXpaHHPo4+vCtfD
OwbXqwkQgF3RA2KQX8eNlTA+OPV/bnA7Z6m8hCzVwjj3ESh7Kd5okzDe1M24SFDOabCFXOQo0ZIv
z8QogE7+V8gyE3X0d1tc7C0p/UDLhuLc7zHlgWon77CfCoyXzuc2ghu7F7RXe+9ykKwsLqxgXwOu
kxBgvI1bIfaxpHMkHbbIRji/NxCT5YA3WfHrlSkMBXZbIxz4sOH9okIqY+Er/+ZV39kUTyZ/rFoN
Vmfbp9jr5Axg3vOkEaXYd0ITx1hx5R14UF5SvCuycrsaY7cIfxnKtT6srHV4Ojs+j5mIte5KNKKc
yuyVONZO2ViWWD7wRUTO1BGV38/fTxe30g4vJBc2TfmsPQZYrDtr3LdfDtGnGiXOaMZyETmJ0iQj
sVshyT8WJHuktLXntdk7iy8I4JZc3pvGw8AjCM4Ky8U0IoKus0KOdbKQjSqAVGjG1fxuGGmSrbPF
gbgSjSg73SjKlRyzk4X2TONkMRjNZHI3fSoFHJ/z6qr3LUu9hiWw6QypfyM/vI8yUAQ0VySmGMj9
P+G/ne7K1id/p8kiOJjOM8EyLHe6x4lmBt957bQib1eBPtPrJpOBsjIEUD1l83lvXpZfE/Dsn5Gk
ckRBhrgvbThrhGBzeYEfHwIg1Lby6GNFKEueZkF0nI+f7dkbT/UKoPdCwXuGzxy31HTy3vtft8EO
3yGzGeXZ7GVCQeoB62bgLy01OOKsFQiO64X3f/DBOhAg0yA3j+pIrilWknziSRga5WHAL6UExA/z
cmiYjwfoy2JoySeDIf/AJNKEyRI1UjdY6eZtuJ4frLoOGzZBxOZD/v5I6NYam3hM4HSLaLoaeXnO
H5fY/Jvyv/9CmOKS5qFoO/o5z0/gC5h3bzNnvHbwBh9ZevbEVxTyeys2rcQ6tspFRo4TrHQ7JrzL
Oc376BqnYBPCv5+R+FonSlftSWnEOUahy0bEVFdpDrHdtAM8TTZhmQcrL2vYgaD7lS8LJbsGuY32
wwERo/ycn3GoIAQRkSEdel/b1JMDqbsST+C1rbjjRNN3vrH8d2zZ9jIBtBvGvktj/U+Sxnh4nEGm
gPhiruLZQxmQfIQH2OQjhNfNW7Mms8it0tpmHOloWjmKXPdxDWxY5rYoz8QCLVo+i8yvX18x4w5U
PKkj5Q16JBRLOUUER6m3sfEAyylYbpjjdpEeRX70vr50B5dnhd1/aR/P0cISGSEkiNhqhi+gsABn
4iXNFhC8U5SEK3aTWKMDdUEQS1yv+k57q2UTVC7FHeG+YlDiTEFHm7TU5jky5eCIJdY09DDd8nC3
VClcWASOuq/mYOmuQGcsrPnuKL9RSx8W3kIXNGSKiwsH6ip9JfUaJWAQGcccuAgw0x3FTUYwN/3+
wndiY1xXXsShCcqU1cgDio+yekHVxsozOo7Q8yYvwYPpmIjzFGPAA7+4JDwcD3VNZP5VjX/xg5+t
z1uOQdAI1xJphkpwPNbmKY5wxR8OVj93KRCXaJ0Jwol7iizX2c4SjGCCH7NVKqw0leruhew6y3xv
/bJyiaqEBS7MWpfzlgnyohR9uhCh/x/G6pZC++oalHXM/ldrcCA0WsY1jq0nWVZperSaXp1a+1Cu
dQHzSLq/doQ4gN3TEiofqczSsTHqAL/mg8R7r2XnA0puIE7zmAci5/QmAgtUtCkERjoIt2GjRgPT
Y02ga+Gwfz2dFwKsjDPPgp55rw5MdSCxSb2G21ayrCMw+56Rl0XlvTZ902/NX8M8wUz5zTRrUUHc
JwImwMbVsiVxiPC0qWD5LydVdbdOFTbHoweW44v1PpnD1GGgx7hyerz77kvWNTCquG/HWdAR6b8d
CWsY6TOxJRtOSTTGxcUKaEDWj+734Odgy7YFMPL8+v0S5zqXcCSZpV1wKmOQirkjT0/6LfRXk/ci
B2t4MbqicboMDbqiEvktedOOCIlbLNiJ3MrqRgMsDkiip30Qvyz9jSFir4TZtA/sLAS1GaWhA9DI
nFgMICULX6jG1h7M3+oew2QqKxxP3HFv6RELY2HffT2wKnhWc3X5lWeVCdbwjvAVodg0QftIjPuN
MJlrB/TyIOftmX25g5O6pUnxtD55U63Dor3N+afg22ZvaTTkRMHYZFci4HULkK7xquK8sxflrWnZ
bOgc5lM9oSsN+r2Prugo0eESj+2y/RNr2xYmb21oi2pkG2ORKfSwJXQ2UkLqJ14iQNGcdiO6bXjk
9IMLYGvs2keR2bpaQhXYFtUd0c4JTskCiXGeVuGh3ULZb1ERN0J9end+Zha+nsq2NkZJUNCSYxal
0EWmtqRV6Ck2Au1AKbRDCqU/kMZFimSBVPgtQs3c7g61bpAI2LYz0yRn0WUoGEeX0q/JgxSDFFnq
Qijbu9aZRVfZ1fJzoLOP7efSc6t24iJoTPDPt7VFWeW+gb4TcUUY3k0ETdlgNl7QNoNqSs/lkvqr
qA7m71l3pXsdTAKoS/5YXO+923oNSRRO42Xoq5ZBa9pWGLf0Uo5HcsHE/jEovjTUzsHePoJs7S+B
spPE547whpnvvoCpz/WYLAnUmQP/5K4NhDSxhKuKkwqXbmWH6qFK3xO4E+LOIunkUMfuVpbtzFGs
cq2NZZ5OEPPiO83btqF6rnfobHdYvdis7KDMaDBquJY+T7UNZpE+r1HbFflMSX0PzQ7/2TxF3dtv
2YUUXKKo9S0PBBF6eCVx9jXj8NDdLjK/qrAByVjXlWuy506uxD7ncl+y2EI+UVI1Bk3zEpzj2qIJ
chGOcbcUxJpJD/eIqZR5+uXd9I0AqPNJorqOSys3AkIgM7q/z/Bf+wZW8I9zKnQPIVS1Djq67k4x
n0DmF+9JTPoG/tEdkkmUcmCeDs7HSEBMRjc/2bU3+CYhPej5nDWXUD64oMU2ny2q0UMhxFU9nuQp
Evm65/bKuVKoDExiZjFCpAGAOY2Dvo2dabuiwg1JZBu77al+CaItNa1VHTBKVpQNuyW5n7ON/WtF
Yn1wQ9KGfvafeAIRInGs2UWI7iT6X0OGJh0DeLnCA6nxqyU0hkQhxQ3W/aTm2g/27Zbjv97H9RV8
xy1IiQ7e0YTv2o6ArlOQzsxlp/HjWOWXwXQSfZiyzgN/2CcEBJnjlnsDF375WXEXCyT7Uhu8Zf+z
ORyWE8PgFtzp2paYlaFRkF/ilNHUWwueaVTPsfpiCx2KTLCqwnMZ+NmLsLc2NaM3jTfI5VL+az2s
h9djMXYlr2j0hOxUgIv1SkLRvBbc1zJ+IIRj1nM8x9+zeD0fALEcN02ncQAiJ7hX2j++TWqaVDIh
67i0gGKqEU3lIclBF9eDC4ccwE4ZVNGmbgn5YGAdo6MqJj7absHXhFbnv3cTF37D53TYlLDA/Vdc
So0aPgRs39z57h1dW1nUDNoVVd8g3bptngFkq+KLXTTTi0FO6tVfpGsfbavGMyScZCT2G0+2EG6I
rCJmOh3bZM1S6VmqgzXtYN7+z54DNCdfYGJWQ1Q64Er5vZYewBaGhGGu06K3q3NM6RcL63UF7jD1
D1tgGU9UMbcVeQt9pBPIkKzk37xuABdchuucWQhdvx+5f1AFdOvQ6J6FUEjQkgC0+/woXUu6fT0Z
rEGhM0/bcNPWhfUS+8lprQimTfbXwYFGkPo+ew09Z2EjZbq52aGfYBpI52QOnMVJBVGOb+W81U0a
8T820hNMwtZbvbcHcxUd5FHqVeyTsF6JPCzmGaFMC8WNvKx+BqQ47ga8S/YD+lCpB5xtI4R3sKGz
BQm9+IYeFa2fvOlmQX0Fbv0sUBEVaTha7nhZZOGkovLU85nAZHeRiTZ01U0zzS4Tym+kaGQI5hFP
sNtOAef9SgxE/CkFE7JZuFUEwWHxUT+wXGIgT2aqdOZMQprXAdSKe2VnCb6AkNkbxNL1tupBiqXs
QW2WfbY513GNC1xjlJL9JGUrLscASu2xjCzvNMyj0n+EUgyj2np6B3gLERvy5bMWXmXJKu14CTBD
8WOGiaJj5w5z53cwmj+XWdexsUIHXSIihbeS0L8341QrTDd1dY9D+cNFyDFggY6QBRECFJM/xpr9
0JBjFjUWfE5WXe79Z0uSoUpi6D+WkMOJF6S7QGCdmOT3k5D10k8C/TniPBk1rJFp9ItsBuILNX78
aKruWR77l6L1NmbK7KGy1RuR9E3vzh9lMv9Oo7yshpDQcAwPFlWdK7ZX6v5mqQdz550FVm6xjxN8
21+bEuD542qYI93/m7K0pKb4ZmDNToaUeEAYvuiFo3yUcHQsteEGU0/cqfBLtiqeGxY129bygBjq
G1ewJrI2IrcgJe5a6RNiWB2h7MAfa49ZjqqR06T8oB7ehabxGjVFWh9LrZV0VHMLjJQll5zw3w53
y+1KtchvdsjKf/UuUktgh4SZozl0XSrqgg1ISDKSdPO2BjHv7zGa1IfHmfjPcYZ7aHrFvWx+Zbhv
zXNcwYyijTUidQBYk36oKDLwFKQG3/erM9Qa57KLSksW6xxCsmSxFhBw0gIC/SxMte4boXC/Vbip
MzsjZ10xdx9cgJYbFShiijUogcBwnPtdBZaou4ApZgLzfYuo0zo/lf2rcskPAs80R1KK31IXF6ur
jvNJmY/zBbZu1FBskwTooVSXYmturJfeBeXbs3zoW+Hykf2S3YEARmAB5fPRythCj697GugJqivA
/juRFkg01iUIzxrtPEP8rzc6GYvT9T03q8Ot6AqqnSQcrjSg6oYPZ5f6YA3y7Fs0qhqoknqqDUiT
pibrotMXZeIJ6L3o1zAId/V8RhImTC2dMW50Fh3S/3TCcHh4CtI8nHcy6iN4AFo/4oFS1/Lxxj04
lS3aj057buEfqYVYrpQCvS3r3jG5G9aUKgHpkXNZK5lb8qNCkGoM/upzV7vsrA4porrBlQjS6Y53
2LNRx/b+k9I87dJGZvUiUmfNEeByhsn2vaZKe/eMBMvkYELuHEqQDe+B8fSh/dPQ2PDlyHHnf1jt
JpOrCJMmOo+BjBzN5wiA5lfm9mcDwQBDtzAqpiNrLEYr1VWIawCaIO+Hl460Ehdkx3t4K9BSVaPb
a86FTEw5M0OgKPC1D66i/J9uKLrkvYkf3HEu+y7E7vCj5k1sTF3c/OhPG2tirXo1ZeQ6th3dV9TF
tIRuDcoVF7PDw0ELfDaLDolTEc0haJMvW7E202guEq9y0SqwZQGwV9VGRz9Lff1JlbhHCnZ8VipP
T8h++Hmyk0v5mDTnJKwbueysT9O2yyaAC5ql6e35X4YD7JyPzSnwtmWbQgp/d9pkAyT+3bmamqEO
fAr6Zp1aXpgzsclUpnp+LJT30S4B58QhEaz9vR6Af4TjZKUo5xQDBIa4wBP/MC6+ycNWPRGs0wxJ
XjyyOxhS2qUbumwOQJgMymdHNTiZ2GUM680/ghrYbaMk0NZRrGCuOMJbObN8bnTD/eHWw0G8bcBt
C+RakHyKUvGNni+mtDPfnv8heaq7g+ROUcn67nIVvwjl+SB05kf37GOb1jPYGkYOmjLYnQr10/gY
JMD3AgSTAYXP7FkNCbSN84BeGhOlBCQuLYwolWbffV3jyHCRoBmw9tikn0qwxy9mOL4spN+555SG
xyHk2LUcjsqZqvww19rjG0KHk9wa6snw3nK9WNlMtQ8wfCIoA9/b6HcQwLYvAg3a7hzd8VZ4fzP/
DZqU62TUJ3Dm0ZVail2MVS76/+z5riYEOvePtAC4rDQp4yIjiZUckRWOiyWJiiHnjbd+TOj6BIeA
YfFa23k8p0RHQS4oULnlLx9HBkVG67QUxkH+y2JC7/+H9ripuQsAqTf6O2qC+/NUuLhVl6+IAgOp
sF+VthofQjWaTAuy1GV0Akc+bgRhe1BlSTRxIU+wm9J7uB0x0KZRt2aM9ouPH5q9L3d7xpY63W6j
/67P/RFqv/X4JBrh6dgL0YWUW44X6uzSI64+3YJolKYmcFbvqf7Wbfo+jchbEoO/peDxqyXFe5R9
l9ESx+5cs397rSdARR48+fmWT7KZ4bKL2RcEIQL4n31FEwxQJzR3zoEyUpJNbogdYMELmWLxFf2v
FlVAEzdfHyFiAV1ieHC1Ariz3VR8hy9ikdeIxDGp4X1k7w9SDQeOjKw2bU1qGsmTk8zUG3ZkcKwB
lWFUXra19x2rjPNNeCYQhT9Ks31oW9s09oXsnH95Qw4qd1qfoO/st+qNNWwwluDT60Vv2uKI858U
qMPVrEYoLeStFTQIGZgAIrw33OaSuNY3mQwYqJNYYVf6/epoKWvRNAIlZBDkZ1ay2Kj2bIPpuKzK
iF1dxLllJCa88qTu2QogPstJxRYF3WBvy1OgqVzxT/mPuSL17FEvr3gWtnMXaDr7JY907emjXpTn
bthk7gt/XS0N6e8YJVaJ/htSJgN6k6WFxCTqECregBgGM1gpIf68VohHuxPa+CccDd+lcvczWms+
ITyE5NKL5xkPwEvJmWqHW+T1EZs1T3fBFCIjsk/QZ1L8cWIhYJ1bVOXK8pDLiS6KLRwpct7AYuLN
AWaInCniOfdXRpo5pTPorfl+lLiAFcMXagrC1xHWw9NKhIjL/1qUEStIMN5IYklzw/yFMEI7XKJV
gdMG7tgKGd5Gv9DCBPz875E5B0HbbptNOlBLn+bx87O+DuL6/GMm9CtZCnZRo1XRJc0JCYP1dSfW
i9WpD9cmKDEC8JlgH8C/nODfycBtc2j+QV2b228loVib//PE8t08BiHJA3VefOqcv0yvnmmbF/fA
5CgcvRXmF/zta6E5vq/ylFSnHE0p4Sa/ZC6AWxJeD9LKFy1sditybdicFVmMNmXTld1pCZwfb2rR
ABEt23V7vPLs+CVROyhrqtteIFiT0LcLCnvHaXoBr1LEtMsLF9dUikSp4JyHRlxQUMPV3ewFlmEV
H+9X2YxNtGlQwYTpZuQLVNSHUcA/epRH8Ay3nLpzcOxiXKB79LmKlT7JHu7U6QpK1gofMGrL2xuJ
8eMeEgZOuuVaGlsNAY40Bt/sz/xKXDxiVExyl7EnPBAxP7fgnz66Eaf+dMuxGIp11nmH32IOiFme
Cn7frin/MbA4vfEbxh2gfd9pdyvOxRevMKx1WZEVDNUyJhVNFPaM5ovzjG6EhmgU+Gqj3REgsSax
Tdml8VX4r1FpJsDBcIRXGce5ry2jd2YEtdg1x0qj2hSDaKr8Vt4nBl4/IqhkHMl6dNom0Tk+7YTF
Krlpr7rbwB2cVvtw7WS2K1ZTK5qD7YGyei3Fa4d0Kcj4NU+x73bciW9mXIZCiHw84xygZhElc5tZ
BPzri3Q37X3k0bTu1rqDRp69evC19iggYI11q+dYsA+h2PfdRPeqSnC97V5PKEda04aOi4xOzrpu
n3Bvo/G6JXCx86XRySbAfIWokAH+Z7BvfivMEJPtN+a4uFmqaq0dObPJUuptkcTQoD0iUNv0DKg9
ziq8D/4lYeFk7qKEtxGeYGp8afv2GzH+slMlywEACu89wyYl/i1SGLaHBwZ7F8OVPLnwh7pYKI4B
6TiPpSBReCMK01JlkGABd9omIQbTz82IDmK9cBi4gZqqeP4+3r09s2olJPbD6uR7w8p2RQLAzk7F
S5GdzHzI5hin2Y70g/qUl4cAu9wZ8BdgNwIBbt1mDpMKrvHq929N+a2E6h32k0mghrQoOHsBxKw7
ykIsH/Av3jes8oesybG+cGdC6igQBETKOiyyxoEM87IbGBsMKDagq3/D5p0v6rbtV6LnUdV8PDg6
EgYCNBk88Sq5OXK3apo5PV9ZyyZ2ocTb31XZ/AnEdeYN+v7TNi6CenCGr/LPiyzHrCfH/JTdnxEa
g9JHDT/6tC/863xKJPjoQB/Rl8zNcAqeNAp7Y3b7C106UrPz79zZpxMSBpuARMF7hL7bOwbZNOIz
EX6rA6ItPQ8tFXvMoKmN0I3RovIa+xnv6Cn109HkhOCkXtX4GWQQ+GhWkEVX8jqRHv8NEdmukzVt
IgRFqprdHsHH2/QB1AvWUmNALvnpmkCPtwyIXQ3bAc4/haqbLie8zw1FrQT5s+rzkTJwW4IOqOvA
H318tPStDHv7WP7bsUuoXfBpXazmLBFjS9e8Cl3dFdU3Nn4Tpi6LASn2TxlEnxRgnyxuXItetwTO
1KSmewid2LfO7fm4wpCzhswOccA5tVUfaSIhqnEpfQUigZMi0WsDipFNKOPPQeWy6QAoXe84gwT5
Ub+HTs1lIMXKT+6GurizPwuK0D5TnPeXkonV2qig/y0c2STufE6L8fP3p65BGglZO3bNCYbYtu5A
OMoegqTbelMwFehum4B4+ajnsSsbYJe2TAmgEnb8HZtCPf1xuH8dImQsWjNhdjnCbUd0hShjrewD
Z+k6hC9BkzoBkDj7O5tHRg2uynTX5hDicKUqATLnUce3PzMIt/7VwxLylEEcnAeM1oxIGn4bCFeD
vu6ALADKficWoLWszlC5f71vkdMB+4Oiyu+jT//Vkb29fxu3YpFKrDwcCLyjitEECXuOIp1+om0E
rHrjvGE4Kr7HkDHtsK1T35/aC2yl3W585LHe18ieCsdTB5WIDBAPdmdxOXDw8o5G1m8/NugifEhQ
/eeolQdllgaUhdDW9VgM9lEUbpTKVpr+wpWj1wqpEBwsUA++qGeaxNvPD7JouYEvII85ekN1Wcuc
TT7EZj2OSVo7egssAr2XWtVGkVMvllCVAiwNmxnc7PXRKW+HaMAwZdze/Rl1Fm+6yoDcShs2UxuW
JAl9OUpXYUI7hQQdcsDxqeaJ8O3jFLlDGwKcOslHxeyRKB12cG9LHl2HGdyzjUpikjcgn65CZB/8
HfWJ0D3NPQsSEBYkfZqyrkIpF1mI4CVn4vnKrUvSBq+uMz1NnCiZv9fr4kY0t5xKQcJHN5TKH0He
LA6qdu78apAV8OgIGKUZzBQJLBKJ3Hm4D29f7KocJTJJKytv4+9rIXZOsZmWQO2Ys51P4HHYxbPj
1mzhq2BkwQCEO85dmfe6V6IZNdaaHol9MIyoa7jy81Wa8/oNtxFweuchw3+pjJOjbYZ10Uo+k3YA
7dNtDiZzv9FJNj0bpKor2lfcuz9ynODwoE2tiJ7PW2kGM0JIzt8mhHeRtq5qiBQiEq7Dp1nDd7ae
QdeVX6a7rm5CJNMJfhhyvTMgmdOm5WPCuY9VWkfhMC7a6w9rrn6cHizeYAy0Cb7NsE/aGR1wiaA2
rlyb6rkqKEAo2bJ2SH8aJVn7H2sHEDPDJuHAeq9jxm040GM3/JWfpHJcQmGh2Forh3mfuM6GKRae
x3XfZ2OZrQRpcfRsZvps4brj/r1mT5WwPeNtNSkfyJoGgkFz8gzUBGasjHcP+YcQC1DDbk6429Oh
ne/6qx2L97P2fS0wTH/7oOUkafdkHpm6WLeCl2S9Wvx0ptVGy+VKtip88YQ5+Zl89/XKfU+LrJlV
hV554TzsHLa0fw5balbSHAIzV/IbKktMALft+SBbNkL9/gaOrSFFeOf4xEFMQF5sI3Upl1S4SOTo
KjWabag4LMHmk1zXoMRr3TYE+INcIgo6B2s6EtlVdY7MU8Jo4bbCtocvd2oJoqvLbTSR2nEylw76
pVqXx4Psgz8i9ArqEmnjS77/NAF0tslBhIhr8pg2ABm45EmlE1N4pA3rodPr9upq9IFoKZk7881q
Uj1SVdbQMDSO1QmfhBwuRGd/T7cMJVgeVpEgJXd3nGoflxSeEfEloIH1wfa8c3zGyZdLLxts1GpK
1cffa/F6uWw/uEsNIih5nkVAZLSyNW1c3u3+EPmEU9fOC4tKCswbpLbYLWtHFyKXVSPzNGXUcpeN
gNzvaOaUIalI89d8YKV+X2o39rm9q6T3RSC28PDNIi5Bh/Ucnt4ZSMH6GUPkoIQKO37VQuY9x32O
lggZdgHLr+3ZAPvR2yVQY4kVMWp9SDPnxWfVLSdEu0/qHpuoV6gmo9u4yXDARy31MdEO7loJwfPs
ZX9c3NOYXwIm/b5Z1eilLlZPIu02a691UcqD4UROCLVRaY6rjVI75yrbQqgwKjT88ZEUDqZiSOvX
pDj65Bruj1FAnzbcWcy0SBsFwNAl8DKQIwfJ945FBfw4VqfFb7ZEWP+smCTWSvNCbV3eHV67Qb2r
AFMyhyx0jtwBNNOSz8WmoP1bxoIf6R6on0GoGp8BLvDjlKUeXW9n16TIuV3tpHSSrSTZDe7GT91X
VpeDaKqIdP51xl0QaaZmhExlc+zFSkFfDgNLEMcXz6fDBYRsGkDCKTW/+3NhGUmDZhngEJDqwHq2
llKp2iAOrWVKH5PYwjMhgeVpypraYj6ypOEzkJj2SCjNSNXXs4V9eIWCKZamjQCKzbAnKXOfiYtN
d1nSsMNv9j3huH1GQvSxny8jNwyyTNoAXDwfby6e5bNhWAwRYvMGNkd+eZRVRIecat4NfAVongRs
Zov03CeXN4RiZ56oZeb7lFTffv+3iGl0km9LIzaHE4jmLJR/HyVhWxyjC1HRbvBzAZQkp9otpQdJ
RyShiHI9mLDPAtU58ITyWIv0sY7y/ilDwDHMlojvDy5MLKSp4OaVVEwy1Kc7OzMGCrbUnV/TvCHK
keE0lNOIZKNEX/hPQW0QdKs4LG/udwPX2jfx+q1ceoChALAqusemq4J+NkQPgAfXk4r+uv5Ws7+2
JYgYOmz28hZypilJ62JfgLKkAiQ0Ksyk1t8jgIlmqCTH2hnwSCwxNrkyWpiFx4TZqMIBMg4zs4+F
2ZZhdskfQIoKtwrMj1M+BaNRkK7TcjUTrPHhAO/LcAPGLzGYJbAN5FQQIoA+ve1X/snjE/x89sM9
SVsbxP3LjRj+i6L7vP2WzuCT4zITBuYlU8jCGNdNdzFnfjekt6O5zBoghO8S+UAZpthu4qmNbr0e
Rjr3JI+oIm+zqCPYQI5JW1YVxIRzyQChtvQO2j7z7cPkVTQvR65gEHhg+PnkYi12jWmaPgYcuUPv
1pQv/GBLnUBgNyoBRCc5N7SJ+ECleKJ7CMYC7S4l+tvBFpJS0MJ6/HxCx2vINpW6FuZAUTz8wDJl
bR2XKoeW3d7U5zd8s/3uA+2kW74jbayR7zDWc7YwbyNpls1V/NoSokgnNp7vRGIzvJDrsXQy6850
zvnQVYuQRYYjcEOE0V18dIQ8/moSOrxO4GypGmPpl99nJkKjx71drBC0zhLD828PHr6W+JVwhUn6
n1l2XWivN/mpTP3l+gR+ZnDxto15gCNbq/dbzh10LdhNpUVIkwZNieg8x0NU80S+WR/wpnts+gHR
eNvFgX0xXu1lMCSczygB9t3KXoh+2xUtjcJpPYcfBlrBwQt940R2TvfBcoT0ojm3uEGEyAAxW0FH
iKdPIO2JbgXmL3TgdEs2EYO5S4zV3N72XoqBJfGnUQkZpRFvH3XolDg7qoPY9f5aPaWxJMaVvjT8
7ALCbhhuioWO5b/fWtd5Ga22kv5wAzWCZ4OosrQShu4G+MulXzUz68IRXmSN1KyvtQsJuOMUy9yu
ikP61zg3fu6xrxfmLEW0s/XHRUNO+f/2s8GjVW35EAXLbocVM4eXxgCt3YqITXNdwQ2llNlOYFOM
/iyY77vKqU511dSyjl6bw4FS2Y8lVY9gGXd6nW58nMAkkOsE2tvs4EHa9GuNwD82cft0vFYB97to
75UJgL7R9bxDExoeqw/PHUNMDUCrDfHozibOrUaAsfuZ/q7P5p/b6BSGffxBPToVQf6zuQWuaiP2
yHImcQ1MXFqx0aV/HTL1JwhGQkxdeztBI4MF78BVAxCXnp6xZxqKxwchibRrNbtvbsi+t0oOJICw
aCS5JuxVhcJr2jsIiRtaOwuq92vpGxVDEr2C7JNDFZyx0CFPGXLCZ14YbtdBu/Pqn1GziXG7DFYZ
+w0mLKo9PchhFSVCQRD4HVdkqaG0Egb5FmErsdJBwNt79jL3Oi4NaWu8lClomJ3o36fV9+IIVfre
0cNu5ygJVTBUKn+XNy6aod5E28+wxUr+WWmBAcA0ya7Iec+L9xaw2iYCPxIkgW4MGwiGXmQM1GHb
pUd75lAtctDBk9U0I++VqZL9Ta6WV6OrUOVNr61mB7VQPdsupOJO9ODOkecAX/DumdKoJVOvGL6C
ty/jV9rKO6HDY7CP99Jc/LdXbk4uJFL1+rVNMXYH4kstJLxCqcDBpxo5JUISxYfY+GH78g11BFLF
JA/PR56SBDu2UW9FdPYSqo+iGpQuOmGOQjznX/BdCdeK80/m5XUP6MRsu7PbNo3vd+Sb5/ZQDx3F
PgESZklwhjnDeZzbJwPLx94fMMmXtmjkFFnMlNZiMqUecicXpFosHwBRPC3FGvvFQYSnlQ7Rqxle
gMRvJkmp4hMRdxOXrGFG4Io8PqVFEptGOU7qZxhqcwAb+bQEZbLlab0w7krFhrcbGm8Vre38GnmA
0H0oV+iK+EN5HTgurfLPEDWRj919jtQV+WEMO4uSj9YKiW2LSBu/arUR8qg6eVpLuBffkjg74L++
2C7AWg0qaRaTJbOsw1Ru1Ck9rrj6IajF+nQVs/DZFFfIsgeW2AgOMJr9k4ZKBBmgMHtJMzYAB8+n
i8xv0peV8W9edLx1YenvSgFXA+Z5L5lhwO3LdJGy65ZeBzoVPNDgj27danw2piQu1fI1RHXt36d3
P36PN5r74MKfkReL4MKcOlTyiouQfbNFjfIXOL0N4m0dfxXRSjlpqzNqShL9Puz29tNrdPT8+Gta
52PUfTlbFUuDsI9575gYI1KyWLgj3h4/liZFCmNh0zEV8XamRbQnyjAGIKlfqAOYnmyEq08g4LkV
iLsmBoDP2XH5TPDYNuJcpTjgfopPez2NM/j1jpRs684YQtxQ15ZDw9Yfj8d+NlrTOwyyzyCJzVTy
M1s1oP7XnEZXHc05ss/lPgzw+bHYNGRxP2wI5tXK59ukBYkps36pWfwGBZxqVCbu+6EnyoLx8uBc
13npHpdgZ/OjkoFx6m2gPUXU4UpulRTJUeyTPDFnkqrg2Rea/X8e1Z8H5VRJN3udVDvuDBcIBkIr
IISv4BSmdss8Sr1x6zZUdG4jMmVCadhnoMueUC7/fL6Y2l0qyOoRvDmGy/Tkjqoj6SQDzOmLKODQ
bFCh1rDtH9gPtf365M1aOb5QcITSo+QqmHu9w2XcPDdaMYWcnY7I9BUxkTmKiZIN6tBElzxHumoG
xc2aU1wTqm4riUwUUzqzA54C1rUET3W6F8yxei4wn0EHFkoU3pFnsZfRAzi/oMedvvu7cME3HuVn
ZbH15okW3P0tXT7swqVKot16xX7lo/XmdUBOFGBo6d/U9GEBWqVSnB93F6OkyNwXk36J0G02dzza
S+U0k3iX674oInk4jDTVQCPEmC5elEBmj+nPqW1/gAQT4PoZBF0FA0j0wNblcenGMC1f3urd/4dz
rEJM6HBIwfnjdEk/xdGHoY8/Du8v1BTJdxEFQf3IwjFMHE3qvsU6V8seqssXbYCC3Z20cLVpf6xd
uDc6SHmMj4h2hGLEMEUNQG/GYWvPtT30lDdEagzrqF1Fw/i4suhWJqvF4UQX32Is6Ia+3xs7EH/m
6fiwjZaIqrRE5aMKex5YlbFh/DNAre9peAEN582ANGfy9T65Mm1s4ofeKn+t9btU0LbDi3OVjouE
osBmAlJ7wZ65+84sVdYWxVFl5DCLAdszZX0ewvSVZbb0LCLW0UvKhcDLMzyU+0RbYHVEwV2yNTvQ
E2K8I5tXvJfrfqfWrf90uLVGRCiGz2aQw0UPkNBq288zQZPCbaULHLFtV7jXEeR7440NWtRJ11vt
vtSFsUuzvOXV5bMubQkAKf5Qx02sY+NYi6gAAb3vT6VY8lLbm2z+bY81VL1b1zgBX6wJ1SpWIB6R
sFMVPs9vkUtVam8wW7c4TRdGm9grHzaBF1hYqYGznuHUi/fg7huCQXm44yiFYCevhGHWwJwr2SrW
wzzZtrtQYf7EvVRqP07al7jfGB1rujnUt62/CfXeK1UO+0bLXVpkJjvmIviVzbm4O+/RjexSsXdC
xGZqVuJ43TGgos7OkoTvRMfSu0FEismLqxrho2+WXtiX2ViCb5IdRbzzrgKluBrhRPf9Cro0zLvY
+edGCxF4BBagipBiI3qRCxQKmmIMkB4OZDBVP8HDQE0rI/lX1pt5CRQ8b4QtNzb6i0jl4qgdxcpS
hKtBh0gN/SbeGurEPF4Omvl4Lbsnt7HkhZLyp/2M5kcM0AICltGwXIdXX8oH5PdjEk67gNkjuSw6
Dqru/NDz5cs9Z5vYzUxnC89Svyb9feQoaM7x7Mg5gkKRIhqa6rrI8/tP4uZPpFl5KgqjxI8dShHq
J3zKPOb6HGRdgaHb3KKufDig673TXpUwnAeYp/yoCv8WNFebCj3sdoOtKWUJwlkEiVbh7IkF3wPb
3ta+sXCPkbMpRwj3myQVlKUugMvLOdims1yPc8d/yL8arS6ZapwpDcOkTKYrn72h9gxG59kqDTl8
JJfG0+5e+cllmfLPOu2G7MbXv2swuPB6tO2DF54m/+aC5GPwPchcsHyUJ8GHsXghiyuZ010cwbt1
QjxP6xsOuJ/8IFZv5P5kl5bT9cgbCProlLOmnyqYwReqXWF07R/mgtICWcVvfE/8aMAUkqTH8Vv9
qpxoHRHTOsLBhhxsyxe20d4zPELhG53lTzkX9sYpUFLEYzpMPeHWE/SYTkaTz6FC4adxtFbg1JTx
JVGk8imegb5KBY6O6iIoXTaPxzGnX+Qndz2QEWBBAY7DF8ZHglNGig9kkVp0lpNlFs2PXKkAj9f9
lGAoCUftJZe9Q1zB0cKzP83FS/KcxmAp4mxHGwK4iktjybgU7OMqUR3u12bfK6cKfIDCSjrGW6cN
O1Hx8J+iwMLHvYRrWtLB8pg9LkIVn8bbBd+d8Zc4qGBbSb8qQq26go8HPpVOySjT14y00Jb9x8ln
c9rb8dF8yeCxjNtGnFi1RGd24O8F7yY9esPyyW11aHe3yCnZ0D3QlXdrKfdeRUrlrBhTlGPPe48F
NpMokiLP6TMq5YDYKFAcqs941EgBiPe44JZ7eFrNroGtOavM1UUdyPhgQuw9XA4WrH21AWM64ZnW
QLey0TpuMMoKMOZARcqaABs2iP3r4bqVZsssL34mbLAZOq0Cf3V9f7vr/iXt4f9s8f/0c1+WV7Gt
TnjFecZ+8ak9y4ntl87AZSPqVqXELz3le9lAG2o16IYjmWb+XNinpdg1b9sWsOCOciu7oePh5zj/
q1wGrHWz792Ot1f4BAYO8t7LKRW/ZWriFjqXt36NTxeKie2dUcsIGmGnR44FAoST0ali4f0HveCz
C7BTt9yaNmVx35iFgFTMGnItyFNmSX/j3bzN1OEOIBYRAYvPHU2FNjbAUAypCvRlS80UacOOEOus
83t54kvqvoZnrjf+A2N8n9gAhgsnPJD/ytdw96n5HWbLtG40P6tUcXeUsmrYSTO5KfZ0j07u2Vbg
QLEQRhdPdPyCiS8K0itba/WnB+TRIUfLfMqvVLCp6/PoHSlGu82EiFCHOMaKimJe6qGgewfBINVf
We+Nxh9twx0S3HsS074Lhhjiq5BbsyusuIzm1aPk7L9gS6X0MhV6m2xgXEqlt7H3y67G+FoZ9T2w
U68mvvow2SxdSP+QXDg8uMXtpc6b/htJ6cOR9XcMAC4VeOAB1XM8s9vWNVpMXWCl2hQJQUnwm8jX
rozhr39xkrdUs+YnKzYp2QAVTTqNBuAM5FQvnaV21ztHGIl61M1y0DT27AlXBuhDnT1S3zLaalFM
tJqSm9dsfwTFfvQaogVj1coMprxVJtIXP5lBTnOtg8Lc2oKqhx7c0YHb1QAw2SMbb4qZqWjGSf9x
CeIlQqF2T8By0ui2jTdXW9jiL17PiRnPnxWwJSNhObBnW129lfW3M/Hd1UjxJBvaRu2XE9IENu+/
5n2XDEO52yXE+2+qGH0gxkU76Wgto+mHPwm3eup5xhQdOZyqXDJZqlDXElUKeGtvO3QdIV3CD81C
Vl3tooAD2bUrp4Z+Y+oDB6IdFsrPPpCZUXmmMCjDERsrFsR9iTeIKVYTrlCAeBJMTP04oEzTKwZ6
Nh7BAr0/QnYpkjeu29/E3PpgMckAUCrV+JZ0Rj0/SgtM+uJOwtKjGqomyQyk7ERHD6H0XTT3E7dI
WXqlZ9O1snFntPbeaWhUnrMSx4EFFctfQE9wMiMQS26ld41fVZF9+Ci7G7AykHhvHaa9RNkUZexM
oKtaWAIfbE8XlHGf2bHYnqVJ+Bpr78HQ6Q+HJb1aQegVNcMI5ZnNeZaJ5A0LqLaYY/SKhME8gRnR
GwIhrYML8qXIdZeH9gv/PVhFo4ofVno2H354vgNNtC7r9gJC2MdkH37kijKxaKIQ+ZAZe/uhp6yT
1Jr9+qF2ssgaPjbd/oyCBhKpqG2F5jcXx00p2xl8rV0IUaAUXSsGb5IJI5FEbc671kE8/XIB+L0Y
tvRDm3e0bkKCp8+Zy6B6uhyZJ47PT6BIxnWdSCTHfkU8h7HloD9+uv5xyw6VXc3JKPXxUag+lHoJ
RagbbUfxIU3om8IMDgzJojTv9l4K0u3sVRIwDWN9QqMsQYaKEI/bEnzFxRq3+jAC3vdEvfetFLZa
Uleyr/qlBjyrgzyGZYl27ZP4DuNpoBh8nVCZlinZUcZ9+PeUmiRY/FXDA23P3iNBGzuNyiTnQMZ0
glEwIXbFbOQrJLJHDFCifGp57k63Oi6PD/yBsUc+C00wxwjCAFQvAw4AHxNxicXCxQdP3UhmfcnN
wCeMP+cIqC8R9/z8bY4Or7ski99mDRGqhwRDhFDa16iHhq4O/RLuOQt+KSGCaOSXN7OjYremmolS
04I6pHwKRCZ9jBfuutkUQ2QOAlUgIsBO1pwCfxtkyuzjcjA09SXaXRSEqnvBTKF/A3nm3UXrZpGf
OGJepGEsCRwqnWjL9digj0pRGDKlVJwGFndm4s30yjiEKeeao5I6evbi7b9LfawdpwsvtAzc4cXn
ZobMBjkv3gBjhXFBzxoAxMyeZ3Mqv1RTkGgmcg6bNz0PwrnhtySEyGmNK7vXh2FLxVoJTQQZ9CM+
oDo9wkYuWlKLOGHucsyupqudb/hwU3pUu85WJAwfIvoUPKlcoeRqCiPM+MIpLQeLLDlIq8rfQh09
eDB9pGGpxJ/xca6x/U1LOTrOIdbA+fu9379Y4N4zo0l04qOx9rgK+yZH107GoNfAQA30wTpqr0JI
fuAiFc3bqukZ62NwYjznWCxT/8c89NapthUPf33P+IhnOVsy/8AKlmlFzcQ4xN+EOzBFxrdqWdxF
vT895pdFRuB9LtYPdWSpNthtrFCM7ETVu5rcI3px8EpWRkv2nXMyP3WiT0Yr16vHdJDnFKsbd4gt
Fx3dySaRnWEWb7ZusWlqiPxHoMziwGIN4nAPBzI4pUvD5E+BUDknk5x2YfDQls647yeuPcJe7iLC
d5ogDXmTEWI6le0Gc8izntOjDLKJcE7sqxtELLPqJhE1oM/+Y1K89gWxyVcst/LINP/Zas49neLk
tET3nDtOimfPzZp3YDkwcppw37YQGxpdyOZ0psS5Wv2/lM8O6PZR/aMEbWkFVzx4H2Jb58vXV8+F
0JaYdiUdR8DtfL8yjcgmPU6jEp9H2TgkI3coFAU3RaoV/oekKw2Ty1R0/YbdxBz1YUvTO+8Ok5qW
c5RwP7LfP1IyPg/8O7/QD/DQfyvAkdb+zwoaJOkGyyEeF/147IKTAOW+6xO+vBQxAM2e5COHAv0Q
3ieysYMrSwYtAPFz4uFmc/NOpa/UotAswXNykHIffeRN0YCoNFrcotuLNmMekhOwJAM9LV7LCO3B
lJ6exgDkRokUSnFTUMQfteGGJ6YZepQXBz/KH94SEwm4UCAFZkHaiaX5x/ThWIEPoJiyr06nkcXf
kHNZxmrC5VGAV0odjLixTxmDpHsfug+41Q3++8nGCfmubK9VsADzAv2QgdJVv6OJ91XSaBpIJ3E7
uDDCkXT5QZW/ajL3c+eFbeXpldm8LzIlQECgV0IQe6eyoC3sJZTnOvEVHeVKIpBiRlRGIdGcLVHQ
5A0s0lGBQNU3+JDaDm73BBrrNNKtwCIq3M8raC84u25g5amq7D4VLj4ywUygdecsJJ922EnTjcya
SEg7PYegc3hLKUr8mvwrnIhkLdiQWGOs/UHDUroLpp45iEHzSAUpTMUrqxQ+FLS77Pt0S/yYEEOX
aT2kBe80XHrV/iEv/g2CMU7pkYj9LuTtM5/7xeElTDd6Ov3HqMATOuWopPGL9EtCQM4C7Z5FLrbQ
Z5sm3EQOnc4Icg18DJMx3Ws8gFcN7vuyf0A9ov7PVzPJZcUHbWaskUGmVyLjzWoVhDVXVjMPxKfR
6vX6SjYWjQGuObuSGKuBY+S/wcoMUcubycODRKJyDwye97OydYyO0W7nwMbUmMFGywW0YLW+Orcg
qExd/rab+kILWfZLPdjaFVrm7hz0LYTIE3HafjdJVDHI7xvvkpxPFDsmj1NCOixmJOvofi7a/Omj
1/It7gNnxz7rWezFRibfWye+0TuiSmrxjJhyMPxIuaK2Axdlol2LqSHm5LyP51D6aKZeRehUoEKJ
J8LQZqugFYlSfdX7UWYX73ggorgcIYkaCsOurKA0Q307kPvWTgMiJrYRkAl+IIHF7BMy8eaqDGw9
Owh1qtBG3a6f+MQ9ND/Wl9IoOL1Vwm0+OKXrmRb6ebmBvHNg7K0o+y57DI54E/prEbrheZTCbgwn
Ter9xi4TUoF54UIi3W9sydzWjG0EWPpBbEhGIVoYpHE2giJlf3QJCg96eq0mHV+H6FokDgPUmApe
Gvd0agQ0vH8s/787/2XmztmfVJhDZZyeKXN196K0n47J98Nwnn32rWxds/lpEPb+ImlNptPMOevl
1GwtlbjaUi6JtM0ijyA8WyjIr+KB9AsxrF6bmlRFG2bripaWmIk9L5YzKJ5Jrg+WzI1GjN42Dy4w
oSYem1pZPy8e+9wKNweQHDeSgQtWgoiatW8r8mqDv5+VwrEbBtlxuaJAZMky5/Gyo9vUkxCynZo8
s9v9Bum1m2rm+DasXmieA11B00C7WIUStUpkIvhtEUzuANh257RCLQg1MonJV2xjW/AuDd15Gnn6
uqaM3qlTZvTW0DryVoDRrHvnjfkAIIA0DgIR9INTU6qUvtvC/rfdKKKCIwOWY0JTn3Qcwowjs+0P
0OMNd+i7REaUhzTCQxQMHntooBV2VECHMXxay7Z8lFhbJPTl4F2HYhMAV9Mth7GDN5eaeMOEJbCZ
pT5MI6//izFGI17NhTHTswCj/p99XWtAdLBXIUX5acAlubmKNFYf2L9qWrECV6vaOuZDSgcp9RIE
jjv//rUH20P0RwYvVYulgXewYHl5G+ahr9ZJKstdj5ueQF4MS2bCnGkj+kpS+jtF35jSaT480MP/
mx/uQN7KhUUnQmE8FMaVaiTf8TRCovNHLE/nSqNJo5XbB/FZBwLlywF18xWCf4khdogE1L4coid6
9OW9JB0ib0MGQmh2W36XJJGZMVvG+6y18q/oPNlVdZKgaL2zHbrU06KmPBdWy22wY0v41QeXB3et
pHQpAVIFpf6et1wkyBwfSMCaBlAEKcyhl/7N/FoY0xe/i5mDUaKoxD2dfiKL6K6jDQ/xiScMDUoY
06NWzfT7JzyvcSfadbZXgsPYaKgWh7XCI/tYVMIFPDfs0mzToSOrSx7eSbXB4DJvBkmkvfO1ouap
9B3W2HHByikh+OP5Q3SBG4KHbboKpJ9TicdeU6UtKj0lmEIgSByGxrZzHlGElgSeLkR+Z+K3phle
YvvaHryIqHMwGCW7l5ODmWnWeZlxOFJaS/FTVWXnRs36A1FhGUHbEeQCMRshtxU907G6eo/oS/QP
yY0piVuy+4QzPhKEExCr+bDBjwdIWks3PDRL44F3wkQDLyR/Uwgxi116eIOFD9Z4/mAoIemoWDh6
EtbtHxrYMbZ+wAaf7AsS3ghEJ121FGvOltO+hLxjL1bo05HQw9NVSVzZhIgMJT+4SEaQPqTs/4cY
EIITS9qhE5lcCtL8TSE7dHQ4xWrO8JbwJu6B8c4i670XDcOZMEn0RDMolshys0zrFJarB5oki16B
PaRB8QMS6hDNygshDUJnBQ6fvx3izo4U6NeP4ab6/JfDRhTZLh6OQxHcSuvGjiEl8qVhYTodjc9p
E/QePTQsBzCOy56Yj82j1SCJyZfe+R/xNZSDrVtSxGdXzCJIDEbWyvbDgqMLaQEy4T1ar+/a0gTV
v+OSnoKf4Qux57gDWoSFZpHcz1aNcwLYWgTii2mNIabsS5Z96B4a8K166ReKExwpkVlsi46nLv5H
GmCaDqY9nOeWOekVfHj7b3yEdUAjVFdzsp8id7mKacNicQNbZdIIqZ5DmtvpYhGRTvHoFEPm4X1V
ABzeOikxWv9729bnGy3ftTFpY74YMO2LgWD9+LC8+kaCb8Mq1pG/beJAwXphFqWhHGMOLz440f0Y
71nWFR0xqvYlhpBv2px6TEHRuBaCpOdl7c3isjsHWHAneojvjSKySzXdWW1YkCWJPI3K2tQFKR4j
baeQyKh4jNjN841/O4hsbdgCUpERqGnVjdyyN3qmeIz2gBftBseq+t/Nei9fXmfL0CSrMmxSo9ip
4JVsHwhmJUnH6k499PPvUQWVyxPROXf93TGa40WooNvWJPfWIdpk5SAotJ84k0q0gM6hYOz3+KUy
yQX/OZu7SNseCiR8BTlKLApgrGBTgtCQMlvCRC4gnIZaCLN0XXKvyA5A+CscNwyNuTEKl6/YZe1b
XlO6k/JUGCX6XeAt1AUtAcv0oJ/yH0IqDvrsUbsWQGnhPGjBmsbQfA8a7Sjg1tr44s5aCJtD5kl0
VJKOBkTJhjQm6OWXlT69PrZ07AtyxLJOjYIhQC6sF5roaBXWzkSHeI1IuPrGAzFNjdh5EK7s2LDF
sRUMpqhIeOOWh3uS+BSkqiuG/5JaKiowkjTeqL7QeEvrWqJ0/c4Tz+rbJ/SRCnE3l1Hj/AJfr7yZ
SkrW2gNOiA7kx0HWePc3F4dfBwwdmlbVyH3QBb/iw81epx3ZYCCzEKqPJlyLW+ILVJ3G9qTmBUlq
bD4dVtgAwRaZrpDa3jX9sOuTrwjj7oDPmSsTXbklLdhL0Ni2dNbx34a+Uo6/AztNdM9eSVydshY8
XY71UW5AGMd15nzby47oX8at0416W38S05DIw/nKokxMoN91BSAe3CW9l/qlDOpXNGXKii+0JOGl
7c7ONs1dBeNLF1AD5HBZVI+1hms9YNO9/o4FHeNDfSkcz6XVuHGGV8DlQNjPoWFPJr8XrHzCh1ZN
kS44FLar32JaEZJGgK21dJjy9z/Oy6XlnXdaXL2/HtNgs/zBO0sP8Wz0rirCiJB16hGpKehQaeUX
+GMMi+YZgire+xBhAioIFiuOg6aOfiX647dLDf7rcHU6+068ASXufvL7oxvnKFDEaEH+ynhRC60+
eUajVpU/A9oWjQJ134grrFDWci/w5aP2JNcSm7UjWRg3yubQFTS33K8YslYu4fMLqzDZPIX+Xjqn
yQAZffGHQ9GYxqd+v6x88S8mY1JFVDUoWIHojMbqbf5m3/ygXCN/70ujOFWnAJM4VhebMQ7lZ2E/
Ys6wBiDOz5bBNgcvnD6EYPDp1znpdfygYdI6lSVLXrNl3unycPh+5qWDSffsnPOFzggAJB1GsX6K
Kd+KZtMKk0qI5wwBGcrekoQBCZXc/HXdUdeeMiP2WzowrHx3AqoXL46nn7OTHSlYF1xgtuwez2Db
5X6gWYwJ0tyX0vSqohNyXVmqgAZ+7JoaEAYjYCVoPvPsbHeuOV8Rx2oqrmxIaTluur2+CDjFXGJi
IDKWmF5bM14F6usaFh+G+J6DPF9i2olUqAGSHTe89Ra74IYhNOZQ/WA1YH3UbaxOIoCuATqUAXbU
4fkYqGGyk9XgIRERem9ql9Shmyng6glM5h9NWKsreT4BgWw0so8RFsuyC/rFcgWQrsh1PiLG6QWG
7gA+LIAbMDYvyB92eutUDtuUgpG/ApxU4T0t35vUdrD6IEKH3Hl3RNmH/6ZHHDj3z5mfAyWqREp2
eWF/Ch0Vfet4eeJgq2U7GLdl927qPQvLOrpyyWf2s8pu4KqQKGjga8MaP5iWlB32X/nclgtkcE5g
Z3reG+9ELFgQj+bq2zCFu6swe9jXY+tnbYX6Wba60QxtzNhFSoMsqltKHmOhiOHGo3dq6n2u6iZE
g6WY9e3EDKfDGnAZbnpVdlJ5PsBYPCM+TYcTud7tmrUb+Q7J/6lqcIRgfrprnNjB8D4YMX9T7EbZ
cffgRwRgDuQhu+5y1kCAVkQurPvHbGF+ld/6px/l1lYqOX+w/aWSwzEdtnz86Bi0v5XYyWoPkIf0
kXz5dUM5Zp9Vo/QtnB0Y4lV8qaqoJKesjIbw2DI5Y5gVQnFJfneHecHuZG348CeQURBa8jkLUaFg
4IzO3Y4sMomMQPRCpCn9SSQXx7zQtZIqeRDiCIrOH7xsfKLCnJ1YGNBarWTYp1VF5fRnOD2ECkl/
7tfd9BKLJ+wQ/cFBhPFo91KzeDhVVCLG9HVKTuCoZ2Xl9otBTCrkrNasl9A1bCskxAE9egQJ/Wxk
ptCgMVZT+pX4IQhkjXXLXq1T/2PsMmpiezh+EfeL0Dd5VO04nB216sPxD1IP3rjHH/C1YDZv6FRM
V2Nr9yoGl/Nr20wYgJDGqJLvUxjF6seidXR90qiaFl5Jbx2WM60o/RXgVyLPW8gs/NYxYdqZ/5DK
5vrDa/FZJolK+wJcB4PtvRSPykOkfwQVXkGxW2HT5q/If3ClkGOP+d+1RbadJ34D27zWHGWUmS0J
SSUCjfP8AfV+rP9PuDEB3i/XRrEA9Ng8nYojfm2vq6VollBZn644dKC2161h1TzBOdR3lDSF1zqP
eZiymx82rrbv6UfbgdBmAkkMc9HBBX92fc3SRn15Jwy6mny5ETMiAs+9oqn/+M4+WK0Sgdbb6nJQ
Z07GLIgBo3RZbTxjmhW9EFCx7plQw0K/LnenuRqQPM1Lmc1ijSJmnACSRfKNlqkRkntxfr/WBkja
tmP6cXLdTg03bCnEahMoaEi8dd5JgRftBYpPUBrEcMQhGC36kgjQ1r9gUr4ra++NH5mGltZ/E2xd
amK1dU6bQpuQ+01fBKJN1V/km6dzZuOjoZMo9vLQ3nf16+I+8+cWmzCCGiCT8NAc1HlkmOUVp5uz
83XZr45kthXRxYbNfEuYHGyXDeDh+YdHYNWUKvyQadLluD0kVEem0JFZQWoSqkae8oqIHuTpJLjv
alURF+W7MtN7Y5yCcWGOt+5/8YCjeOf3zaHUh6/4VAgKeqkimJwivCekaS4x/M91W74G95qXbPXy
GE3zIYYR6TsnqGxhR8FvbEMKFdwd984exvA+cIt6IZkwDFbE9F6BK2A7lTpf5ToAg/u0/BRvSgWW
szw7BQP0+9vX7SOxtj2AQAcg+posSEfVWfy6iAFHoLdRCr3/Dh1eMUD4XFyCHELqs1aBl5TsUI8x
RZi8sBMnHrUUgv5N4Hqx3AUayh7TGSM8XZkFHkh4s6Sahg4sYIsPOBhGqaNdrj3icvrEVEStWFht
p2a2kUc3tgPRsbmvzyzd1vuTNJGhQKptJOws6N1toa1U+Ragaqv106xRGwzUsCxCvwjbtEB81dQA
y3RxBWt7E3juCPk9dq94frmSpabzoENZzOtYd1vOETR69Fb+qP07NQY/JpdkMlo/KcoaCO6HsZCA
xnE0Yh/Awmaq1x0AQDbwwfCqRqoyPn5pVF1IClvoug+JXVRgKoAqr9b9X8d1DRbtCWb1soade0Pg
Bd+mghCDsoXjygKT9TROw+LRXmRgALQ03cEaO+JldUFS2yE+1EkvftGCiHiJAHZQUiqpKHvbO9YJ
odKJGZWb5iQ1lqXhqRVu9FqCozS8tc/9UDlbjKM6ljds3tLsuc58fJHkNB0qbXqgHj6mXIQIgs2i
INWm1odpZ7aiu8RYnNOEKdIDYJxEQNJwa87Zv/ONuBjxbVedkv8Z/9vIXu3I6FWn3pdsBFhAPpZb
o08bq7WLFiyi+ChQnL/qACLrxEqHg1Gd4F25mHzmO08tFU0QJNb/intzPPaUmVOx6ZopP7vmij7P
/D877KrAuURahBmLCpkx6+ZvgrFSwat5wJZTedZVyL7w/MaKiSYdllt5nX5+AK9x8LjWLkXrqIiH
zm4ffjHdFRnYGnaHGELKhYpjDZJywvlKRI7PQ8Idrzq7XpoDiI18r3KKtbvM0UBsKXDJSp9zESa8
AXobpZkG2uLeYWz2tASv2HmqrcQRyT4QS2gauAEKt9Uqz2xDzfgJzWySR65DjM2Z7GlxlgpX4Pa6
BSx0xTSRYl8KW/h69FA46sWAeHFX3QduVl0tOs23nxG+pmXS7XGYk5mDgJ2Ue4XPMiem92pHegv/
jnT1P8g0ffkaBQ7rLZKyibYwCB4XjDqnmOKcQF43jyArZOOUfUXse9yDfZ29p6I3QH7PqzBjw1Vs
sQF18oU8RG9n4jF6vvzjPxl17d8CuVRQQfmBZ9FAqSaiTfGVhIxJVYhvclMpcERECFkShV0f8LwA
DSsFNskpxhoO2SKLH1w9K/3Fs8ZbvN0dEzKvOOYq1e6+j5dNmEy0c2V2gau9SF6Bi4EvTQW3qypF
tK3cvP2z9byFFk5WvPcJEtZ+8p0OhXboAo1epgXjmgAo2P6gTJ3UPUUsXjYZ+Vubw1tiLiLTWPJT
4X9RkXe2WvO2TbkQvKFmigQWarnhPZSbSgaGjq0Zp1fDYrj5Vk8fe3gp9bjDt5N5W1sWMLhOI+ag
rTSZcmtlUgIcdygGB6fUBA3pumh2dKg2QyDMVovE+09ZXbJ46ecinP7SkgBVzHMrkIgSzI7iyv9u
OHsNJp4OSGI7nIEk0mH8NHJu+PJ7YGp1jr/i1qmBvgP39gEFELP+7Y1HH3T9XIQHh6u07PdhobbR
LT+AktnPAodiJ/UnRK9UoUNV+a5WiGgkO+SEAgC2zDFmL0z+JKfP0o5+oEBVjyM3eiMT5fVj3UT+
QOO2Pz42d0/5V7PQgM3nmoc2wQXNvowWQcMlMnTVus2KxOcX/bpZSYPwZpo3isvbhDV1e/17XeRj
n0l0wuNxpzhf7kYcdy2WsjU3+ciz2yp5ebc+cKwz3u0jp5ZCmH7ca0Dh1TqQsKD5khs5IyehMUWo
uQDCaIa82jl82rLpCKjnM+yR3KIhNMNd9coRZMvDXOxABDDoa+WQzFUMXIT17Pi+8wIoNtgIagFq
6ZN2CH5ZzFE5yfL5eFgo2FWyX8F9VE+2YYZp9ja1onyl24tC6wSJUFNFSp5ms8hwjVHiNHfMt+Bc
3rIi82P6t+pgSL7K5uHXEblisDUMguDce8EeQMF3t1Ab4HrCB857/fNdQKefIvJU353TyuyZo22W
aFaVsqBhPRDEkCsfcjii+ylMelKfP4DzpOBPQAp1IzXXihkxDZ6RJnamCivBgCnUkH56wnRFPRMl
IXjbzekd+V3dhpPLqyFKJr4gn0TJKHZ5hJ6JUrJI1n4XULQvwoIC66u5uxsNrtw0LbqmJ95QHcMS
GwESiJzEBEkKE71xRfBrnt3ie60+2hO5XlkqwCV40f17IdccE3Q0GBxnfo1AOxxp9R8bJFRgJpTH
kWb01G0HI47WgUwJ/kox9g9l+U7YclntlawFfEAoPX73yt1EgFE4pNqlsZtFrOmoMyuRXDsx0WKt
xvMgybx8yYaIDh+Kyylrzr+sBAGQ/Xm8dXUoS+FNJecSbrFjnZ0ihMMa8uJudL/YrOyr6bAhOjv2
Q+b751m9fQT/Y7azaRC+oL3Q71zspdtfhVtK9vJYnmLpQ/0otrD5tZhm1zMtA1ikdwV6prfqsBlB
vA48NyOdsANPTmQ8JqdRe57q7Tsjv5lh/LV2tB7SqTj+8WanH1R5amgW5yQ4C8djqmPu1wcJYzSL
kSEI+DxnYhVWKApjXYFf8dgUZ+FgTcVZ/g9/bpfmbw6JJkggiNNC3Og33XiBEx88qoiDeJAwwXLE
lHPQVEWK3bmrnOAnxkyPmdvWZqiO+o6N2xzdNBuLwdod3SaxNenlvhFnLydXY6PBp+yqyrEzE+Hs
PNx/BjFwqyVSVPcJZ7Mr1myw3EEkS0vUkvJnOdPVsMidypLGWYwDon/fmnKN0v6+kg0AwXa+wu8H
KyPKbglPj2W5AQ4he0aXtQjhSHC8KcbbPAlzptSlENr70cIcDRbVHo1olHK5N2MNxRwRBatEXN/a
yja4C+M7XOq2NuDOq7hoBolWgJPLXssH9qCvl2XXGq1gsb+Mov+AcP9fbdlKgT6p9nbJY0enkxvd
H1V0cBSp04hdT9fszO3ghDqBgep0JOCB68UAXRP1NX6fkq2bYQ0y6zUvTnhAkiFnFF/FdQfZEGCU
4Q4LhnZNkl8wDj7Ltapq6UFlfbslGMzyM4xmrptAIG+engOUaJJYRyLog5T4sBmn50PK+ZNixv+a
bNRqdVrkd1sPf1f2APt3xB6amFvzXc8axRsoAawVfrizyphO+RPkJIeptIuwd1daWhXz/X2mcPsL
M6sIi0di67axOcGz3ExGe4eKlIHachIkyE8spk1fHkkr4NoavEJs91n/+0WsO/zyURNVYnBHoQJN
+ac7ITArG+96xSVqCimlZ27hN7EFpid//eXGzKkICDsYjYcj93/jPUuTjBYuTmI8krqwRjIvR9O/
aTexHBrd3aqFSLpd2xVbAjzBLUeTIUj/X1x2uyJi2hJ1fGhGgB/s26DZZ0ahuY61HGbmFTk105iF
RvYqCptoEeMnVJ5Dqh6brzBPaSEoHoMRBmNS4LhZLHcE1I+LEO8Gsd5KwISrff0eYHeIKtm9Fnec
9u/IcChnh7qfUEktn7vu9b+m6mxXeOtvgTaTrfnJqLysdijNY/WClo7REiSSRi76TqjpRluH/MjR
v8zz9asx9KDpCCdoM0I9Lw78oEK1T79cxZ3u2thhkPZ+2F+Cn48rFT8489bps+QHMN2YYcgMn1ct
xmylMzXvfGcNh66RUY62koJXW7RA7a+xLEbM08gi8EcwcZabKekVd1GfK3wp/lufooPUFjumEPfL
iUvMbVJHNabLgLYWTL15ZFQmU+BZOOk0faEDisl/f3MLwENP5Me21l1jueEWS/L0HalGBdZYrnXo
fF7nGYv0QeCuBgv//6DgH8y3R8djjqVcyvFMEwh2rymIIa02K02L5Wrz3aFficI8XaO86gCtnyfO
k3GiJc6Li2tiJjS2LTCqDsf7DOFNXCtIlGzTAmgiAW8MfkjkczUb0ng++NXFym2xA+VqlV5fBpH9
uUbYHShgQsb3anqV+KoJv6Rta75vjK7Sl1i/TCKRAlYr39n4lg3GSkGEVmqQmml5RA6VaN5S+93V
V+dOslrQ/p+yUHFQykwtbA68fotixqs/RANLdEk71niPxs3iK8ZSSGGPG++w0XEmxDFMARbPeZS/
TOOsUxy4vGy86bhMatMLtS68jdsPGE130yRr1TuZ0aJtSeX4MEIdLfliIzovS5zlEGag2+l4FBgb
jBXsAg4+K62XfKEDgbgzK5wQJXT8LfvdckPuFfbN1ffN0fWLc6r4xbvEnCDyRccLUDfvdvmpf8Ly
kmBg64YlWVr0G45mpVWG4KQNqSFZPcmeKRoLmmiykRL4yOa5e9kadDneK4LXnmhX3YTMwcpqLyh2
7MR4YoD6Q6fQLabzhXGHhFAXvkbaIvc4GY0pgC2t7+7gsHOR/gsFpQpj3vHWteiylp5VgT/ddJuN
6q8lcsL87ICHLrn+/AlSjkRiS75iCRsN2WA4Cw2tYt9AjYZot1e1jhLMK8rO4g8+g9/HMoxfvbIw
pz+P4xF+ccu8KGjLhfPbMHhFBZpWOzR9rnnYcIBvHX31cGpM6VVonYDJOGgRI1S2LytsByKg/vzv
t0cGquL4pXxUMsMrnHw1I0dfYMmw8I10sr1BP3lWpunsEeUqCBrpN/Z2Xsgpgx4r2Aa9DrXKnxnu
qHrKLlQuSnwCKHMUZT9i2awrHMOKRUum0m055+WuIqr8oW4epmkodU8pRaQ/llU2tcfPSansXoe8
jKsux+u+EwdDP7PI/a+s65y61FM8W2taHddy83GfM9PlDTA0kAWY6qB64fq77LJYko7EDkXO0AMV
zCF87+2+WMg4FAFTcIg/1IG09b1tdrBrGc5Xzxe9uEmt3S6UmVfSVxL7O8jLFKg5AAmNFvZL1yS0
NlSuwn2qWlvE/HZIhIoTHYe0YPuR9OivpupAX3sFy0kzSLSSYDghTHFbfuHypyt5eX+tc6CXxX9W
SxMCjDWxJdiEH10SsCOfbk1bEjSx6p9OnbW0oaPcXxG6EVFDzQZtKsYGaz7ZkGxL/0WmI03gxQrV
yvQOSesgP6melsQ3eJtSLSyGkepyWlZmPh3zqSlXETkaox7VXymXDV5/Wn3Ii4VPrfphEkQE001j
8p0rO9uIWz2JCA28YWPau77G9hAM7f7+OzSvRKwskjhHQsU2ssSqfYTJVSz9KvttaBK7ia1GMM24
XCcdRj2Ldxtm1uHNYcRx/ciKb4EGOe3d8dcpKUdTwjsNYJs0mMQJzRwlNmFPdV9sHiLzzkmpjfFx
q6afkUt8+7GaJDiX3KnRlQx2oKOVipMOCTbGF/MW66Fptngac+BzcUlhlwin+OKVXEbH2w9/iuhp
NXHrenR+rFITmZJ2lPLfBgAAsvVLFMc2BTR17kAF8PDtIkxIgSm/PA+pmzrAEHF838BeY/84UQtJ
dk5DKRZkWZeezAaPSMzMjlSB+w7hzDKzfdev6462jAs6yUUVgS3ee3rw0WX7+4dX05J3iPpf1B+G
JsgqMWRu4r1ncyRAj6dpMkzPCoECWNkpBV2TCBkVP4vjhlcduQEhXg+nnEutSoCsU5fg81/xnJkh
8pYgQnXlvFEVesnYDtr9Y8ysQZ6HO+7PizcGmgzwXPMWyLN+oaTBkYhMvf/uLL38bkY4pabN05KC
8KI/4Fa4MO7vCIEjslRWaiIct/In0Ehg0JLPk5sGpXnXV74kVy0Q6dpHZclnLOQFSmjG6xHvJnU0
MaiLZCPBAKrKE/Qfqx8akRCOx0lmqB8bY7CpNluunQ/NMKnG0bneyY3RXOUby4ZRb68CECxMZxf4
JHlUa5NdPr3kXpbNmcW7N9NAEYmcdCCefgRyxYcO2UEa4hxtXZddjiTEDdzPXkKc/c7K58mOPnLT
zkbJX4T47afABLSGpSRKnm+VuAwJ1Jvg1XADhsjuYBnL1ypK+SvEALwLTG+JK+sFV/O1F8oaaCPB
Dlv/yo416JCLUFdl2LqXxw46WzWSfo5t3CnZPBOpYBEU5Ye8wYDP2XR1QJnyL9JMF+t85ECtGghN
fvKuAdLmAi6faJt7bzwlV7v/NU+fu9cNZ9CH2N7kO3LVD6H3Nukib3kH/E+wMkWt45NQ0w+lrbin
5kT3TuBity5LnxBsaZvWrgR74nfO5QTCrulqKzAebUF2ARtE1fIoCD7dqUoYsjDWxYjJgIR/u4m1
mjepOuTLtr+0S5tcloP8YLQvT1OKThgSi+X/s0g3tYY5cRZiw9FoE0GZfrGmrWS5abkYyamRI9hi
2lx4cjJpH2wpAEIHHfRUxGocvu2j95wyOtD8X31DznyR0HEqt3MRP+kp7tJc6Gq8aR5oDtOVyY20
h3lim8OcvxP0Hea75ZnFO2KIF+gXarNs2aW21SzT7Nqd+MhDk30em7vtK1SxVeMFrf1zcVKPN8zL
ZdLtZJGXX7XUWMRdkYP53u3PQAlegFFff7ZGGyQsls12dbulFHspM9HcvHuXQd2Xkoct9pL716Je
WnHsXcmXXGDcs409NEtxKnjDlzY+JhPU09g3M1Ei76m3DIoNe6gh9aPrw4jGUcQAxZBVzMwbXVM5
D02c9WwfHio7BsCi+St2MGMLfS0oUHUiJ4UXIC0FL0/oAxAjgypvP/gQcBWFmy3NHTGr7iysbKnV
Hi4kObDKO3OZIPJPHtaSJNDBOOQSurU7kGJg8Tmt/zhW8yoxZiX1kMtBpImsfRySDXLzYtgLBE0O
zolRUJXgvjobYojpJWNOe5gJ6x9rnUH/jAg9AeBgwAK9QtdQh1j8dlsBRg1L1UYKQbtP4SZNTliM
0tBzNU/WmRYgUlMbk+ypq7+C2lBbRvcv3/btVxxNl4W9zsRd6TN2OhZ51lFiLg/RlVu6Eml2L1IA
uEw+mkmHuzEog7JC7osr7iO+VNmsv8yMVNQabKEqvCK3YYoZK03SM3NIy2i2SSjUyzYpLl1QO8EA
+lgZggV/5DQKdcaOnjvrW2/iXAtG9wB0pcm2fzbiPdm1Qzu/XkLk+GkBq1oLkm5QKA8r0DVSny5H
XJH5Jkqb1+SRPzZduq4syzmQNd6waUsmniQaZ7EOrVLvAIQt8Ira7xBBnZBQTOh9cYhUFNozzhqR
+IiAcWsXvoet1ikfrBDYhCKxt2Y1axgKN/7E0bgVWEuxnxam+E9nzu709rVoenGqPp/ivaODBSNb
dCV7FjJID6VWjyXQD86ffYHf1VdLI0MNvLg6T0OIvPGvfeUVcG62iTe6j1o6K1KbRogUXXvjnw0U
2tfEuBCTxUsgYyWcML2U69hnhDLAcXIHdIwHzvQ6n+QE6WRXUf58/1RtFXnDl0EGbI/RqtxLl+rF
iJLen/DekxhqwBuCS9Op0rWLrEM7S9GO26XYSzVM1B9C6MuPnRUn8smC+c0t/HlGrYsWDKwpHcnu
H6L6/v1PQ/RVf4eRiOE8Xl4Jf39kV/5v6r/l90Ssyuxni9bqdEuHMCmHm4/Qhra+7Kk6t/uQv3lh
4HoS9EUiqbpL/hhzM8xy7CTTwffvaDKdjq2Mk97f3An5QT4HqBgoV8MqcxgTT776wOJbmJ7y0W9P
jEQpNvROwH/NlBX3YZI0l8QDeHfISyo3yufazvEroeVvyG72fehNUYoMmt+Dxd5ZxWAQh0PCIpPs
Foa3Pg5ifw9/+UWxmqfZpRRZa516JKLYwuvsSadtHizdYslDBr8r5Di5vWLZCcjllv1yiZGF0lcX
EPZeAtuKa1cVeKGMxKlfSS5f7gPa/24iBzBbWl7Cy2R/UsCBx6bVJ9+weOuqfjFWf3bTU+neKTXW
Z2l0yoNFKd8OfMmhbpeho10IdFaiFWyjpzuPAi/LXDCY2SVlpIV3Gfqtna63fctdj7sarduJMDyk
4/eRtSgCXJ7rvkaEYQdMfTuvbVxNPf8/JBrC9PyXf9UTzbOrl6czsyGQYys2/0taLzTd+m3KBkHA
eNdznHTufJKAShZjJ8pJTEpOy4py4dy74SHS0mkRaKNJg19QUlHPYlvx9mWsBSAqiCmpHMV76qBx
SClKYvqBPmfUzIMIgrxDqzqTcWZqdiWWBekdpqvpr2ZB6S22PC7z+P6CVeNRca9MvKSffBVeMarB
xrcqJuRevrwDNOQ0Rzpa4buPAoFnCXECxCH6oE4cjKquSR1uzWHU22LLhjPDr8iKEQjJGQHaJ9G9
6yMOnSLtH8nqhC5xW/bA6XWkjnJIcmCiPKnDYfjXA76dCeZzAGAdz7CyPT9Mks4ccHNvOEyiL8k1
taTvu6zTGQtJtkgllekaWiBsOaZpxvce+7dVfy2Z20nhcxi6Kwp97MwvbV0klN6mwQHDA/Fufc40
iyS/qP8a/tIjLqmJ1stQSoYFSS7L0rcKey86/igIC2jmwZR1s6yz9Py8swfleE0KHvQ2i5b88K+A
OzG/3irC2j/qyJrIE5EaRvmhgVmUsAK43lVUgo3KPojeesCz7omOKaa/yi3Xsv2PXipn44DlOrHD
r88Wfy7uCKN4zhRsaftweq7sC/yYkJnnnd/N5ispcFe/G/kv0zM/5VQClJyW/cxRMEtrESrOd/50
GdB0cw3O/otIobi7dC0wWPwkrA/QEQxH8pitXMG6+MSnHitXRnXu8/HZqNR7SY1pIm9N89yuNOnM
BbukJ2zS6sjQ9pcRJJiZ3ECq2f6nMIVCUjsh0k7hF1VWvZc7tl5hZz+tWvSN9KSZF14p4HJOOGgR
y/oMnwGba2HEic61FNjVa+wqm3vfWC+ZU9CFaxteWdvvCDQhePQFzJGo147dar2q9RCbXabCNvWB
LQaPdCij3oFuvnW9nGbUqghk2EP1K/uaVyW241HYAzdpKU4akhPCvtdRqGSAX9oHWrjb8rsHorIp
x7X9rULOt3vHGAbvMWNNkzqI9yYZ99n/QPoTC/+rPESqOLwN4nZq6DkhL7d/yJqdHwRBmmejOc4y
uW1OhpRvlYG2oMJBiZwxCMlb1/h0GBC/O9d1X89opHlomYtZMtvPXMRT2djU8oGsRCvJpw4e9ld7
3ylz/l1GpU00rUzlhHze5UGmBMa1zZAf9MEvqq6qA/fBLl/HpWClzulR2bazvlIpKJAe/VEUyAcl
j8W0iv9JfcYLTGtKdJmscQgS7IIUKVtnqbxvUSbre4+sYq/euf8p7gINZaTbH44zYfkKgzJIrbqD
hnA/mlPxo5t5ZR4k5t8B6BxeLW/kvjVntYiLDgJNEa62kVProCz5/3Q4Jc/mL6yfl3oNO51QxrMY
Y2Bt8lo9aG+il1o0RfbHS+wnxAJb/1L/p0wf3XzSlDykB2rS0lrd/P0wydwmTKD3t6B6d2Uqua+R
bmcGkcujP5/uZsqQXKOGeZrF1pqx51adKVJdnT2GV4YdE4MO1R6IyWSIO1+6geVI4gxYJUQBxC6b
8TzQ0lgZo47iKoj5I543JryJFqgtWKPTq5jkCETqy0uRgTNMYoyQ+F6ac1Y143l9b8No2a/Ns7Az
madAUV1gpz800nqiXGpOFv8xXvW+QAIJYs4VszzgHaqLX9dQQg2oEF1/esMQzQpQqYpKBf5wlefF
F2Q88N3D4Ml9sDp6Wfk4ZsWF+DXOkR6SvdIFkQlKnA5JBmHUze1MZ0iewVBBAYz5quVpECeC5oVG
ac8yQDxm+YN4KfoH8J3ONXVn/eaoJccK8OJcOAzT5lnSHAW1r6fOugQ6vbvcZbFhkMOIuBALR9yv
oCYRPu0+JU3XCkZHKCr7Rg91oBaXOmfU5n8rESm9oC8KutlAtIsqenrwoRvo9SYu0FeGDC+p88UI
1n5P7Pz8HEb0lHN6d+zIxIjh80eCY88iNMdoy17fOTJ1OtV0XwcL3UuS1TvwH7yxkMoDj5dsQhEC
tol3s28hDvid+Fhfj9LCzhFbYHyAT/xNfLqnE7WaR0V8DN+dFZzZpSPL8++eTqvtOW08oiaR+nRJ
WwqUaf4aTOQaV2mN9D7quxUzULU7TqIl1BkcphcKoo2NMhOVectKbso6iH8zW81wW6mj861pYKDJ
iIT5zGb40AcX3qO0sjSVRqF+2zVZeBo0F8cTTmZwOCzoFbF0n+CQChFBsWOx5VaOs588HOZc8bYD
LOoRcFSknuZEP7CcNpzP3gFwHTKypdQu6lC0UPuSzq/EwkzvNEXGRG4kIXb70zvBhXqDQnJOJzf8
d4+P3GDpPdExK9a6ExoLDNAPRk3KcOW/iehpgQ/5trkcfOYLaKSKTZUXlH2KC745IGZtLI0a/zkr
DQP49HI+Ebim8YUA4asj+oCH0mCsKd+MDQxXimD7w8Xy0MavcV/oQV8vhMJxE3ESft6llmba5t04
NmnuWDKTm9PEYZPLGpXtrd1EZN3mlmfvI6ApviJJseP3UX0QExsTPbD26yiHWoehtzKrMSfpJckw
Hs6+jL8htX0kvspNxiNXXHsAb60srlKzqCwrTb5HNRWTxPTseTW3c7oBqTqAlQQeVzfl/zTojNY0
xiWLKEvjCjpaJro+C7w+3Nlvd3oXyQGh43Vj5uDHddWgO2vgXFeiNqWWSUMKjRyN+RNZZa6OGjSr
b1ZsflPY+bK7FsrPhaA9beafbR3QGjPcIa0sphNlgGvVUlqBHR/HSuIm+lkZWSohEo4HcM1Yuypg
A+PYadh6YxjFrnYvc7klAvqcoeEa6T3srqu+wyv4Q8a0Pmea+NdoWxDHHCpx2oiAFvBLjrxs3B4m
/bLJzVqvPSdUmZYVJCYeqxPVh8pzdxwkqmK5saFPK4nHGnW0PPfPAw/4CphzQNSUkljFSEtMS/zV
8pj12UIruueUfgBTd9JMPOF374cIXQPO4X4/zwyIVeDUswBxdvLtjay2VK7gBTmxp+WDfG6VpWiB
dUQRiD4DQc1phcvdyV42bHhNzPlyZnGheaDNrpvZbAo2CHsqQjWGPbgPPBBdCfRDpKZi2zOnXcO0
Y+IDyWBCEDK52T68Mxm/ZDHybKTdEjTGWhtYlzXQ74IydQuW91H188T4OjiJhuvnNCKiCOlt26Zp
d7K1zOo3PoH0S+Uq4J/xPWJUYbCYz3m6yG41JdosY0LMJmSyI5Oy8QavSny2v2pFbZbHOv3lbbgU
q8nNSxmNWcqP8cLltky8fytKVvarN7YT2fO3+TZn6j1wyGARCxouu65X8S/HNENLHejibC74eFEe
2wu2EFD17AHFd41RoxodSM91vVVJdhxbnaWr9FgRtIdXR2wJtRmFFAcjt3FfhbgBeo/zjx67RrWY
bniaTnuvOkm/A3Xn7a+oKvgqq1z8G7SanT/ZmZeAB7fgLLK2sWxH3mT7YRM/dk/zm23h45wIuDW5
SeDLwFRoM7I14EVBUasjdyhls1QKebhzA7u5aFZwKAvaRMTImbCune9nfa8/SHbk+3jwC6pheF57
SZnc0QzD8g21SgN9rmQfu9icpswvgFkAj04ngTW3qvYTYbb8AUvaJKRugPFeKQTdX7BM3G7GSrAs
O//XFeTEEGxB1ZgzxYYS3dJWfsIf0jM30w4uX/yAqgvajkN9XBHHqEQuvHbKxjmAWMfF7WrvK8fm
Ekw5ebb58O6DjWMkQUXRrhV3TLwVXJw4Jfty0l5i9Eu9ThMtNOfDlHUR/vw3NiAqyPQB79/me+IW
m0w31YatyHX66zOLxb/lB0uk/GUNVF+J7J0EaZgzIjNpUS89ek4AE/H39olD/g2hRLR8uQpwosD7
3BZy53sWCI4u0LCM6H5HO1I8BKhPtOeza6DaezChYatugsiYTYd1C95HKBd89kAqLd4wk0yw62v2
XULvu6NRXIDUdqc+2IR7qAO/H3Ht+zAf+Jd9wmbFi8THllOcfwGWbC1/iKLOCONXmQsDctu8XA6q
i2dUHSpn0fe+c2H7dYO99bzUZsoy6EEeuqpLkCEvS4LvxpDOdu3Nz5LK8+GRwhAs3iWsjjA0STdn
g9zsZv5N0rOi0dqRS1N00wJ5cuWVrcGdqiCpQY1l3+ikBvRADnqm3D1i9tyKtpAC1Q0oL8AYwHTi
WXJ/cranYLjpi48r5ycITocMY19wdUt/6INheCTvyXKv7bEtMHLpM34T9aof3ogvbwvSFXk9+x0B
hMWtMgxSkQJg8LmxqsZtmZFQOn59uBdcKRCD0IkHbADd1yyPK2w/Xeh93QylSoXgU4iSBLLMQfor
dC4dLMxUVjRuzXM1NfhvaRtfQqoaxP6wBzriCxcFMjq8+pmCgEGKnG0zsH2VaNAoXEvjQjAZ+ULX
fC0oj781BK44ROjY+ohW/ldZtFaoquxOcEdBMMmkP4nNy0tOWE+M86WDdtNLuk8NnCj4+Rgyq/7b
ypcjxxDt2E3O1FnjIkkbN7Jx6fNybqnh/WFtwf08tfSsNM67QSfm0UYhaXJcLw8fKbwI08J+0Lfp
GuS9chkK7gaC61FMebTQc1jZyMJ8g8bswZ+IRAUWx8GTIRrqxA7uhO1nDoWY9YwqOihwbL+azLYB
sNfKS1GDuQ/uGKyRVS7r9YoHbNjV88Q6Hi4yY5WAVm4wuoHm2X4qfv25hs1l3kwQzX11/3DcFEy3
KfQoNqmc0JpOSmd39b/sEnbelWtfi5OGwG5K15KWgHPPKC+KmgfoOSwxDGERk/wvh2Ul+WK3+1IF
qrQJDcd8x4laF8IqCeYGb8KWTsD4nBsDKrPSKtN6VetoFAKEt0ikbXEXbDNMAGnQ3JkToqLg3UQN
vsjC6vbzqCceKb5z2LMuzcjIEGzBcvQopXrEra+y0MEy1iYMLd81lysy90Y8MQ4TnTXoWIBWm/wX
OuYuqHtGbZs+mV+5Oqa0nj/JeusoVE8j83BKEDis7gw39513oGEGMBzNbdjz7tebj1D4jMieCDhZ
ICqcvT3PLsaXMyjCa1RAwyM47j6tAou/jjX2jin4+N5Wo6DujYxAmZioIiTy56WPq5JpHczBTjX4
90v3N7vP2zaQj7yskH0Ngh9M3ZayQpO5v4ezGpqdUHwAsTj16SoN6JCU60yd+jbV6DkBxs8vfBFV
1pMi7X7NmDd5fIz7DrUGuuTuXXmBm+YJn5UysusNuQy0ilSe47sB2/2VY9KPACd1xnEmq6Indmpv
nqC295AbHl5CtuHFIG6KdR0Mz2NlhiDF6zqG6CMUPyYNStdq2PczNVSJNX+nw0EdmP4XX1stEm0X
Jz1d9wysSrrxP4z8r2qgpSsoKyZKQ0aI2PlMmgjLEUBBAKBLFSHTyHloiRlg4AI/1shdCOSckD3y
hFsG4T6k/Mbs2Rs8ksBPpXCjp4y+KHgb3zhN7Zkyp4LnDaieqlIYT8lspLRYwDSwx50xWnHpPAhX
4p8ZwZCP6EOyzimuBCdtKyYYMo8PgmhR9rdv4lOjEKSTP10gXdYZS2D/rM2Ffk/eMsQBha8aUzq3
Gy+4VLYAcm9JVI2TgJwOuir/SHDsVTxV63+HAZSXQWGqdgSbRKQQmEb5PU5jxvtfnsILgx2+piQ0
Eo+78pIn0bHP/2W5qK62wO23rpRtPIyHhIYxdC7L9B1bATUHYdD+EiYYrmruDfyq17cc80PBBFG2
cF2Unr1PT+EzENeAjW6rBfKUQvS/9UC5JeZQhmKVeMy0QCxt+pOHXevEe4gx6UraYs2jrALDFykn
WYOgJfVsjWU1c7CHGCH5h+clZvO28PrSoNdoj+PXwKI2MFCbdiFM97ejbqWtotkJuYP//mZWCJaH
mVDjo/QQgUTEIZZGO4yVfe/hxtFpxjnhK8KVXsI2JDpHnB9OWmG4LCNmnKBxkuG3UHgPShOD3y5g
0ujqZrTqVdwj4Vg+yMpjJYXauZIdCC84BYoHxL4bqYCifE4An6AgaKiEZoCiHy7Cj0Syrp5On6pv
sGu9ua1iV8uDBUQ4vc+JfXK6AkGeZ6pHKdOrXp9VEYmlSc8WHSZd95WwTJ3Gc1rFxiSjDU79mg0P
+/0JBUsxQpIRUDIHb8XZjyV9LkO8qraEr6tVSZIQ/Recf6L0Ve2DQEO3BFU56Ned9H+Rt1kqHEvJ
0q7JctEkgoOYp3GqN0U61gqCZqjhA5FvLCD1rsTTl2xsJUI8UFNZ92+VAU2JNiPLs8joYQacwWCm
uuYqpCCdjoqgQAaNdxQFQBJdBX0+Hlw01wvA0Y6zchckpyW2H7H1z3IunSMdFK2ZM6LE4rIAaD5x
2/L/jDgXX39mhXXZoZnNGhj2DDnYkBW0T/stcRnbnqXl0gQN2JgggUBOUgPnnV9yE1DXcoZBJSCP
z57fLZYwd08qli9Rc4voIASDA2YJ0RXf3D5UXAdN6MI+s95cHi17D2Qp5R1iFKR1C8X0LCTfwKGZ
BhDMd6keur0X/bEKAoUND07xKSBhOMPsSSQZ2/dWvcgfkHyccK5y5rWEeBr0dNUSXpHYQVX+pvt8
eqVwtaWT51GUWEMT5vjdzbaUfTqIvgw5FpMvMBsye2OnpgBuk1Fg+Miq5tDt+3s9/LUMI9dktrHG
nInW/E6qSV4OYhaGQ4JUHTmwPX+qUXprCYy1u3gAXTbnTZ5RAe7MvhJAzE0kt8my7PMekopJ9xtF
BrjuvDzizV4pmNUWTK6J5ydhNxREQbtCnqfkwVXgMCMRv8AYJA8aQEBqat3K1Q36RsZxxs3NM+jp
mmOnTtgXmsd+vXfiQh/DX5cpB2xl0eolANjhkXClwOSSt3soqORftasl3d1jwjYVTYEpaEa8tlgz
6UPB7Mz4eIo5X5ETgP+gzkULsvqvxz6VT0cDaGhLQq84j+2jlELuglHwKZYAX3fyoVkfPP+eLKJ1
3cp0s9RAyBvkTZW8F/Kr8uiJ168kCs8SuVo+abyXRviCutIxMza1jCnv1p7F3R2KNBfeKJbSDsZc
bxtYNXhCR001TN2Gj4FBnE86ikS4HzxhLgUL67IEocvETjoqTghYZNa163x8i+Z2FC1H7uUp/vYB
ft9jZha07UvdaUjBnKrU4EcqCJvqvHCY9xYQSLMtV+U90IKRlnTiqBK8bIxOug4M+FNkj0hf9nI1
/b6JruPK+GHO6Ecg+xGXSf6m2NDhQpVcQonvADdEaT/N+2CVeZvhmz+xeAf0SuQn6o5tcYKV2h1z
N8Eu2x6M3nBf5Z5e4zkQPe0KM0uVFBcvPj+Z2F/GYLJnFqAVFm17pPjJUlgTBJnVcjwfcCuZcksQ
ot5AwBtij9zjC/k9A559Fn4hnaPwpSHfj5K2gZeWAxqGPfhCvli7xYUG8SZIDTbSLz5PzG30+I18
AodcfhqZA0tcUScdBiQxUoYCChdswt1WTHqcRNh31lmNVzOGsTNpywyWN5DFcg0RHuYmKJu7YfYv
ygvDwp/EaKeG77+mAetBq5GTBrINM5s7kOTQfshBpjTkt2IQGeAYm/9I6XzhYAbZbvNeetHZ8r3q
LsImYflExKOXYU97hMslWh6r8Mat3kuiZuLRLs16DDe3XSK7vmOGYh5KTCjYFujCVkYP4upJ3IXo
OZQqg3+cx9kjRYvWwnqv3vZxrd9BRec8rHBCav39+6H4C/CWwKsFKQZyGGbDmwW5DC9AcYU7byIw
N/yOz1+VR/MgYD4S90Y7EfPIRr27kloEMT5JHL6eC2jchAJkXOVG96eLZUxtTe8Og45lf635re4b
bBSlOv+ND3bvmgfenl8D9Z1e9Mx7fdVXI6yRfu37R/4mzO2K/DmlaFFDovcI5AWSVGv62G2uAvZS
4altBeFl7PF4sLp4abxKFY+P1loavxdFXV9aEYzPpYTpG6CqVvYfBNOqdGFVKwjk/D5zR4qEcwYK
cX82mHUB0narpcAgz1O7+IG/jfxa/Xu3BRei0YgwbE6awITQMpNnaTZaDs33azdpVJV6iHInGmJ7
VFUb4Hy8BSO6mlXm96rFV/CLpMssUeiEX8Kj/IA3WP0RhbVyPR5FSdO1aGurgcg9c8wJwwFzOQ4B
3/JCGHDy+dxXzzuCdMTQQFhyQ5cE/ZCCn/5/NbVyu62fQXxIbRj5l8BI/penD4Ew0Fe1D4wcmolO
W9R2lTb115smdVlMpfx2WYDTUqDzIf/xpeldbdPxZFu+VosoJcykdb9X4cPZ2eLpx48km7Q/rZR6
EMhOQX9KLQcjk7m0CfrEKq94l5u4khSPW6Io7bPjbiEtdtpV7wgI3fpjszR9SQS+MpPxXXCCv35c
l6HxkLVhEKdmrHlTFvOHomZOzqtrIvBkyDtge327XyboFSne2wAIkiv0QlKSY04Yo8BfUjUEP9kD
FieZYFCpptUwe00rSGGdQ4GmMITWxayj/G4u4hv8l/1oeIZ1Uige3g7Ai9WLyEQRaeteVnNtOqz8
PA7pNojMDRsq7IG05/LZ1au8N0ccaBV6aoO9mujWk3x4qI1TAdZNC73pvfy8pCaDJxFCHkakvhP0
M5k/vK6g3X42ol6lQm2zVP+iKszcVHhTz34L7mnQ46Fk5zEDUSJNoDTj9Xv0MfGkERnFzJfVMCWc
rkgJpmry8Z5vXJ8/vnVx+s9Yo1zvVvr+ayGpZBZt/PASUznaWx9+lxYztaFU2rO2Aw62xfVJhgFp
vMYVspx1G4+53eP4qfgk0jotmhwAa8ks593n4k/cCium6oXj+wPPbVTPUFeNlY+5rZV8m40RNpFQ
enp9n0X1r6pRHnhSWkxus1paxmTSfg+ej2yo8UHEgcYXbWUAwHfn2snXkaJT238nwedeJkUSNCg0
QjrSENZdynitemiF4TQc/6wmnoeRilhelZ+CLRFRA7igz/YhOTUQw45EVDUzbPRk8MatWgCY7NGF
ItQUhTAxzim6jhPI8xHTYhPoHV7Ui1RqSfgpL+eM+Ml1Es4DLX8vHxdF2qVzMjtufAbosrL+HZvX
bcqyCNSVibGJKjgvdw6J8DrnzRSJWnjboKqhBuupJQ0NPvh13nUlOl7eyU0MSgbjkINHei6IrbjG
gU7sEyFft8U3Nerbo/+09LX88Byu4uQZm1omthk0AFWaaHp4+rqef398ItLjy2PvQFStBbOvbwHb
uGns/WGWa7LungGFdulsmjfUsXbKChu4U3X+O+CXrNE7HrxWT9VV97bLo0sOyeiCulpkavC2Ovvx
s4UhhI/nL85/nyTmy7QFJzo/JUOLRcNL4n0IYpZGKe2vauJwErvgdOE8TB9IckFFn0cqh348enhD
U9crn1X+2YYGO6xGYKqJhWuY2OVtbIsEUA+mYuztgn5L33/f+XRSwBdZZb/BOoDWR73/B4Ix0vqf
II+nQ13TyHStEDP6fl8xnHAUHQ86O1xgWMDustg/rzGqlp/zP4iPPXK+yJ0Fr/1aE365PiCL6XKe
Kr95T3PZmubf9xe6EFg6EPw9AwkK0YCs536ULYPzSsuxrdE1lL+DWGhIxDPOJ9Zk7fBSsqjgxghm
Sz1vVsnqp6bGKPyTALcBUlpzVs09M5wnTsk1W2GnqEJVM9sXMxs8RS9xaY9TXMtSa/IQkx5m18Px
ouYdBxnQ44uRMTRdyLTT/K1tpXRC8OQNiL+K2wEbSlVL2vjCdueeL8TYAPlVDjf363J183GZhpHx
gcBjsWeBk+7rg6ft4Tv+JLPBQVIu4C8wP+t8Ri1iAUwPbyX3V5I9mS1dTGKxgb+SRWotURH/6yni
R8WEyBSZpAutsi5olr05mFe77HFYzVFbRD61oyas+SUv5Cod9CFz+g7jpeAoHQtBT4TTRUpEWUha
6A2UGB419lbDQpOy24cNDnie/YCLitKv424VhAs9LNwsKgtk2r0Qi6MNbfrPhEa1ysmu0TKY0dRL
8cPMCzKrkgAb+0yAtnWEjxFpbX2depEUcimUrZLeT0LaVrQR4RAjKPhW9LnsN+Oak+/w08L+B3Ta
z8C+fOVJVtSdH8LfHtlhI/ACqWeAHfxyo2glz15h1ZFimyTRwZip4SoTdsVhF1HlPD41prp9iAsE
k/gg2wXsN4/991sYGGUHBz7K8HwOgzF6/mWohO3dwsFDg6cXiGn3CoH0/EY8cHRdv1eUM9AIxfAM
pHBGOWQK+867AYLXMrR8i12C0uaY5/H0Z2nBFS2GncBIIx7rYYBOhF3/ZApsL8DMNitUwoq5zGYy
ts5hFFJUnjjYk4Ysg3zqP3MHczZBhlYJ33vF9qf960PGkOj4Pw0+KD8RLPyJ8gD7Bh8dmzoyTvMg
0kxgP0bhSWy5HNIXZfh6KERVBBBVDY4M96+Tv0VJDyZqP3SDEPheYcOKwvqT7yZIA2nUDjMAjPUY
NPiovv/6UovLPcNpCSwEaLlNG21c95dhhiJMlgepX4BzbEohdsD7R00aSniwiwlXDMJgk6OLi7ne
nmQjjVMsp4UFpvdIC6ASBn3JhGz40zfKOxUMKVKyzTtjAS+hz5kdRb4OOubNUM26JtlWeASntpFD
oMZtJ9sdMAv8hjnar6S/A1MKTg55zxI2c4ibVeoSO75vCeU4v3mgeasc6DBNkELgAcdNz6m6E+3G
/zRAlAV2sFwXeFGFa3uwh6yR0QtIoPxTUGsBVD25aKu//FhU8r12S25uuSOCAgeSktlBcj8+YDy8
gGMEvCN6U0shZ2Qo2gx8fW+/eIaybZN+wbXvtP+MkGEiNpUHLmE+v97yR3h5gyFZfBUBoF0DDGGj
AzNVFkWbKsZFIwdYBKYzFWKQEV8DPkzZ6WLuZxjtF3nUekIWWXRZ8jgWN3gGsScDUAGD6Ye0bOqe
TOftSN/nUEVop2d+/MieR3eonlzYaNNQ8hrTRR0m/mm9eC0wGMH1HixAhtxFiSdTvt3Zth8yzr9d
X61nrni3FxGf6Ir3LiiqAf1LMCKbRdvhcfHS4ppqLq0L5Mff1mwWIVwdpGji9BMJ2modf5chX6tw
Ki/ChCqnv2LKQGvJ+D1lafSAQqL1J7JwBou0YfcwFXQC3l438hhQSrXbtp2Z4G8wxnVvmtZBywbg
iCgogVS2W7QpJ2FeKTmRJZA1C8HZ5VKfsmsuV2r9liP2hUH4CThpZqsfPY9qc9gl6emVAxOQVhTO
DJtBy70wma7+fFDbnvdMlQBmv27A9gwrnHpjNfKDbyyZSUptd19f09aAdJ8u94VfpH0GKdVTPhwZ
EPcu9/4uT6urwuXGNrgmH5Izcp9/l5u8xFqu7rapxxHagaU82VUw4TphYVz4LGhIfnf7a/Ag1Aur
kHnW2HMPgxcHGc3GnbN32SIMrD8BoaHM6OdviJ71A6BnI8iJYPRVe5UWaaWr1MbbRl1cPrZdOS45
eEGb72ISHavtI7VN/ecUHyLgps5n1QwXiesCXt9uOWgv7i1PqnGH6hoGAGfVLw0OrGBCn3Q7hrVF
YohiekeQSmj2a5C+lGS56GxTiZz/kbuAhuPKPAgMz4z4wyDHznkzwr7RNWEugPZQh01ZQRm5hdKp
lb9ayGbgDYoE93TvVzilwBkv3pOtrmlQogCrcGONyJTN/0EK7djFJz4Rv30brnRlHNYzRWHo3FUT
ZgHhZ9T2FGLb+ucGXUdUPk3MQIT29U9GbVNhvVJvQArXy7W/riqQrVQkyqvR+xACkxeP9M+xMmJu
/1wsZqZ6DxuQLmomqVji+dYofqUmnsNZHa485ko2PgSdRBXxdxmSYOiRwBXzvSz4H8vMomO5vjSt
aGVwPnbMdPnoDgGzd5HBO+6Td7fpcC/dfgGAcrkes1kHlxklxWxHAtdElSxUOFhiJGLY9jquiYke
0idELwzjQE8wDaeAKexNn7zvV8yYyJQIVS6I7Go41Z0nMYRtN1OGlVxR4iF/k3e6+75ryqUrp8Qg
lM/dtYHartdJD9kd3LDo+QBmU9iq/YPNEQpbQmwbIUVO8dOpIPGCgEDBKMDemC6EdMGgnq51wHf4
77ZJr/o+rCUxWLOZrJHv3VTo/LTK8Ip0AGQLwfM7Rfywg3GCgW/mpEmEimQGLALhZtCuHNp0T4jF
+21U9lp8GaxR1hMP+R+XxZzstpfqVTFzuDrgTj5cg7g1ZzO4vY4SwL1E2DLr3P3GIWO/CQjJr8o9
AeCfkJ7dADWexdFVWCo1y1l7JNmLj5OcXe6jhoEGEUH0aTfE7OHe9SX7noRKqlimd6/UUM+nY0vZ
+C2db1+qOyzJ6WL7sxww7ey4K84FwgH39Qajsb5tjucr95TkptxS49mMRuIHih9mg/5yZPNFBuAT
tYIbmyS82d/dtEA77+02vv3gZCICqf7Za5gJGOS+9WuPqkD0ZAIn2+rNvnCIWZ7ylWLwv06KJa1N
8Kjr7j5G3Z1CCf8Jlnf2oPpfN7w3yltaieQ+kdGlbxmKXAFj1IefYrSJEqlWtU4IaeYscDZ7qI88
wjw6LphXoupWebdGk4T8MwdSZ1f9iZREdoNEkLqplGqyDp8Y7f80yqEP0DesfMvpAXFfV9loyPW8
YYEa9OYzNFn5wZdZx9MsLC9AeAPqBjsmhtFd/vNARqje+agcTSIFI07Cn8UPFFDdqNq3YuQKPV+x
GybNJg5sb92OmgsiXNLs6m1TCDM35xRo19ISaxUHIsliUtxkG5obPM6hEvb+YOTXYkZ7ZewCl7Nv
n2/d06RqVpAbulTvmotuV6I3Mt1FZEKsHDgyVinOYHsxftU88lQGyu+CA5yhUzfOnvuid/BSDtZB
NmIOaswrxwyE4C9Dbb5MMWffZSaVjSxUxu/uhqui5IZAYPn5x9I1oc4ss+lFNVW65t7O8Fvszx0y
E6Ku9fc9jstEiil2/owfU5SC5YbyBEmhv1S+gPoa0PMPycHyegghefJaHd1dkB4/9gk+a4N/GAzs
2CiS9eylQx3Y2Blr1C0o3DxTA4AazD/xuDh9pRGGKKvmQUWqhb+8FybmkIf84cPLej8dz7P4zQBB
/hdjlENrm6IQqvTkXFK8QlPvyRniRQJvTglvJ8IWDLZr5u3B3hU5DZv6zi+nHcqN/RixSMFLUEdp
xjGwehOOsXGr4aSjRwICiQqTSjvyZ3U2ZHEpsMesuZL/VcBWFA9M/IFmwjOzJZ6+/pS3nt3O+mTH
eBHyXWchNwIXe7OvV4OxYH7acIRR9a+QwTjO5J65qfgrE28zuSDLeD+iDlx6Dn7iSDcU8HvicDr7
5xZX9wfeh10Tj3LFOFszu/2Dpn0XNb6QkEOguHjLUO5msdQEwxKTYsUoYjBoJ3vNFM8ZWCJwJpy9
Vfy3FvFJKz/tGvvMcCdsMiI3LFc6WC+XDbJQ5GOtLFQWWG4C9gx5bO1PyP/Nk9n9qE+syCboIMvk
KlWBe8eirfQkPLaxLQgkaB2XzpOCH0xNBTi3Ze4vCsR1dLyhgT1WX7Q0Hx339AlVdJZ9jeTMqaE8
NAZ4X8CKCwXsYR8tsAoFxOykE3lbGBPsx4qFwXEdjkIE30Yjc38us0Tz/tTsdtMVYzWLQ6DZLFTC
QvH/hRMKlt9OQgeWMX21pv/p9okql7AXfUbQdQtzUuY1VBe3jge6cTsORtCIZr+otFNySSwGvf0T
L6jvUm1XtLv6jUQxR1EhvMY0hcT9eJofSwGR7Fn67JoIofz2C/TQEPP7DPqvnqGtBXrduLBRTx/E
4TL668y5ggjwARhv2J9D0oIpba0QSTti3zoASN9TxLr0TTy2ey854c5zptpJlTC1/9AAfB1swOf/
9awlUbPWVyZgM5jlww5fZLtlfNkjSTmp6Ch/25MvEluEKwkM+AlD0E74VtbFCuM7szLMUOxYp6Ja
gj52dCZ4qHlXJUBekTF1lpOf9kGnAPCbTrBmpYXJpRhf/jXDKmuTLLlY7oh74r9flEjzQOesfHGD
VTorx4Q2jNGotokgVvdHq4qFaKdk1UGxctOAsTUc5lF7N6VR8/m88TF6qUjuAjg3KFUN/Nr74VsF
CIA+H7yXX5TddeSEZWy2egsL6lei6SOLiyrxQtj4TLNX7xc5yyQ3NMB2EJgp0NyM2KFCYF5ykl+Y
euO6j1liJqN57qt7F3qLChwuDq+Bmc0MlLB5sW2MFSHF1N90tGvBMofUCaIvRczkNVp+qks7eZmJ
7VeUtnIKbpnuvgK6hmC+oO8S1J9/GPl9xcydu9/8SCIxz11pRg/ju0pwTwLPz1HM8N9VssPwBpdQ
cFjemHIjfagTK8lVw8cVyk+h7hsCy2FgFRlGlXEkKf9pkkMv1yyKTGxXT00fyYp57K4NBGtSDRQC
m5m+axS81dDr09h8+KWo5bAUqjvr7PdQBWMP7n7NsZhZHuBuSbFkUrXNupABpcolIx/ttCAQXLRI
uI3vKFWdQPWdcOBvcsnI5mLDMuh8LJ/Nv/pSL56NT+rmQJfI4KPGRGBzawHXdFhBmlFH5FpLMusO
OG66sCj0Kw+zk1bNLPRUhhwDqZ9SZ8eBfvse6htsWXMtvPCiTOEvqrOQzi/6/wkt2HhKiRirAPYH
4VMWzSRccYR/LvMK8F7BxiHSKN/ijWbATyKmPyLtPJPWnfDCtsLtJ0d52zRjlr8PSWMrO+oqWs1d
/RXYqok6D6Wwf7IhxHtpR4Mb9aRw8SSVrHXomNuLPgAvWNYfNkRy7rB+II8UgOS0GAvPAyo0g0hf
Le5FWvCdDfukYm8UyYMwa3sf+xVejNiPBYpsA5FTpMeE1iRfWhM8bktiRdIpQGaiGaJGz1/EcpZ7
AGFnY55z2vMUa1HiC7dYk9uQR10pkEwcx15bqKLF7zTp55H153BSDKGfTfmQZJsU53H6ZpHolYDK
YFdDGOBjLOTAaRuhZzyNiuZ8SzSZ14SN77XqRMUcitMHWBcL5DQDAPjAhIp4KxjEAqfEgjwMOC99
mJJW6l2dcZv5p8en4LHGZ1TK2/owq07BOobKmPjO3krfFs/NchpATYIEgXPfUndaJVCYmDxJqXb5
VVZW3MXcpxUQMnbHTCMRdyx81Y8dHzJAm4bMiy8dEzs2+Kg7y4fGsXGhP2Q5nDSjYiqQ4kbzacve
RPGw/PEBrRVJQKJqSTaw4ytNRwHSfklcm+THp1hq80PxJw/VgvBpsPnX4KKCL0w/pFQ5LYA8EHNM
IJF+rg7LkX6CWjvhbpLZwnvdL5al3cwtj0N98AXuObYq8Pkqoz6C5Sztg6jIT02Zc51JpFPw3iIG
AEQ7hvMJ3tpwkdAp2bYfh+d+NJl1CI/x2y0FU3cKC33u443bnXXKPE1Yw0iGVMKtaNWs4dZ28+L/
ulRXglKXFiYy+ey9KQYgGudUqOwlMDMkacVlfpYLECOmhxvDRZXuy9/PSTwlWP/FhzwTqwx6CMGG
Hzrucr1xo3WiIHVKiwGfeQTueTlzNbNALOIxvCN3Gz4V6Do1i8LI2sxaXj2o+U4qOJ8UUXLWdSNH
qYUIiMiAIwXixRxKiFTv+kAfZ40POsAmpxtWGLdotiUsAjWRhaettsdLKqSdz0rsolfWB9rpckmf
Ile1V/0aF1sxiW2OME3sxPHl6DgiidXeq0I299lL0C9KIqmFGbNZdCp9olD2tE6PxF1j4lMMOpD0
t+HZnFWqDCLa6lMG+BESbfdSLTWN3XXU02UEHO7Eb6g9Yj2p0pCtLyn9v3xQ0PBXwbjSGitRCa/Q
Ha4jLFE4E4IIUtBH4Wsg3sx3nIaXX0FlAsqfvC13QlqX0etm+cBymJiOgXsqIffqRx9amtso8V6C
r4VwCPWkIeKziMgwqQnh8OgwIy8+vwbezpGNsR/ZEuTGZlJKwH5raUQ8P1LGHilTGrbKZO2NZu/y
gKPtr2w1My2r9pYCsOd1AXjsfvQTjyaT0t3KiFEpQHceajtPoNHzM+3sU/iSGdWcwmVm1pS2dEot
OLBAQaQY0fdaWiSy/SEwslo1knehupe5zMYlFZKkzXjaFm8Jor07bIG3bjdF278lbgwUTY414u7D
+8UNRFBgTsbKZBYiBaT5OEXYusvYwzoKzAv32UZSDiCETFysj6cxh3MDtzAGwfd6KcoBz9SwIAMU
dX74vrpmo73QdmbvX+FZozQdZ2NqKJ1eVL9uf8QQxHmYrw3SjMm5zxL+NDC1AIvU5qNOCL8b4UIt
Q5o4y16Xkic9qR3ZNZLCyFYnhTh9pl6R3vkhZhi3VqmpawM/NiXrP9ZjqQJDkt5zqK5fcv+wSL37
uGXdJm/o+Z/tLny3EPWoMBnU2fcNYYJ9lUs24vT3v8oBN3+RwNRKH8nntFc5Iv+ja2h59dECy0Oy
kiYeYUBwc5e7SkXvTpWQ1a+eQuNAilx8X4A2Nt48g0rSDGjByyZ6iMcq6JBvmB62I3SFQ9dHiP3S
+fG95L+f3AMZ1mv2d7vG489COFaaGrQ3xo8UXL4dGMV7/XzvHm+wy5v+bng9kVaNMahGo6kmPiXl
noHM5QCFgQHICNN2PHetuvOV6xXf16fKFwUx/6iVazsCDzKLbEftnJj1ukap++VFKAGbeDQ050zN
pw4tH/QggY1nTjM+sbqAsWKihP/eXwGdozWFm2c9dttDcD4RhW+EJZB0+7OZKK4utGp4Y//R0a1X
dMCtLLQrmjPsDcNF5J8bNA0Tq5P6uIS5uL6Z4rCnJABziAPtRIFm/pwd1y8AtmSqjh6Z3s2aXo/h
eEU09MW6PpNzQrRFWCcUQnwks8baFeMYr8nGZzUcJ44sv0x1RcVh/ZwvrjGO0KcSzihwKqcNsETU
vNg//DJ+vRPzC6pQwNS9vzpQTVUMdyGPhBG+5twB1+f5jqaPD85786K7RTrzejkNWKEC19zs9lpg
2Y3Q9s/l7yRwckXXAa0sAS6//MIWPd2V3Nj8rIoyPwuIOhRr1gIRmfaeUjM+aN57elzIwSLzhztq
aHL4Kf/QTKIHumfzPDzx4WM2U9x5X33l1/rzNDQjys8dazDwOQNW6sjj5C+uBdzQCQQ9vZF7R4D3
VL0FV/iKVGnXSj1F79U46B5U3fo+wXlz0vlvaNQeBUMGaZWyZW543dHhqX1iWZEhxTQme5r3e7yV
sfBkYAPpiC799tL/9nWdX1e78uqGzDSURxVw392KfrHvM1sEX4HSgcpURrt0PiNjZm9AKQtJRYhw
T34IETDGwSifO557RJCodeidaAEvi/n3VWVTpO/sVc66/V5KOoLzDqogutc+/4TpqScb0MySVy0O
n5wsA9xp34ZApkNa4qEI5039eUP1SUNA2x10nIYCLUK+ESKJeeVKJpQG4R8/5U4F0WwMsDOt83u3
1+rE42/aVvu3qJjYTyDVNcUVNZWSOibh7iact/aYdonvDWuHnTh12OXxUgZMYAlIcAqZKKVdT7wA
7xscMKc0XlRoRZshPVE6y2+tBeh7oe97C2NpVBSHo7jT91hBh3LzTeNjxjtf4IkLTrpNJ9LIHyAP
DElfFQylE+i+6k2H9oRPkmS4Evr2Rqqe6widnI4ivmZw0DVz+6O6hlzMRxjV+raaRYZy0la4g/0L
oJ5/kvTK/4XM/duN9wvCLkjUFmqYPCxyIYhZGvxB5yl2+XpnYHRNrUeXdkWdLggguHW/rJL9LYKu
GwzxgEycDqQ0HeBWYarTqTUfIPsVkq++p60xNDI9Ma766d5uZ38Au8sCvj/qHDG4wrhbrgdqSh4K
zE2jKjJx2vaK9zRP3ZZTlVQBi0vraZ8E+Tge5/XIsTZHIiMrSSNdABMfWmjtx7njCW48O24ksTuq
Mg/sAwIukBhNGsJGVLomGeBiYr+9uYxY0rrwciSiwThkKsaDOgTfCha8HEpRRgWH17m7PFoqf3Hl
qvI2NfRW5NZrH/ZptczHsjlsJa/tT35HxDyN1nZsVmlB+bkdmk13IkbSbJxX7bqAQ6xjvS5sXBUS
cpLQoqxe4ISD2D7corICukMF0/6IKZ3/UYAYgMUNYHTL1WH2/sb8acjvqyw1TZd8fFRz8qY8skcb
wAV2MC0QZ1gqZDnMUjk+QlHaVARVhEhEprTxZxyYbmFW3kyprf/4XyJLjwpnx50QfKJanpr09YFG
qGc0HKp5F5jxTRfyEFuz+QQldGvHiyHPsB5bVM4bPrfLiji2tUJn1PHzLJYdgXpjXCWHgmkhlJxW
8IlGB+se59aiGJIjuAxpvleiFdh6DsLUysYtQz9qjWM9TfvZYSB/tptrad2HRJoYRBoKgoQyqWum
Gt5qdRki+uIZ7z4Z1Y3G3BAqZf/8JB3Go2wbz2g8L3GMMfy6aVeekDIGMI9lmt/xXoDRtEnfx2q4
rEB8VR7FrJ96hcb0+Wt4OJH/2BU0du3gVt0FuqeFVaq40tqe2ix9O3WQJnWfrKpv5s19bHdkztdv
xWaYZn4teOcQ7y67Ti879lIWQxdXsHJWqlqGmbCbXsC5kKb1YcmA+QIyPWxOpFcnQloa2sLpahGX
NbXidAFvXQc75tSYCxp8f1P/GQkJ4Nx17YBzzRkgqpLfeBPz6prbij3EV6piyK6Nr/Fx0hDL8B+K
RYd+CgqAi4wWQ2lzDBKc6WdjcOPn4S+aUx4HMFcsP1fI9Ia1kzSRbyJypf/3L03Hl0dn5jHynQ73
C5/79AhhhDxpnTvNRBEz51ccOajGrFazzuqoMshPGRgZVZtOykvCENLUeRw7dDNGEjH3NAOq32bj
IuoAR0GCX3VHxAafgweBMAoRwZi9UDTi7jovEdQAluZoOHkLQAP+x4uSuyaZ3g7MIthgp2sEN3YM
DYxcKS7oezlXRKhBra7g5inOyunxPcvTBYehbdCX7bV0iXLgG3WYTWcm4kMO/vUsOf9ixTjzY7P3
sj/9EFN5+j4hMv7ebDgpbE+CKyf0KFZMhcnTZOaGh7gJ6PlWyv4PmVpSXRQuMOaFtlMXTaLkA2Hm
/dqEEzfi+Klh8Bww3UPDJw9jWvCiNCnzUk4aoScST2EXeU9PeQ/mUa8Tv6Lwb4HFTpftft74sZiy
NnKoDWSvaFczgaKGPsjWERRfRCODA9zTW8l8p3+ZN4M4xxtNJ3x3nIuFojhjq3YXOptaRBH6jWWS
pwZyz8Ylukb0Lb9ogpi385yAJxncgmvvJpl7OUPxCXM3iHaK3/cL13eVowqGV7jNx0Mi71e5m69P
Ewmg54auSp3qxxgpGjlqCcpUO3ou9K2jgMNmqhwfA8KjYfNipwIsfozyn6kGIDggZFnY52H7kpR8
0BrQ66Q34uwcf70/XcmHi/ozk74+rG6DDbLZ6hbYIck2zeSoMjCbtfQTyrPql/vW4uxgno6mdK7y
Rsn0myBZd31hxHf4ZIy6GCPj4TpMNdSPCh1hokxHuPbY7UDFf5xGDQSLcm/1DZrexcyMHnFxbEnF
Qq+0keZIMDPlW2O5ssGrQ/xZ3M+pAHnZe1j5mPl72HM/82Yi/cV5pnlozzSVSTdU1Nx7B7nz684q
wKGtw4ouv5NF4BV6yJbecp99cHa5w2qtPQ29FHNYGReRcL0cpl8cX1uBtIRQjI/58SyAIn/GXjLr
2URCNqiH6NzxmHAPSC+sw2Vohy0fM/AnNW2W9buDPYXq5oGn9p42iVmnzn7gYEuh0UgymhwUtx6s
HbdwhWmtdy8IfwDyTNVNWrfJ3YCPAg/ghIOCcM8lj2GeaFRvBXZMwF65phUA7mAKEo4HV+pqvtfQ
wY6ey9XNka588QK8FqFU6nKezkq8Uwa+NbMcsqBqBltVNtIPya2YnoBr/7tSRcSt3NdakEiZJ4+6
f4kVAytMBMQjXP3G6vPxHi5bU6lGyn0cJ7VBEZGshS2CmhBd8CIM/jUn/5NB5DSrPpyoLXNjIw5H
K59nI7WfOh/TAUoaWU0SNTwMrbEaUktdoXhm5MUqBZ2/+sIJBP3OOAcdHwUsVlHVaa03vNV4bv+M
l1hMP9xqG0FawFYO43ePPmGiUx+RtCX69njpJhtNt0nG/u0do8fFaS2j9YMtcPU/yw9u3y4qD1hU
b+V7XjwdQz8xs9fTB0Hc0T7NW7Acp2W15nDT/KSDh/ZNQeky8oMHzhy0i9zObHg89wl+LLSqPhXg
Yc/9dXhb0HIrPttU/tMAfCMD3nPPM2k/n+cDyItTRJ2LqMozUvmqEpl27gJWAU90xunEjssj5XFa
y4ORmo3M4RH9tXTSSiTME8rshCaAkqECJOZMRLACwDFx2N4T5KvuZ+iGENKkhFu8n5yqw7CkNJc7
TkP50MX3KO8Wbst34eXeOO+aYGuJZXFFokI06udBdcjUMWuPX5rvJXIP9b4JakW3r34KUn+50nqp
5iv/Mncn/0aK0HQs/0cAb3BU6bHrrvsAiSKcikfVhkb2Ym6MQ6YOF4nzyDf9MCXJttr67wm1q/PD
4wfBY8UwiX/2vobUZkaZ6xlXjXHMUeINeF6q/QZ/CkYuemZrxY2Ht28rSl9YKjJrEmG8QW2xYO8J
D5BMYBE7yqtQbfNCMmgOK99JrYik8KLuVNlvz42W7DP/QhncOgl+bncfdlLz2dLdG/yZY9IFnywu
Hl7bsEHNxhcHQcAeRtF0sKh8igPjomJpslOTvKvo+3CwbP9lT68BDsHvqZgNfpmiiJUJpentvdNO
ufy/OOmhSEbnGuxC2G06rRXwoGZoP6RKU6mLennZ/v4XEfUQfPFa6LWMMdd1Ql8xHn6DGl9JW2WA
TjHQKPnmSKxAEP9LveDdey4ShjYQPcwih41lbpsvnH9+AdsUuAdRcb7LBudr5d19/PJGucHsnpvG
Av0T+0vOXhta3dfVdFNXEPJcwkeX513Lvw7faLSvz7+lqVd7gunYgYEY6XGlmsWl/6egY4JERvK5
EcHPFlwxa4myGj2a154kRvbjyxs+7DIyD/Sgxtuq3vfHpw2Q4L+LE7B5mGpzHI3Y9kxsYFvbL7uz
Nj0t4wS4rJNALjjI9njrHWCQrWbAPGo0I/CnlujX3oYmY/X3mQl0ftXf7VaOE8W20IpeiggXV7SX
9y0GGbAKbuUnWMmizO5l2PMm48gM9N/SsfHPCaxXbY4nDTkyw+qDxKhHAqJah9k3zos3dEr2/Jkb
YM50SMlPWuZXsI6OTu3R1J748DKwHC9MsD/eXgzsF7uu405A9SlPQMJKcDyjOYVLwEPXgA7+1ZQe
yz819Xlc5Opmo5CMAsqQ7fBrMSazuv2ZWuNG0Ra/9cUuMn7B5kIN5+/w0T4eUqWiPViXTbtsCMxG
JSzgX5s5UFDfADglRlpPgXYRG/p0ykggrGKbP342f0ItKy7j1WLFRSDGi3t5fY2bRnnFBCbHnDRv
RD1Vn9o8bmaVec+BGQviaL5qcRjGQE6V3Zou5e7yec7FCvA8wHBcQwcMkFBv9/etovt3l1LyKRM8
KUtpfQRIe1dQkaEOIS6opvMJnYXLTe4cDz5Kpauu8j9BMokbAVHGxXIA67aCGQGjvrY+qydw41tQ
p3SbmsUBdyUCHccu91QNcnf3yA5TZg7jBEtNH3LWoHG26xH2YSZMUoWzONuHDBYqajsiMw98rJu+
NtC+m6KKXLjRU5XF3Rxos6w5gfVYQzI6NG10TLjNuDIOar62uYfw/4jKimMdxNozJez2s7u8qCti
8/raq8p33Jg1HO4vspARROurN/5a2BXwYPYqtCZd2OL/m3KKQDliiBlYkMbSZEZXC/M2P/hdXKbs
58peohODqTPF4cy3tP2sv8jUBF2+u7QZuw0lqcZpQT4WGKdX9xOJFPJ2i3La1pebaLl5NdKcyk+i
OBPSvK+FtLc2tGNmy0FKDeSkiRPG23IAMvE8Ly/q5G363QLhIOD7jTj4aqeQCNzxdFZgBJcyQXfh
cMWpjaGW/ag5OALarLIIV/VFgpOcrA6NfcyfUNSDXbxXIGALVBHRz07n9d3uVErQ+TkS+0vOTuwG
2FcZrTASNqfARpl1jVzkRx392wMvb55jKVnBfT7TVTrnhuY7/6/KoMu5VncVrI30dyIQ6L8vKACT
amsMPBMVPv5rThgZ91gZ1UUxuOBatlbAQ1yEf228Qonv8wVm6kVnMjA1y83ZCliaoVILkhR0+i/1
BN5CaSxG5fky8RJedjjwq1XSpYGZU2D0/LvD0UKornz88WWCJWvTRD018dUm9rerDBj5AnCM7PSL
5cZGu/0e34BvLggPSdgMXV5gfWRC2d/Z/u+dwSoxk7TsLQ7uaTDO0ZNmPabd57S5tb4jM2Wp83cr
b3mmwoI9PeGg4ib9/7KFjB2rVnZx3VqzcK7sbtPGZQtCyoVZ808Z5vIMX6MSbvspge/oRb0nCVaj
q6Z06tdSUi/aNzWjRTQcDq12mc1xiIidb7pWMeTjXPMBfl6GIx8wS1CbDSiEsx38f4M5DjdhdG8V
R8QIeXmWsS8iFHXFS6UByBaPh/Mcv72/VwyywOkY8ZLOgdkhN/TUd5ts+sI6ZEptTq95kYrKXvj5
hvqCJQHKz4B9YfhRhvZYQsKy3cJVHIvi0fyP3jmiNhh9r1eFFs0jW3Rh7H4B7j2rRlBbiHZEC5JA
Ze7xQtI5946RAZhPU9nB9YA+o/j5jDDASRu46ibryAzaUjwGEf1E4ia8tL1gor3UqY3OiJHxw5Aq
3e13ufbQCKvVcIYt8k+nJns4Bw4hGskJZTR2gMPBuVTRmxHZ2K16+UZINRCNthaXAagvwP56rDgx
XK54shlay2xM2uxyLnFwVZ5EHZ8jfKAvZwDCFAdv5IlrSwlXFNK1RAnz+TTTYWr0o2ZazJ7kjDzi
BJ7mYl3QPNpj5zHbBD29qEpGSl2QXg6VlhYfpHRLbDTdThOiDYFi5WUFR2fdw46zoVLOEf3cDCKH
GsBOxHgWr+RqgtD5StZ5py/5ZNCSAz0I4WKdLlCWuMCviT6eDEKpOzZowtQ7DXoHpKk85QFHEW2a
Xjy9INxP2AhzfY0ai9ZXDbbIA684Ic6dH6OmWbCsF1bkFQv/SJ38iQElP13N3ZZFiLX15TTND3y4
yu6djgeEfN3Trn8KfsRqx3JUB/Cab2nE6U4oHCskg+n38p4O1cAu9GZ3u0wDhqcLQ2SRoOU6U9OP
SvgeAmU9fFGeD9B8d2t9wzL+nmEhnqgqpgecMonAOWyy5uvlGx5PC6pSqtftyNCOqZi52jGKOkE2
0mo2bJSQmy+as0n+2KauDb/uofnSRwCuIjkHZfGcLHFop0eBpbawHxCI87gb/52qkdsj1NdQGe4T
8nc3bN+MqZjdn9k65vqdDaNOHsyphw7gQuSlwEkozCSgUQsxvV3jzPpEB15KOfNrEgucjpmc5xlr
pWKB3CcGOGPk5L6z+41ziDxaaacq93URnR0oeJOCAOE/UDMjXPFJucQ/oujO8QyfA3WgrAbCbHIz
HJLz1WXR8k/Of5n9S11pbenxFLzSJoPzoAivb/g1fDo6UqRnS1m/Z69jqq6RBcQZPF6C9wECr+5R
PRxyn1pZNWMzxVqKOceKfF8L442SLlJjzvk6FP86XmQ+0AaU6HHaHiOJ+NrhA5JI8W5AlYGAAwkr
xrPTiFbxUB7JzTFcC9KiUDNv7P8ndHN9K/gLa0RxQ71L/ktKPXhcbaLRHjnM8/a2a5eGCVcaM9+h
BfQo0zNltvWuvScsAxxmV2E/eq9JwBbN7oyenWzKJp67Jaf/CLuu1yUoi1u/Wlfan5IqZugfnedC
q6R9vqvXDo/gFvwNwHx7T/kMxkzJzFb7/1TVekTEHrkF4v9OSresNt3P5qr/4pH+soz9XnGUhoE7
K6Ucmj6v/Y3DwRMH0SBlg6qOI7qDpqOWN+va4xeAqZsPJZtRK3t/EE9T4QIxjyB6/IDz9MJGmSh9
SPpBa1+PxoHHYbRnslZidP7jDJCDbxqlp8q3OPoWzAFeuc0OzVzU8WeFgLPMpBbfywlhfX2B6hug
OmHcMLY/Desukk6DwMvSTeEMUlpl5BEzZzKhMuQ4KDK/HscxVge0lIu8K6fVkLbI6wuV5EjmGgVF
jnXDgeYfZ9fnB2fu2APZ1LQO5Z4ivkE0gfU9vsTfR9dnUWdRAuXF6wmBv4e/uNea2oBVZm5s2fyd
Fhs7Ici6g7WzoSqHOzU4aufCQFaXuG+sLuNVMONnMGHKwKQzXPyg7MecB89Ll19M58zY4XqvxhCd
GCLdszJztgBbTA4JTc6MhEkf3UaC/jLMjXQJpZMFmm33BvJbpKQpDGza7rZJxuPS67nWaAyXrTyp
jQ4SB1HIVYS/EZCh1Ez1CKkLls79MHXVUe7fskb0GyKmL/X3GdrE9B6gCM+rZXZBnk5VLiI+sH5U
neQp7CS0rLudYALKV1CC2uaNc2bsXm5Id6N4vGF6oAV62L4fFp+TkQnVPtKquRYiye9Dk3KKPrWa
nm3oI5jORYB9zs2aXdue2CNoHqBaqWWTEFzLtbOzuPFZM4RJEqpZTNiJii1oHhsIZCJp3GdoOVzx
WUQFSVHyyLaNoo97Mh0RMnI0+BmSQm2Betko/acYxYs1EDVFuzFHpgCasFppPVHIIDUCHFtZuATv
WNJnGkz/4ce6dr2d6jXc6Vy8O/DZMPw4UCtmFuVlrxYQJFDZQgDTJ7z22DSXIHO0FDDA2HtvVSaz
HPEBXkFbABoNEUxVT9sKkdzEQ6OpcdqdnT8dJH9rEJk2xyLqDvb9+RwLCA0WTIig/3lTiIlycDNH
tp6cFcNGFtFDwiMLdyp8azqwoCP7XIT1SPeawcON2h0Q9pJ+ikDG8miySW/rEh6HAG59eAoHOWx1
LeAqU1SVMrlJHWy5tp8RkTBXPF3RF4vetcoFOl/sSNw34QrFcp/9iJhBE49WLDYTAjvB6aNCma3E
Humvy04LERxpZxjy3ZPqSCpKNPxgFNBTbm/lo9FrKJZF/0r6pZwAAc6emJP1h07l0Hbq3dR3uitV
WDVqbn9QJunvPnVixgfg3+NqtwgxsAXuhXg8JpYNpglVxero14dzpzpJRmXssrM96K/KPeH7XrRi
hmeTybvISI0+dcvCyse6GYRgOczi4GAoZ14IQsIg8bg0FjubS5LXPk8/VszSBt8vi+cY7TUB8qMG
WxQKumtlNkba+5B+e6GZGk7sZb8Yaqvf2CatA8IYgLDVz+vbAifnNSPiTby2molU5kwSNgUAnrjK
7AvvyU59Uu1j3IbFYZRjK4XUMUb+9HiNz4r6jktElSUFSulAduGfvzjDufGATxZAbAGJUn7aOBAV
0IleJpkae570erC8gF+VzpT1xV2yJ3l274SYumb7ksL7QqLcpvYY2rMluMywAtQ/q8lIh0dHF/t9
bTvObSv2Ilg+onN9btYonXzfkZJxWHhj+dqHv4zEp0fo+gEh0VFE4UemOMW0tgtHFEATEj5JsaEj
iJTHX3s6Z/rJD/dDrMg8JwBjZzFRVwJjpjvWv5LoFokVY1tEtlVTac+sCjESR5KpC5cIt/oex6f0
DgqbPUwl/nLbdkpgofqFFOwXJh02viFxBesBnj8mypV/0MwR4pjhd4owgbINSUHWHbCxPwq0ZTkI
ijDMzxQVuirv7RTyfsKAENRw97L+Sq2t5YlVsiMEtsmbgedYzuFWCiKBYN2jQhDJmGVi9Ob5xZKK
4fWaKGe6q5zqx+9sWCVY7Mhui4p+Fu+ummfGFcPW9jnY560IUs7ONQkQ8JxLlLky5AEQCbEZ2FBS
V+T+6tN5XI4h7QAuCZoVUUiXToUCm1oxX7IZVVQrNdKzNjVuJrFmdM9/FixsT2zZsqM8QbZxZcmd
7JV7nhVJ8D2i24pElWPidwQMmSAIHKWLb4OEXjFlIxeoaGbc86NtGIR2bmG1627wfQXrUYpCCllE
vI6jJ0hq08Ay4NZMQnDU2UbTgfeRAcbf6qrtsxTwIMcsgL4zuQlhz+SqPsXA60MgIeo4C25ScmEA
4xgouaIq+qjkipDINSrttQic7j+IhXP2ET0vIL1I+B7w2k/xyKL+MjJlXXLSzVW4ovMpxdccv0ke
bEqUFTi54gbyH8cNNhYWVXKXIptmmr5ulpROO070E29HOgYurSnlyR8Vhpq44OO0vrfvpHKe/AMp
jIFV6oon31MtPNaFWWQ5Kw5gZTMh/KM2m3g+4X5mipe5muI20ZjUYtO65jOA4+w08XF91L32U2iH
TTlGoogWQ+KXMkdCkNWq5T7y/juOztDmTiJF7MYkM+6iGVxvpUbWYJRLHmXC13FDb9dOogFo933C
GSlpo9r38WOaC+Rb4cuiR+OIArx5P9BVhOEJIjIGsV2ah8yOUE/EobarK6B1c9F1F6eFOrjewXhu
lORdk+oTN9fyUjWFBd1x7NB/PCnox6ab8g07tAY3QOVprJkC08nILTeqstrSN1pYRBi3i10MSOrl
HaMmlTtLucNuDwCDG21SrynjVBuE7Lvo42LDQvfmXMfnsvpXlby14lhQaFezmUKFTG7mJ57Zn4Nw
uHpuIdcHDMlY5WOFRvX9LkPOhPaxbjeEbyjEjGYHLHy+eOABcRvmDFU4JJrA1OrojWza8cjtdpj1
iadTdlyEiEfs0jLQqrRPBt/9m0u/rRVzMVVfcHg4JZ8qrgI87fVPgRAiWpwRKBKWXiOlsBp/nKCq
AEbu3leY2TTdZSKctZFH/n5xvujbGuZXmTvPrxopBGfnLPR+SxNwC5XVEc4DW3b4Z/2R4zYT64lH
xBAwAKyCi46vRB1NAbdoFqDJyEOCINlQyb+Wc1xYBGPfEgx2xqO8vk8kkSFdkAsA+wPEttV05uoc
0D6vKBU1Q7t+X+VETlglKs1Iap+obEkp8LQV4C9tsmwwQrD58EQief5mksjqeu76oSx/6CztW0Qe
e16d9nT/43W/Q9zY0xSKJ5MggFaTm9y0VGnSQ71/6hDdpidInzq3pypNgWKuf/3S8EpRiidjGGlu
KHbhssJOLyPvKPOfVCUqTKqt5M0glgi12pxOolG9QBjBvdDVsA7I+k41jiKLVlxB2KJ6oUa7FD02
HlPsU1x2+RZegmgmqIEQsGH08ioUx4E8UWoImkPheWxwNnDvUNUJ0H/oK7gKbl+UVdvjpaUiVg0v
FjdrjwpjNtMxnryTfkO6CQU6j4ncS/+YW3P8Bd4DIaSVfEUH5xCKMOywfW+xMbQ+J8tyO8Msvqjl
yhc9R9GKRPLPUDusNUAdcVBIb3M5FzIXxUmDZ83E/OqUsrklV7mix5nF53fLKIIFtOIxD4DSypBZ
FnocufMl27WdmWJiWFFHh94+EUJ968FNZ+sCrSh5txgm/rPmUWuSw8leJ5SNxQqeAMG4NdJV+80e
0MZXtYgZusw++2hTKyFsqlEzjCO3ekzYGaQz84MjFI7ibAyMRMgHFl191leGnjMvK3byxPtSF/gg
ua6TwpSwci/5opAss+wbFZQctNM86MONrFTvb37mGUVlXpSpPC5PYeHdIoQhPU5i2pIyqnvOvIKa
EIMHhmdrkOOfQS1N6Z2USjF5CuPQmHJ6vazbI4CvGi359q9ZG3mIEj7YrMqosvP3MAt7IJ1Xt2Kx
DbuV6NUcEIdq7IxLIanqSz+lQP5Jx65eCns8R7KMlDFia3wOrr2RQpryf88A+XfcnGxALhpzKiS7
bGtpFF7sPLiurW4ag7e6hW/pshlqeM0F4Goo/VSsy0M53aU7d9BD4R36gl9et0L2u4wA7UoC9wdw
DFzD9/dVOIMFcbsS8ok+5zjLei6/HBoUAn4rNHEsiAu6ST8PCNkGp3slEttXXmtSqvhlS9y+OZpD
SSxFPNjgW1TCJlmSxCFSSVR+7K9Ncx/L/fcAvY+Cpm2o4xcc5BH2bnLPl6QoMDauVfM+WOBpM9QA
jRAgY5OMNSwtmnAmyHqT7wD5+oUyCSNVGyvBavBg6feaihVaAEaNtlxTjorblNMkbFowtbEWKpCz
4EF/gyVQURsB0W9lTDkKKyGuglk9vFY8LhDpyaWph4tKV9KWhFJbNG0T6YKK4IacjN6uceUE0uo7
QCUsSoxhEUqOCZ8cmAmZ3bTksl6kLGCCY59HMOX5xeOJ6XycFgU7Cga7o514NH+YUuKwceZCCyCo
2tFy5tPrsAZPFimjQFnNNPlYBFFA/Y1ZuifeTtlK8R3pkDvnUMpX0zK+ppxbd0d18EE+0p8kdb6L
4H9Eg4o7QtW2YQf2AWNjFPfxmXjeQGF1UHNNHZaZqsCDG29E9kTXVy1K2knWyGu1TS89mga9cAgV
2m615QUo+6GfZeRkah8RpsE5/5glVFFAuk8kigR8seN2QOltE4/LXdmp9kUtbCgXBDf89x5jNBK7
wuhLYdp3Tx6JTb2Jx9Q+HF4SsR4Z8ENbxwHi9qS2wrG83fHCWIMdbAzJJYfvHteJAKhDpqgqed5c
vl24TGwa4Wth6CIaczNhNtyAEkblk7PtZgd3DDG8tsRuMIiflWMWkS+XYGrLTAT0u/hYz4tU7fiJ
+ieXjYJOEunW3unOcPVM1z/o1QaEKxjE//NXMxIOg38GPtZhb8l/uCII2wSbFrYY0ogdJRKfG68e
ff3PUXgoTIrbcRsHlu8oi94WF0CENA9CjGWArlbAOSGdVZ9AlNNHCPKXyLgXlRvOVjTGBLp+6P9D
Pb9GV+KHFe4YpxqYooew7S3QdTSyMTErM70B9UJR973FPTJ5URtzPlUlp7yP08HabpwKjGJYY6jQ
u+0hazX0Vt3/BTWMB92c4LOcW7dQqz/LvmxmJU4OTs/C3SMZPS8fzsor3kAEaKTSF3Pq1QhID37W
wYu7TO0DUd3VDRM1Gfu0O//bl8CIqJvnVyEQ3EIpm+Sa4LXKscn5IFohLCCk90lZD46iwe/pBN/c
YB6D8j9C1K6sbXxwgnq4IdV+r5otmWOPfdYQaV15Nmf46NPx/PtFbVYf33hon/NDPhArw01SWR6b
aaaUO5ZHl07LA36Kn0K2mze9u8QbAiFREEeCYWgMqxTFkWMchYuqJeYm8rGa8pDEpAspD5Cqtwmh
+8UF8dBHnJaSc9LrcaqK2AiAlgSlAuG/mj4elCsYPzNEQ320Txh+Ucl35DruHw6KGTMV0OPnX04t
Bb1XReCOJMJ9SGV6neGHbMc2z5dkS8gJbQoifL/xYZzd/pbE8BFz4bivn6LGsgifaXCJldDRC/cA
BU56Qg0cyvwE9qEH3fMpfZ2/Z1vTyLNEtBKnwoW6Ll29ckikwPQHg7+ik31xfKcR/fcxUTotVZhl
mSlXonqXapiAbl46kZLrEAzzeD+vNCvN7lOPzV5F7ULP8QHdRgtXuYbxDwaA7K4bUOT7J4i0jyAM
8b3drq+E76ko7gwtpdpItN04meMgVru+QztYFgaG3oZiqJmTm1L62DxYPJ50ewFPsb5c5jEVgVf7
zQkf95AlUpzZr/+trmto+lrWnnxHduuKR+BsX1EcURaB0cKVBD2DumxBs6Pw5CXssI7WdY7BuLsh
aGB2Vf1k917powvrKNrhjl8fOkft2O9MRlXArMJcMBlOZzXQtM7FQm7m95ddC/WLMowc6oyA9MJ+
kWSEbm7+Mu+X2HItb6/Wfk7YxMXhRVr7o5gEFjdY2tdtOn070ZVnVksDM2kPHBK44zZZbxKMoPjI
fsc7gA6/IJHWfixGt7R3s70S4GBtyZvb0TGAIroaE9llaTOuCwGlqOV3FR7SrdeFEqsUl7SsAATd
dhdYQBhnizUHunVGXcr4aJRFLVURCKPB2F4AwkioQ5kfdacvUm+fXYlk6Dv5iy+onTxxj5hxNUCD
KKis0gZOLQ1NAeL1PrfN3Rg1Y6/71mbNQEtjyJ8ngegzkXMe0kuwcjpIjmf64dFtTl0GhzkwH8NH
eFRHn3wh/T7TPB0rMRyGCsSknZXg4ocP7VBDTYOptJHp1gR00mon3RARK3EMdmA8r2Z0hCLK7AG5
YHTywe5JLqJa0JjGPKlc2Uun4mKVYynlzmGdVJl1Na9riNX9wfT3Y24V5/Tk+otkEbUhkwI+fGVM
bAa5oQCLoBMLrd4jsuqFLn4/+B3+mUdJTH2Qj0ImzrVSmmlbynMFDBMPYw4w48cFpxi9qnKA7MUt
8vp/0svUHr7BXVmU+U1n2OZSJcTWhtpbObEw5ioUApeVPV+WYk5nGjBkLZ5SmVfXCRzbJFvgmbox
wa7sZUVBEkEQwRLWyQSnF95O6veAb7KyE1aF+HSC/07zUs7UPcphO9wN0JPEW/FB+oY/gRzSRrq4
f7uyE/eJKUdq3OuFM0Znxyl4lgkDa5MdY71bqXESgpiZ+MggKmMryzB88uwEChi4YPad0cXWbt6H
GUJk/LlDoZb7fgI6I+qYxUEDbLAXrljDhMRSi7nOWcGW0uc4OI+o27B9j0uD6qQ0d2hUp4unmY/k
XhG/uvHDpNH1SLuN/3pgFxsbLLIrozwqWQ6+120HHS6PbXJtzEyqaHKun8s1ha7XjtxQLZmeabm/
cC7sJ3wPrURMz+jM3beznsjlm2HIxzYoDXpw2Xlt0Vyk7dKDJG5xRoyoe6H2OFC/ww1Xvx/7zdQh
d8PIi0An0Rr9DvAXRhCfDITvpqSY7MKZhWSkD8bF36uPD1sIsFEqt7Ds8RTT7TtLgsebg/fFH9dS
kZ8kQbAFVYn+GiEb9JH9l53L/RXwBpAQEq9YYneF61o7dF3JA/DPOI4xeljT3MrdxklE9NorLo1g
AN3F7kQWRtQHIdei4yetKAzP73jnQf62CQ/SpOPpzOo/M9qnBdoLiF57hDjBjxXJBqKlI5VOkGhU
p3By8UlxS5yvPsut+0CSDPaC1gYKa+VVrusQWbMElP2jALrX48fADhOEnwBNpU/O/bTTw20eISi4
Sah4M09qth2JGdzM9IA4n//HANOcS7MIvOg2vEQYtAxIqwXQRroaEhQldoUsL+rYHWTwr6q0QSZN
nbwo8aBpDceftyeYylXYkp3mQIBcWk8JOM5T9mc8648d9YiMQlkr3chCs7g8r9cPUXYZjpe0HGXv
SJ1SdGbuTzcjG4x2A2V1hFaNhwS1KrPt6Gi9GfvZTwK4ZdqQNbKFwAH7DGwzo/M7f39V6aBH5e2u
RALg+KxNyK9YyyNg7QAmY6c7BAVV2MnAvna4A+TOZpk1TXJMgHAPbcawdnwWeER3L610qakBIVLm
OpyT7W+ncUXffdRQV9nANsM2ThwHgNb3XV4KM1hLDp6N39khqijvtutcyY+Be/0wYzRVq6sehcKj
Q5CuHyiT9Uzss/JShAOMwvY/V6VQNlouW1SqXRQkxohG78t//YHbpC7GLzI2CDbqd891z/+tnG6u
RFzMKKzg/DnuT1Ir9G3/8lUDFdIJU7c9vA+fBpQRwaKAMvWairGZ3pLgeJw3dO55fmJBdNh/juq3
XXSnDCRwhXZFdVNH224qYtH/LuaeWgCHqDrm9bRhZgcmo0+N66UPRxjmqm3x/C+r7/efR1STfKpj
aPLUwj8lvsrOYHbqrIoctH5s6z5CumJlluveOvAbUHlK6Lt6QMP2BvBucIVfkGGLl22KFwvsn2AT
NuJM3VvWTxrA68QV23SXUuW5aO98XUoogMpVGR/F3hrEC4dacYXkZmh2y8SBIQddE96CvCH0w6kM
q8UeHZDCD3H+LvB01sAI72E4k4lvbdFxbd/c0ehmzcw5ATi08G1611k4jxB+t2u2vx++PURhBSue
FUao6Z5vYwd9Rv9grV5WzZ3X/eh9W0eS2n+0zraLTqcX6e+dREaO0S2c8t1pE6ccv5TjqAcpdoDr
xAi9l5j8c9EbkxOxWKkIe6cc268+dLtoI1KONqH2vgX7wL0G2002m6uFTdERdbX6tgq3U/EVecmO
NW5awNYyqipWu6pJvMSZgautDW4ajAksIfAVpK7M6CJ92EMTtd5EPLDDL/tTnkqFokzF5yogvg+A
jxsdPDT+y90o1isao7PJ0frDWi50Kj6iXwOiBRukeCsXn+00bRvB1jWkA/ktVhApqsAAy7IlE4F5
KgScdvBBflF1zsFgMRd5r1UGajGYOngJ2YBQNT99tw37KnOTvEE56BoPo4mVF/YOazL2RAdo6Evp
JFhRyR2a9Qysn+WoAzNv9pwVtzYCKP/rvOWQGLA5QZOZA3U7yf814/EG8ba25lnErGe1ke6FYSm6
Kae0nbBaFc+QtIztstIhhqfi9+J8Sp4R3o3s9D2rm8VLZr/Qm3mrdIa1phk+Z/ek/7Y/DcFuNj0l
wQTlU3bsxb3GtAg+ie0wyKzuhTyQvGZTI8XrT9ABenSKP6jWdGwy4cc5NDuf5gK3AAk2WGn6ejI1
zKPcxQ2V7sb3vqdf9Jg2gdulzEpR5G6cTuEdYoTdxK6+WQ2ihDp9uDJa5y0Fx+VUXhSmZAvUA+MT
+5VR18UQBbyeg2KsnTCJtJukDJQwXviCDz1WZQ/GNRGJBnkW0wLPvYtogXsNEg6Rfi6F1wXpUA3A
QfNF9XthDfb2OOTAgNeZZ7xOfX+bx68u6pUaftzCZiqXMjjoikPZFVhrSrD4MhGXUcnGiTUg1NHa
NdG+mWYZ0l3uqUt5V5Yp26XVRPlu98KW3se7MNGGYlgeCM8bhfIjhgOTVcoH5yIWe9aC4Y46bX9d
usBb/9gcrRF1wJa/hqkMG3QmRDT88BkdmXmxIHIni56k2tqJ5k1v1eNxVMQa7z4R2uizKcmIEOKT
AIZEvCNEZM5qXzQ6m8TSzISBtqBsW28SMK7BfZEcT01SwgbsURPpUcEqC15/Yy/XLP2Igcvm4f5J
vJk6e2AHNc+iz4DjimHFtfJwSjpPuZwr4tfh69ysD4/RTdrs4/BOsavXTE7k6R0yZ8HKJhRyim12
TtA7MqSOcNDMtrV5EfNOqku3q9RZm4aUmJQ8+PptK0kTRJP6jlaY3hNZtIDO3Ef7tOIxyZe9eIvj
IAIcqeYQlYWUc1e+yYwgOAUUi6196fUHUa71bcdZlAp5ys22NNOLC14dPLus6jVnRzw5+zeeBEA6
Eo3y5dZBLNoHS/3yVXmzhr+GkOhyd+WQvxLYJcxyEyBxk75Pm0HQpiqVCk8KzSyWZJHYtefndFtO
lmFHNbulWEyPOQ2md7WO8Drwh8jIluVK1ZqVxhRxc/76vDgW0iSdplLjT/yhnek/gN63aeiwTeKe
2/Jcta1j1S94Yvf1vwzheah2ZrTFonKyHBzYo3tNOiU6qWxBAjnBoVHENjAFziAzP+EyBKKmjbXV
MLX4T0JjjkuaniVPhuWGWRw1aN420tOkB4EXgcoz7AnlV37FbcltqfcQoR+LdA8RDHhRGA0L+CvW
Mmv5WjbwlHFRqWK9yeypEgi821qkTFcFY/Oktug8cHi5IH3mnB/WSaCTQlMtTNt0xxKz9xuANmpf
WpuQIiA/8grP3/IlebY/Lw0iOswQ9h8/1CLeENCVswVJqH/ocGdr32uZmG+sYJF/kplhT7NLBCU+
X87EsIYZHqVp/+tcLos0GxrcHNcs9LvOI+8R0WZtiMm33ssKv5lEtQ4N8zyWqrDW/PGRv/j1qbGt
dw8PUPz0Zxp6edBKYHK3G6jQn4jKTP6+FMPAaNIy50yt5ax+4g9o+GjY5ebcykPOUX0EIBU3GEEe
8v4WGFFk/NX8a8DRHDoYvioEr05Iap9Rh+0Z4Pq/0IvPZGCFU92b99yik8C9WOSGsArgXCe0F+SN
6DPMY9vvcN8NoWS8/9G7uJsfFgjGQ1GIqKCX7UzBYWXwuQGn+p7x8tW3vqoo0YhsHKAH2ExaKPXQ
554sruoXjawLhNCrcOdmaz2NNaSpImkYq+P1SJoyfCefLf6q3bqgr5guCdEF1WbyZUeuWqbVd62M
KJLC967uCqBSDy3TBQ/c8qXFingrSssiWuhUam4sEny+1XYDVZSJc6P+bE6mcQRwxQkUhltdUvbv
4mD6uiItjM/KZXSCjOJu/Lg6r/nPVa0IPOvqpTOhG14IpJgEYnASCmIY8OUD28gx0JWSAu81jFjx
38ZJkOv6EP2IR7hdjLhcqCkp4jnn4JwBzsergm6a7h51L8Uy0T7zkwiWlvaTVoa2FVbc1REAS+rZ
fGHS8f7eX2cc93j6GINe1dz1eH+IeIyDYXVcalRTTFuhLq8P3YBZmo9bqHHH4J+AQoU8sBG+judi
Ypn8I3D1lTx9Jzchy1D2Uv80tcZM4Nv+idUynNJv2VyxFTshlPknPl2POh2fIgAOhZSY8pFbEJ7I
4+WpY6k7E+64dRo7nxP6hCM/StsKXg0yl+fnvSZNkCZ1uxtS/PB2xBj71zu7lK9QttXyzGH60g0q
xOwflTwfmvgrObIFacLV/wbkrHqjxDGzcr11v4ekPMVdV8FF+nyoQ/LToio1fpmzJVVfVVS7uIeN
5HZMnxevBg0rehMjnpmxxxtCUrHVYYEaOBnBVhs7HY9wSpVfUWBWX2HCOCyBXHEu8TgkJMhXbiGk
UBC6/MTS5iN7l9cr3tO6YJaircGbpnTuLJ3tNGGou5IAlTe+OAgzkLqwsu4Fqn9j8Wj0HhmPYSxr
uQegJSLvLcE4aUkyFiFOhxKJStJG/0++lAeesI/s3oPpBqmhPOcX5+1FmL49zYHN04fpDfGQtDNq
TR6wJCI7o/N0O5cO9IcfT7jvOow5n7btw0Z5cne2J0xJPZJ+H9OnOm0BzT6NUvDFQeIJ7FjBKKKp
GeunRDvOVybHLBpSS6NbkydJN+qVfLWf2bc2bkn2ewcvETYDsTlfPt0PoGS16yaz7Y/U48xK7Owh
qu2WqI7ZvycH5RZIKDosA1wWK0ixKX5ShkIO6gi17Sk8T9aUY3H/rY7tRxt8I5hV6T5cnq1B+8Qu
KUrTNt1VNKsqkX6GKqlGL8RxDh3j2qbVf/LjnkeAVEKQMFeFIPDV22aRJo4SYpwc/D9COZwOjmwH
UHJoBhCeH2Yx4h8tkDtGuUJ/7iBIafL64JWTa+1JtHIyRWbs0P8X6Z59RT2QvlPHzIyBQRpW7pA0
05f4zFfFk+8hIoYGywg1keH8fdJmupTuOm+vpLM8Dv0PIDIBLh2b0C7kv8WMAYIq1MKQscGq4c0C
SHvnYAsSkgMudnbAGNxA7Ifsw0SV9eoqQ6YGlEmqWzdARUJC8TULBA1amzR99Qr4wT5IVnsCNJs+
Qhh5EBTNH8uDwlENkh3sDqI+iXoLYhDzJna5nE2NAtd+cDdfjBVAXWdCtqkniOleT86vMdxOI0wY
lI0attPmIbPQ3RxY9zj4lEtC1Q9qZ9HyGav15R2hfp6zuQfEoIfRnzrldNnsyws73WpJxO+Ol/Px
twWegl7dPbtsiyVu4cDn5fgn0h7ctAiqseRy5pvx9O9VsFUGMWobgeEz32EyCt+g1aJvMDJrm1Sj
k0EtH9UfjhH9R4QpnMynxGu7eTFOceHgDO2rVvBEF48a4J2nejQQ1WuR1iHIAfEHSuNRpySqa1H4
JfYeDuMQ8CMJDL12sbWScJKH9ETH1TCr6zxpj4GjAYNZ/PeJfMfbUf1aNqhxf01oPWnHDdihNozl
/69gyJx2xQNHQRSBG03Td3okyb9SARaxdlcgaE0FCBZfBsvzc1b3Jv5noyjUG7V83kXhlIc3XsU0
V3anywd/+l/TqHEbY08zPPrgKBbvLtDeFnsckj8L4a5TZ0FEawQt/L5t7Ufw0SomK/NOJuanmYlT
xDKg317pGik5A8jIzEt+md8lUKFMJPgSnfkrhrAoMjLtHN3sZnGtP52cvSl8OiBB5oZW779qvxhO
7NUmCwFb273RD5HF5+nfwhzdoVDBBZLxPcY0274YGt9M3rMjRhGjwLhWFmmaGEv2EebiFP9bTT5W
uJnAyaLwCkQ8Pm6yVP2VaOckyqRGdp9dQAtW3RO3Wcrwj+xDPQpNWcdrfTmghQF/s99P++fHJhpP
6mNsgsx5kCkQoJJnP+3TGGoJb86YsMLqbokIoCcsEHm46UgRyoDiPMgb8Uxtt2RFiGeamk3sn6Ph
2KHCkj+tpPaKEQ7F8zEKOn+JmZR4bXIwhCjlLCU86Qrw/JSBF9UWByqphM7Jbplw8pINLk0fOElM
OJrtdcZRlC+ip5ra/CyUIeH2g5JtrknW+d4u1haoTyy11HOhJQYua9OIUshkA0obAJH6NQWJMObQ
eRdBI636oqNTEqPNKhENvZnllu0+QkizLlv26flq+KHUOmFurUzyxL4/JBqU4edmlA8nfTIaSzSd
/oZleAVqYIgoIgkM2inz/Y34xEqz1ls2StiLJZmAwczVsaJEO1STN6AWU7NQgcdpXcpFmgEyTDuP
p1ZkpRjanAiLI8dydDM4BPTkaHcXlqb4tG4EF911tqSIimPx27BnofLoVuc+zmNd7Vt4tBzBwvRh
rwKiYbAXtjv74/zR9XKVfOHImeg3U9Zv0A4O7snVGnc1fdRwOAvI6iRZo/f/TqkS8GpnfjDGag03
k2FQOWQdcmI3fBB4TCc4olSs98012O/ad8AG5nbHL3FgC5odQOzRo1j6lxN2fBRYnicRY8WYgJFH
bpOBRb25+6rMogIRE/MrYzrQ4tpCFPVI/KqCZKdEDGOVOx/GoeA6gxRfsitf+MEdP9EDNXZLhTIU
mJReJUasd8p5eUZWwxAnuUZnVfbjT5GGtjGS7svzrj5gBNfzumDlutc3i6fZWKvgUEQbnr7m2fma
I7IClQluPxpE9lpxIwRc/ZNob3p1sje45ttCfVywmhK8pyZHmQsP2eHWXEKEQBmF8H+hPZyBBVaw
0Zv73KTPxhdkunMi2tWBjwoBdDzl0JvbCF/hzL6GxQW81juu3Hnpw3PDAIBVCLaWpf/GcermnmrH
J2YSEs0NLzsfF7JNvg9XS7f8SUCOA6IWH3aPxzkiQwZ+qEGUR9vkOWVyOSjmZuY47cg6A58FGsES
9pO6o3LV1uA5NJ3ksuGdb3ZgAKxvjCGkmcvrCJ3z8SGTfiOBIahlBtp6J0Tm1z6V7mOidSgKDWqs
+4ZFwI3hW09W8/OXZ6lzRjIiKAb/2xKrUzLDIbkiGdev8Y/+xw45EXNiDDMXpRCgmuC1JqniuzTY
4cvSR4FLnce490psXv2wUtmMuFBttU5ybPwk260UYG++mWCPTT5KO0SeUp2rdsww9NlGTqN8DyEt
InVfAYwrkWr6Jz/OEdqrea4OT3IZWLSlCn2HdLmuUviK662ZjmZUjCMR2xQ8yMGQm1kLs5xwnE1a
H8UHNJfXYzdNB8ojgh1zs34qM37FrJDwXW3gV8KBirB8ri1k1KX2IIJhCNfkGUFKuMd0h0zVny/k
o2YGeJMzd2JLit4ivpjNsdP3/ukNOkhWmMzaMbsktt9ngC3YTPucXadVKIipljF+Qd8mbIT5xr7r
n7XKHoBhHfiOkLFPVto5oFqIexjzazambqx8HhY+ejsZq4dEYl+vNqYJvkY3t5P1/E1aII5R+7A2
gnbKhsJnICiOhpvYdDSuZQThIAwx4dB39HxBMrHLhLHcV3GSdVC98+zk+06D5MGregffj6UrU0sb
s7wUm5kFQLqIzJSJXjVXONSB1q34wj4nUdhVTRuyOeBL3OwwsFjchk5LnxBqoLgK0NJVw9dpQ1iA
E8eY9PjFUIP9TjtLAdU0niUToqkdotoRs9UwS8PWd8vCRwh7RyiIeaojtRmZXxdu0zk7O79C0VY+
AGmYZYkWvpvlbyP4xnwxnORgQAaQSrDimigIdDRqM0AvOK5wuW54z4/pXkjh4ekYILt3fX97tLzR
Cnh1CPHmI6nXnYKD5k7BP1h6gsTkTxyTPVQLJD75GBYqqtahOuXLUUWdwiO8+X96KCWUP+5EWnN9
eA089MHMrwu0ftTA+xRaTCx6HpWzmesjWarJmNkAS7LXGRRsM2zMMUgYnUsAlBNGfqwr5431VohD
WMyZbh7/E7xKHmvmEhgyvg+9DZr47pofaOAp1oKGPyjuS6lzKQxqYjlxVfzT5ZM9AK/PdB9uu5eu
CZylr1cYlfcFHFMJxyz+yhWHKagJJfdhkOeEhXvQcQ8ZOrGZ/SE6BdwkAUZLpBTsdsVStqyE2X7I
3Fxqf6XnE5VYST/5y6trFJo6QbgWOiDuWm1pcvvKTBEOHu3/t+1YFnTZgKQ8Lt/e8KRDE/rVqjOE
1d16Pi6qR3+APr3Ut/5I1hS21pVXQNEBHHSDWEuX5gL/Id/V/Y+8HVfJ1I9pQuHSqBGRGj6j+yPj
QIoBJB9JuYlCbEl0Bp+8mRqvlY/rLviq5nv1lr48C5fBNe8ytEZB+6hDLJsY0N18g93KSYLaQdPt
D8XT+Akot7l0WxSJZWrYp3iSt09SC7cO+H2YBMeXmBmxAJbCKiEV5suuZvvbV3c1F1mrlawwpzR4
m2Gfw0zriTm1x/NJtMcCP1Q9h5vOoDYtZ+Q/66voKllL52MZNKa+H692kHnOCN32fu0bVlw4c0tZ
feMiyHfsa0m7d76coniQd+Cqa5jdz3gjb1F0S8rN0hKWtGnurrY8dbMJ8EcMhiWlJx87sL3cnyVl
MDQJijP1BnIjfYxQAuBbKFD3pSD3G/CjaPd2rBYT6CBpucpIciZW71HM108kg6lnEbZ7NLKSLUYj
jrJbs04H7AkmBfOyx3bnJ7kgKNyb553DVGYjjV1ydh4LiVGdGXcwsCXIB9539hlEZDOjqfAowpVe
JKqy11/O8VmML2P7EOPhRmdUEEXH44AoFtw0rRWKsP+Hu5fRC4etHusM5gxXCFRNIkEuHIcEws0v
CObCZRLXpC67FPjyUPSjE22OBdQ53PG9S5UW5FGHuF86RI0yGE0W7PHh6++KKS4667bd67MihLyG
UtJdMDiH7JXBfKFAIKVsENPURIeWHT6ebNZREFTeNMtFPmwMVFVZKlcje0h4N0I26+LSJ7Gi4mzr
ZmPgO8BIeHiGDiM1CkcZLu8CZTswrVlfbhdR8/c2WRlRl+jQ1+mExPLsvfGgC+zXt4Q44Unx5ToZ
WtjO3RJ/LUZ9gAvxVbXmPqDT0vubCIr/kVcB2rHIbgWMyytN/ZspZtdM/DUkBrUyMdsfunFIKSXN
pIz34CBLC/3FO0DB26Qk69wYYmJCgWKHT8amk54168VqCQhwlyVkwYMmSj7L4MTRXZjvyDGI70AI
GPFEi4i5pTGNbKJAnkORtqPPlB3BEKt08qospBSNLSVRmgNOjBZGPieVsIBDvrmTyBETyGuigz6u
/RJ/uCDqyxHlONQlQKG6edgftpzkh2PCmnNFSFR2n4ZsPSMRJ/U1x6GRY6ltBUuKsoFhGQeaZfSG
UZgKjuc9n3npAl10ZXeZB/jHEZDDKEy4lp/CWNLLGcQBxqHNd1+ePPIU+cgc0Skbwx5SBhxwGvYX
ARxEozU3YN5NY0wGybvPGV5HEthloi1/XlSksxJbc9dCufzq6Q41KiZYNalp/ckth+zEGC+ksThw
RLF82Z5hm1sCfyUzcVZahSe31ifUHJ8jrga4GNp2xcxktI9+g+Oh/YWj47uPXXUbxN/pxR70LY+D
iapl+ODPyeX/1SWtrAiXbamB/J1rrTG3pH+oyS+tj12rzZ8D9Yz7NlzJK2BudRNyK/Hxz5QzxvXJ
o+/ZhFBLsi0RGaS+hBDgtd4+OUSpTmqTOgeqK0JGPN8R3go6g18rKPkQ4F7203UyuSpZ/it0DPmi
mi0bbmbetM3YhmS47Ic0qUGVNj1qbEbw7U44JGZYRsLw/fgUJhZc8SVxcDZtk7s55c3mCxCduLUZ
+HJq/IVaVR4OmJCEy/Zp/u6rgKWNllrGhEXGGS/0EW5m8iiELD6Hw5YrORGYY9uxvKI8M2RQm9fq
boazMYBSI60nJvvFh6KzMGXY5TjgI6Cp9rHf4U/ozeUI+5Hyow0y69XzMw7GnZquXJ92CIa8h1Mf
EWofc60U0C2KV5z88MBcN6G+snhuRXleiBWYekligbXmatRKtBQ8F9Nvy+DA2XHcJCpdTT53n0iZ
X2CIC7xB1ps4Pg6DMcdZYrAX76B2ngi1txdBZPs9U5L2YVzojA+TYOgJrM0lGgJ1wJSqygtllqU0
90bM7AxsMl5sdDMCNTwsTIlt+W3eiLIqywUN0wXbSNoC+nD3L+0ozPHMHYnIRk0F0/RZCPyn7meq
a+SQJRFyDDjrlxpxOQzeY7YeJzt5wQ6Q1Ib3fqKNT2RIM4Wd68WnV5ndUVd4Fbiks2/ZgzwkgQy3
YvoRlCU1FVmkabe6EjHt0XisGaTOwKw+3M8JuaBu6jXa7g5uVP3/uUj0SCLLTlleszzBPZpocTLj
xlMvWIOQa6VSYidqoHL9dE5//+2yIaSWE1PVjvG5LKvm3wxKYg+u2BLfsTQFU/4gCcpCWVvuUS83
ZbWpHi34BYTJcYXZeR1IiyLcvu/9TKVzZNznEvClgsDjIz0OzIFezXiNkNv/GAWjZAILaCLXe/ck
tf5S0aFlWseFaNUVBYc/7e26H6uDaMVg12YU6Fozb2JqrufERRUZyeZFjlr/1xR+i5tap5ixceVX
CjCJu8zYaHvdTJg2flrqxV3ZcyU/tSirj95ZdzXbM/pdf11J1M1OwW2PO2q2qUysg5cnjjEOokkF
eb9gaEP47Pn3oX6RANDRPTzPs/yDcDg8dKlWPZgW1mLfiP4XVPbIKRxtl8v8QN7DhfDjvES2c8qc
RV9hXqqrMzCq+wsP/g2jf8uwxSLpKJk8de7zzDNsyvs8Crg3AmfKlinDUrJeYfFXeQu1ps2+H8xK
inhEIN/DA+IZZCfkyTXs/O3SxnDVUnWann2syaSQOBlTmAPTtrtshzfjAg1B26CumzHtyOG15jgS
/X1sPno6YbHbGB1Nsdo5y1Vs/vGqxbU5PeqZ28qqAYsp36JT7jfpS3eSFh1u9k8eBY2Bg5n3Jrl4
WKJAruIZ43z/ierRYqnMDMRbWGDDqWshXULBJ3pUauac4sB26nyggPAz2FJMgCavL42/ei2z1GVQ
eKTTSRXsBZPQDJULCRYWTGBt3bB8W6kcbHMLZxIb/BiEmwWXX+ukwT7pFndy9Ow2slvP8UrN1dC1
jLXJiLoUY1qEY1w9XdNKpls5fD0VS/umBGuk2Ldqzg3vcwCYCTt883+cRlx2I6srnzryWWSp100U
0lgHkhf69hseq38ixDD53lnOTJEZkRVorIo7alWc9CF8nu70O1Zy0UpNhkMMjePlNz8/aLgW9/59
qriJW7ENd3IvzHVT9SY28f6XNJWMeqaIJRXoGgG5YTHVCkZ2Exw/8yFX/kGvIKVvSZY5zD14nFSL
rSREACxdjmYL7kNcR4poRm6Apq77wcKkvtwThNFEFiOnFMfqOKt5Z3uqA+1fh1pvWJHvzWGInG6a
I2wVlxtdkPx9cDR0bvtrvyexntXPcByF2mQGHxN6kCV4fUHNBCWqi//XB39Te2DQRzHmCyaCwqge
OUM7hLbySiNo5rj8C/7oKox8AU/sod5KH4P8Jsksh7eMQM8T0ItmyKmkOuSmR/9wtdgIkECOcj/w
WAedqZtlu3bQVncnTJA0lBpgpYxsXGB7gqQmeCPUDJmDkO6lFiTkUtJ6p9inPllOHHKdjdLqt0za
1HXUp7zJgnnA4e7pdk+D8AiuuyOrkTNs9Wcwzs8xdxh2I4n+acXbLl3DRAfhYkuwbyflAmkQY8kV
5w8w8lEAau/sk7Pviz5UpVcwkCUd+Ux+QzksFr69oNI+F3yLbkZRdSsDZXEHGsAmV16axK2Bw9P0
Q729kKXe3+FL6IRoqMtHBfFCjVqWd19/Mht3xCXC1E1cqdt7vDd7TLYEBXQesVH7CaM5nq+DJ2L7
cq+cbf2iKU4s/67gcOVXNSJjZuIou613UAssp4tKUXqBTuqAsmsGZpH+LYeujgDWumHGkNCJL5DZ
OpOtWCGXHmyG5V7jziDDOTbVCq4Aci70umgE7sYmxwysjN3WtG+0r8FO9rKbO/A/IIpXGmAJ8FzD
idIUQbMeHjofhzPosUGwoghvhz4HDI5QJBYH2sf9UC30LCFRwy5+GR63Z5zOfOI1mu68IlcARePV
vUMWqaeIZEB4bTBH1QB1O29+IvzoiPZW0jCBK7IWRYpSWunT5NchlRFY3JULG27ZvVQDFC1sDZ3g
DyOo9zg52cgGw2bO6oKICGVFPYcoIcSFHcSt3dfVi+cfnr3GHD13T1JXdBW0pnvExx6Q5FhyZ/EL
6ov0ZjMyDgGxwUA/ZFDZ98V8+RUvCzVstinSUZaTPEScJz7Jy3JOBfsSintXn2e8YXlIIClQ5yai
Fwdgb/6f4oMpB0sfEgqOG2lDAwXj4cbZQylt9Kc8xiv6BBvWHSReDIYMtOM7sp8TVtwche39V/g8
c6giAWliA+YKvfd+Zq0fAxnn0O6GQ10PQYm7/S6+RzJABA7NQMOWlC5GCwmr0v7psFL8DnaVQChz
ST86npJdLCwddWtw85I8dtriHcKMYClEQ7Xsk0sTMDGJ1ZjIsxUInGbkLCDXpgPFowYhBgfG+i7b
VLIhkegAc0uO8lWTp6tV0hi9Qxfae3hRhERnAkS77IO1UrircJ7wg5JWtI2wbtqqGvzWZs7iZSve
jxOH/ZdYLfdgUrA8z2uOrjCrVwHjUV2D/abSL9v85VrvbPWcnIhz/cV6jsjhtIu6pDYUssV8zTMC
t0751wPJr1vsaqd5XQZSqG9e07JASrFWZ2/sz6pSmoJ1zRbu4jWi2Ei9B6wC+iVG2HBBw1pdKhDw
hVuAcLdaKm9fQcMEesnR8eQ0GDXFWOjPeZI5IgCTFafGyQbcdWxPTAi0VvfgulzHqspB9woTrxdS
7npS5lfsRQSb6D6t3qlEotT15Jtors+YFOIU7frvMYoULhCVeW1LBX2loUmK6USFY+qmTx4cgSzE
ExJ2ru9uWMlRevjj62cDiC7fm2fyz5TcXr9ESSTpvPu099JaZraBLDLmsJUWd/To7UWX0sB7K6++
7FsMhLrMD0dx05eO2DLuD5Hs4zz0ZOPK31tt+a1G3MxxcislTQUB4BxEKnQY4MdPG5terdptzZNs
mkkHAVXQ6OPotKgKWBtp84OhF66T4dPFDfekPZRRonlEcOWQjI+f5rRrKFUHSccYn3rLAmrymAfI
IUBcZ/qpyDQ0b5Y0twEQt1S88+i7p5qQm9qYaFFkgCvNe4rU8O0NoOs9+39G0hMipQbv92r1p2Yh
6oV3BtTBWWn/FWmjeBxGIfSyGdlJSJB1jmtCwWa1uI/ihV/fEFCqhEY3NzXI7PINfLjog6jqPMGN
UtwhIHHXykfjbfOz2XhQCaWuRMuixoKYdxYEi/o40lXkAU+7YRFjcVs+lvxA56AEyyQswddBfQIX
YuxoKPF46z2kyWAQrH6wAdV3D0SbI/XgB6rvG6llqrLxLyVMlLpNSpgCkbLifdQHEmN4ORaCb46b
qCTPcl2ZqslPJmhKYtP9B2Xf0ApEfIfd/Hyhg8iZPt7ApfNlu9ykv7C2A2gKA7MNgCrZ1lIZol92
LnGjta6Ay5h4TT19tBlJGeJbOlNTdkyb2d1g2uXT+3wjvWSMZEZcYFBFCtbMK+V7O5UpYKxorH2i
BlKNyaIEm+7X7LRje4iKmGbTBJDzOp9xmGZD0hsyJlwwWmsmx57sNnLflecCEc731+hh50vjhe5z
6Qg2MTl36z4F5PySryHoPIfkyQEAEUII862iTWFFo1Aaid9r5nwVa046qT6PNb8sTqamaCDfMBe3
ryXB2DvUra35IYiIQsOc57+uy5Mdp3YNHthfZRZiUmnx0RpIUhnQCM9L/dAj9N9ejgWDVgIRJQal
T5jlU2BFPDDrKONR6NTcOwmurWuX7CUaSjxwZQlfbYtYN1eKaNeVXejVzchxjTT4m8WVNOQlV/BW
+G18aXwxXmhb7z81dqW00c+KkMm31ejqgJa8XmcQrn2iYVOsemF0IenX0QfMg/3cTSkI76zx1T6U
Ak44zTZsY6Qr0SkdeDEuNTVlAe0MJF9jAMIK7ta+W2IWM6Ei4JpYkUVHUdsZXwWtNvMHuMcL1e8h
RfxPUBD5jHnh0Wed57hkYNQ778EpEKUBFM7UiCMsW7B/LDyIH8qqNZquQbr9slocseAxFGW1ZV6b
ENQsmpycRtAYS6JPusa1Kq7lbN1U3O7nWNbuuLqDTtyaJ2Mrbg58bGyxmttPA0ukEGqMEWYHm+d1
AQ2WA9svOo4238VMkNMTHi1fkT6RKHnvTdsmZ5Z5yeamGGWd+IoSssO1D97umo59CUtNnbXLxr/B
Ip60ssAk/gQa0XnMRzS2TA5HvgsHgh6aPoQENQ2e4ukLGNoCcy3BOFwUfrx6PGdHnR+cTKRN+JRU
YnA1cMSZ+IMqGiyjak7K/0d4vx1QZopVCzVn9FOQH32cGhn0oT+9OdrUequteGcQraBk1tYC9iHt
b65PRxMDzyJ6zD69EpteKsu4SpC3Q/u9J/tf34M3M8YRRx1xbpFZd4GujSv3zWTyRcL/xkvr4Jjt
9+J/+2xobbji9xNLfrhIY+z+7M1nK8F31sxvzNSqIdUl/YrQx50dR+bjN4TMz1mMU2Y4HugxTyaE
A8WHgd3yqbxuRLDKJr3tVVGA0c7aOT3SFMf+3UJwSAwjV20YkJyISRxS9lA+dXMGRITHyZ7ou+ba
1y5EigxRCr74o/2eDW3IhjEBS4BMmm8gosgra98YpgvwpS9Ab/dNJcNhmDsEema/TnIdRg0BQb1i
atKNZkWrWXWvoRzLtWCV1CPJFGlHKyH4fJ65djYxZI5ZqUNwdNexaJ+lZUWvbKGK73DnAHX/ZyW6
4ZQdce6kBONDmLZKUZXvVA8CLt4/XavBPRrBoqZdKLhmkqDOb/bIPHFRu1eYX+Lzpbl5wPqONhyF
yh06ieK+B5osRRdxZh38jpRiwT4QHRWm0Wx6YOK8rJnFkVyH5gSv6Q9KFBOYa3QNgyh8OsgLOeRh
ZbFH633gGBheqgz5tq/+b5zcIP5dDKNWILnq45q0YHtCO+01gqsoGgHmhAez4D5bLW9U+1yqirxU
SXlV7ukNj4OuNn/w2WMmKIsDL6qSqj9RjUbuet2nsqlRZWk53peRLKGA5TksHow8I/00JelccgJU
VwVRZeDE3HEz8Uq+TenjUnceOcpxRpBVoyd2UV2JWeBZZHxXlcrOTAoXK/IDFIh9KQKEagBC4JFD
k7O5DNOhXC+MzIi2y3l0SVUkF85LX6Fa5Eukq4TqfZKG0SnFLjhmvZwLuaM8IcWnv736RZR6M1/f
N5VZk7Qas2+CDzG/PR316GWSdj4+GYxQoe1QmyMG0gMrYfyAU+t3xvOyDA+mlNjtiipJw33NcfCT
FXpeEbLe99s1XXPcod5iagDdtSAbI1t6p9sH6/a+D+ekJQvyqB3Qp62s7WZVBiEwgJsD+EzNNOf2
F2Bs7EoQAeNZ6DEM+7hDSKaTjh9xWQxa5Q/OFj1XVl7vlav46tuKedpFuQcTayfIdCH92j1ns34Y
Tzw5YvQrBKBmyHr4qoy8ctRsUh0mXZYcaj8dFTv8X2i9FXNj0u2LBJHaVjkaqX7gkcL3hBfuZWNJ
fqNJavZg8F5Rq3cnHhaCvZNiYFmlGma657JC8WlxwF9C0polUPnY6H7AKIfjVICybxpGNB3NVxda
fuw+8QHmEx/76kYX2daL1+WB+O82ZD/cHlfUmz5pxdovMW+ImErnzgNe6HXKUfzATxMYqmHubvA9
9I+9tBPgZnnzedXsEJe0+89HGRuzrc0Kt0D8xCkfxU9Qj9MB/Ka4vp4hdp608m5qh2oWpAY3rHmy
F9meZivpD9JIdOsa99IBCtxDZkgUIjMnx9fODZkKu/2LHRnGxkjVzuMpUobE1zw88XqoDjEqQNKu
kgf5k0emppaGHegUi2rBkjgD7H234VpKw6mpWqgvKcErdSLVzOZi9JvHFkDYG+44DdYWEaaULb56
NKzRM0YRAzIddugAwDA0RhX/GvDLI0ilD6z8VwKrCNY7AazOc4rf7531gjw6xc0VzCu0ac+CERsK
q1sMdElrVIwP6CqJ+T3+IpElSkZSLd8wezJ3UO8o/4RjmHe6F6y04dYJcOpv6jge+bB4UiOxMroq
6AYtEBAIzWS9PXgQBzA2NXJqrhz11qcKhbm85oUXbhAac9PZ/LMXBBTgWfnwQiHxkT2too6pCG2m
ygS1j2McBY63llsJDSKt7Qxf5az/Njk5441qUUhR6RAUUsx6YL7r2WeCwxHI/nEQbDyyiBzmkuBg
RA/oPCrADw+srgaYVA14fbICBoMLo3QT1+Qmkv2DNitaUY5XK0K8VH4JNOjPA1nZ/gWmvU8LxTRt
GLHnVo6W75bwy7TdVOVYrv55AgC651c+UGoKlTpl02Wix4STLhar3jKhAhkCymJftv6dlLuMzGwb
lZL9pHoBBrq5pPJb5bgidTHrjjroAvsLgI2BuU0Q5NDKNLRr+2XIU57GDbEZcI6MOUUHB3fKGZjn
wzdUwLXXJWuwSbea8B9+bUHLLvl+ZWuloXIt0FZ8Xz+032w5weHMaAXJd0Pd27mtA44Fuh5ihKJL
g1MLHz1EdGrqEuNQW/atpFMNj73R+JY77111U0GO7Z630To8GFWsUY68Sa00HzZoDOWKb8piWvAI
xUZijHOop4Tz2fA1jOghlTfXmatTa088gJk5S4CWHRluf+CVc9iCIMl/OumQs3VomPYLRZNq728n
614VPKGLXEcpDfmhq+h6Xu/w6qmag1CqP27ycOhnUnPeu6nJwxJ67P3PU6TMFXPkoiKGUt8seFVG
ndntOxl7X7cTvSf1xXzHXWpyV5Zk62Sc5YkYk7K3wNPS8+TYn9CvcBbuD6WGPyaYy/tuDd1ci9fb
UbbwVTahCHg+LsqRCDK9IG9p+PLp2q8Uit7U1UQI/5FTVnsQpQNBLDfVfgVNIYLW3W1VCa+6Lqi5
Ieo+Tj3ixFiJ13Xrq/3u2LnjYj9fR45xSq/T/M8AU0W8zk8yPA483QO1dChJY34wGcQ2FhQL+wqq
VXxjD52EIDbBxg0Fe/tKhIRaQTjngUMkb5aBaiH6TKeaTLBUnnmxG5IKaAX1Seyh9V3BZVDkMovg
oXr30sBI8xz/AjTYMkrswRfBlHrpwVCAoHzIjJvCk93G67rZ29EPZYezU8u/S8yPatpKnEgtNByX
dThgXibS2Sqaqxra98Q+R5NM/KZjn/O9Iyx+aXlbEt5mSxDYHvqJtpk6UK7BULAyl5iTV3xKbGtv
A/Qu3jZSgGFno3NIDkTB969ARD4oEZ85JCE/yareWBkPpf9+UG+M0XYd5W/4bX4USm/z//yV4nUt
/Yu04bSLHCJJTpKv/v6YS9vg8FY/5Qyt618ZDgsARNMP12P9rUfbioPBDfY7uced+47ydm+mbYNa
134CljUpjcBRjgPu//FK/WAcTpqIAWfG7Y2bendOWAD33QUGxx9tk2FcoZwd0smnWxfUOAUBoZS9
U9TgLmzK3XLTYopkCILAkfdzpNLKvs16ywjVDlGtn+LDaU2xXaxJv3h7G4tHSxPcDwagBluG5Icu
J1gXBRC/fvS8HTzltyCGfYEyHRw0J6N/GavICJDGq36Zwiqo0+E/amM9eU3cTGA48gitTNEVEz+i
L0HoGu+6kBotM0dH2tEPyf/JGe6VD+4tIi9ksXHyxCmbwlcZ1Sz67avEgqLRI3K+HPhe9lEKBPV6
PyrH7ZnfhY44s0c6xVDzs1QNzBVM7NlV6oAWwZVPAvxzgh87dEg3TH9HLFl1tdONtIr89bTU+tVP
1KXQhlNAfCgSZZwPzYrqYUhZyMeZMwt+W5exUzIIXM5vYuMXu9qC698hBEprjLpvPQV0psurLrIS
HGk6PX0SNNmIvIh0A7ZaP4wv/+lym8HflFKaFwb0h8DQMkmNmPYX4/lBQE2VycgNaFs9TxjtlThZ
Hdq4xoRfYTZNO+RIiqaApL7qX0eSIGVDom5GRg6SlxtPtlvhji810EMbfIfYmB/6s6lyhY+9hCk8
qzQEK8MTcIp7CHYomxoQuXh1m7BH/hIrHAldm1z7o5kVqvdaop+IhB3rXitzUSjxqq1W1sPtvoLG
fZIx+0zZsfxzQSMGuZXQ2yb0Fj14jrkzLGsLfk1opnzGSvbMhowk/PSPtKPsHEw4oXsYv6g4NT+L
OLYIqXF9XmHGkfer5YVX+cbOb5nckjcC9iUVGFY+mYeOdWBYyUu15xmE1xO//0Dec2uQK8TFtWgA
ApX+n/jYr+k3rUipgyKqGXiDB7O4wNI6b510UserQL0fgosQVZHKnmGu/sjpw6kbVMxo/1h3zhtg
7yDIvZb9NcsE1etP07GyHGbaXpAQfZp4mSHGPmw3cl+bVIxuUMM0OecZWBFauDVe2dkZf5Ga5jVa
b6cUfFzsOx0AvEki2kPj9vc0zRnevvdNgopyNeK/39bnr6BEYThvhv0mdXuMk/6RxizYrUjRfr7L
9FHEYeVkVo+rZog3hbtfjwFSf8XZDC0sfhk0Wl+HXhiLP9aVh5LolqRXjhu9dnK+nsbgCYMeo7gh
5mUAjFUtoGlnVz3NFbngMzGjsby5Ve2dcxvTWFCHbCfVs2p5wiTD86LRHc4wHH/1HQEY3evt6bRs
Uvdm+Y32mlRAF3Dt7SWw+qupThXlK98DSjLCeDm4buzOC3Ny94WsHq5PCVMuH0df1EpH24Yeu2Xl
QaGWZMiZQjJsYcoo/KhkHiU9geB4HAeEfVnoCD0SZuDAl0KCc2NHoc763VdIEBLdE7CY44oSnenT
IklKauQiYa2fUBRclDIsSHgXxXfBGHcSwqkG3B0wZiUGD9/hpmsjHhJSpdS9k7E9RS7/zTk2iGt7
QeVUUip15FTCpGc8NOBUmY7Nzs0X7RanoyOM/t5IiD1Go34QBUiSeONsnUJyKhzli907YoO1kZBK
t5qilZc4fjaBDWppqtJsXcrfBgQE7BxjAdCf/EOlqGQOhq3fW/v4uqEuMcbECZqV3hkKgQuCNxnV
EyTCtpaGEp+29PTM/d692PbC/uN8bF8bfkGKHMUmR9Q5velc9+Pky2AIhMloZ3GIfrnAmFjq5kfm
dso6tplUdRb6Lb0GyDouSi+wAsMU1WgRwk0BQd8/++MSBTt1potoYnlAT2U6Qve+k6KDThR08JEB
9Nd8iZgleZXmcTeUlLC8gM7SI9l0JI8p121qSn37eqw0/DbbBTV//bVDoCII/6fJCDhdEV9wzrJm
wRt5/9vCjmUOAWKl5EWdgOexxxOH6r5qUHAeCsi3L3RbOuPR0CEqZSANUVQP4woRlCkFpcE5FpSe
6enHE6PjNqVvujDLHhn/xUEOTzreja7hqyD+2Y0krKTGhCtGFVeMXO7FKcYsBJf2aQy+ztsuttpp
14lXqL5laZ20nOjd8jxe3ihD8GWm8S/AkmsQSACD5Sz0Tr9CZCCSQZeAqDHkqiRUUBQEBXi3apgs
olFCGP8+l1cpaPqklHaZf+3LEjndx3SbBuOZRduC7lykOQ/KRpMcKtH7NYWlH6HdJt2ZGBTPPVaS
f4wNoI8rH16pBm1fN0s3JbqulHSlOn4Sm6mWfeO0CsMkfQCaA6biFtVxWg40wywFiKp2hjdZlT6/
bQeeuYXhjbKHKwI8U7U9/H2vPLnZXMDl0iXOSFzffoL6t2gpZ8703zMZ2GXgGKadPd3Ehxc5tklK
ngEfBMdk212WuoYUPcSMYeu2nPvtPezvPOV303ZmjdjROFZrlYTY5Em+2k7tHzimSGoia61qiQg9
UxveaTm9bxbgFXlU2HBZokYGc3YqreIy5TyQs7sYv88lLO1jYm0yLGeRXJr1yF2Yn9V/Rfbh3ssI
Htn6qyZMzH9/NonPDQjwPLMnR7lHvnZu6m7QwD+LZTeM+232nXGjnzX3nsPQiW9MRnctyo3VtDMC
eWyL1mxeV1J/KceK5fN7UddeHNptiORX9DFZJHwHxeOHLhDReo9Hz8kXfMnBRmKs5TditNV7Y+EB
ZwsMoBm6meubmTQN7mIV2ND9hPCHJec6bFJf6LPejqBSCuZBP4HhhfN/HsWe+TD5Cd5Q+3ecRCKj
20HEyRvtJV6krs1NLn3MKJv888iR9K3FLYhqrWWv3eG8udrSBYI8rx87S4l+YBvIYIRiTqboao7r
tJ66DA0wjfzRfwyKu6jWadMhl6sutJPRUdf/+VXUDy1FAyQ0AqPScd0GaXjtF4/LZhuZKVpvFruH
H0yM2GbICae3/FOIfkpB8Q7SxFFJ0g6pE39xXb+4DMBOwc7TFQjiME/b6tGOyv2tGmglfvZId7jS
fs547bxOXJ7SesIQB078mKKntEuLmZmhiVjmcPcEcRv6h40VFKOTtt/gdw68O45JMWSoP6hSeMya
+EmFbOKN6UC+nM2JKRGJELleL7AxAYE/BhYF2I51/aIgpQJhgSX7ddmIzd/ZZkneeMSUpemeP00w
9Q+6Ue5lube9+opUdTcjPLgHgGSCf/yfl0q1OR+x810KrEvey7n8PQdN63E0OJCgjFZKS7BCsb4y
41Xql4Fdves+6udNNX6/72dJWw7a2uRQ/gfFB+q3WcwYWxq6zs0xOgknNDVRP77VTCMkxDit79ZC
eR1LDD3HJGbPQqBX0sYbc4sDjFhPQ8SU5PZVCyoLq4Ajl4zuGaTrBROlQwVCDEq98Nobz/q8o7+Y
Mf9mOPlj5Poan/EJWE1PI4ds1b+C1C6mNJXkIR1N06gjcPRKfvBVNKuI75AtUE7yqEBzP8Cy4YA7
tPwIzoIGheD1+wFq/uMaxyXK3L6MhuGJxDM1+wCsY2IO2nsmytDmpgYtTjVaj1Zx625l1i6wGu+1
uftQy3He1KCEJBHdD5GmeZdAX4OUlYICjs/HWow/EbnnV09JCnr2luXrbdF12BPnesMxGXGhea/v
YCbEgv5ooogB3+HNjtwogn7xMmiIlQ0HWnTAU0IubO4gfwwF3Bchx/pX7pchNkO5SxLw4k0wPeyM
F/KUNaRedn+S4lvOqMP/SSKuUvx1S5iXmDXByuwMb/QduxcYwvPWBAkutApDTV9IXeDMwD1WpH4G
ZM8dJTwBjYGAJA8YzIZlvRr9vYj3N78AWRY5nMRvtKbQXnBVL1DB/pvsJn3fhs9KlhppMkfu1KHw
tPdV+sfervRr/Co29BwpUwdpbKVJ6J3wEenFPNsE7KXhNpz8eX5TtZDc/tFO0Flcm/t2fFBU/QKF
1zyKMgbrby9uGFPcN6PV7eNns65FmZWfhtoaqjc6KBmTOg/detpMR2Ybmxv10wkTs1EG+KzxLNoJ
bf1l6z2nu/W90eAPvSatWr0qyhn3tOeLbOmT38snnWMHVq/FB+UKmmzM4X0G4zwA0DMlNgOoAw1v
+hDz4MJdGnQS8S5wKxpSG23DW5cOjW3ZYzlFkWO8UpJft2gzlP1C0X4lagJ4SAQkZjJ/liAEoW2D
6xxZ9i4MrY3LSXMesIDWhHjZzvsgRNYiVM9j7xTyW+XygpnJUf2aC+AxCPZzjVPSgCFvHJ5hvfDg
jJjtbXkaE6UcKKS1fFIxziPxyQpmWJw3VeS+y5SvkmfWhX9q6bb5Cs9lQduN/jmA/YrNTO/UpJGR
ZpwtPSlUHmVhW6Gtv68IxCX5C341sBx3QKbu2/kzfP50j3ldeu96aFAYTmOtIMXlCnGeIi4X+Wh+
ThAN3ZRMTO6xj4Lv+LJz7g2x4HzSyhDL+gGeZ3DuCDZ2ElmqW/GTVsXbHREoaceDE1g/r2/v6GVs
u7n4OJXN3PzzF3ispsOhB6x49BZsGgguuWIbfTFDePDB2uKkVhw9IpNZNh2KV/p6xxBkuokTSj/W
r4mWYSjvlPfwGc624/5aZiFsL3f7JzMQN9GPRhybvLKFerCcCNglzUdWMIhIzvpnf5nyRJACY+Fz
Seo9oQItYSyAUyJ+RVB0KAM10N6LRLmOrMWbLF03iJCuNlHK5w0B4Zi4zDQ1zYi8YSklJ9JhuniO
szcRoxrc4pirTEzjRyM8+tZrv3UKoqzesKzfZUxfkwCHpM36qetX+7Ufv64u55RZcIlcFGmOXcB5
jDWuFuCpm1WKavyH8AYWTpmaHVXojXSkFzIuWA9m9IOZ8SH/kDL4JWXVTrJUbtMbnj+coyfsyzqx
gCJlwx84XfqjXCzMpnkMNYNIpebHWXCTemkrxNlt8/IrWWF7njFtzm5GEsXW1JFAE1jRdQ6CN0Fm
OnVUKFmom6XWlNi77m3QY8z8KyTuQbT/pGTDIQ5dUdyF0OixQ9ii1kPaK3623JiEgat1qaZKc9u7
+9vbeJIfP0pL/U/1lcVOYl+EgEAYxLJhCjNFRCvVUblNYw/knmaGN7MCRtU+cMi57RVhBfRUK3hk
gZyK5pzqqzAgkDMoq0Tr1ci3gowWJPd5vde3ov+T0RZorSHF7aW3FGNGFqxpMilG91G4XEnwCpDu
3eCjTBmLNhmjF1mskh9mXyEykb941ZbljhkYdPr1gGL6H5RJgKfhXt6KDn7+gQ7nhLUlPLxLF/AN
0t6nWMJTUoLCFvDTtJ5o3ks9M6iGYbjhOGnO78z0Gb6Zbmf6c5j5WvG4JP6K4LY1Odx7MN99PCiT
ceImJU19SbEr+q2zpfPsY/afMHx73HKwec2RdVtbrY6sIxdwyWbyt9IuYQR9g+epY9C3kZR5S8aU
WfpOVB8SHlaVuvOtJd6hg6//WNojxdGYBZWRPljBTJQuW45GxUa2GrTTzn8XuEEpKLRZHHrEf4MG
ydDbd5IdScfw6EY8B58OdlwKS2aUfU5P8u/pd71+AsjgIlHELYymw9mhmFVG6sTrsvtLTX4iSVGV
0+C+y5BaMTXwKth5EVaQxb8hM9nPDrTv2ghLVF8BF5rgrcsL0V41h4R/rz476qZrJd3bw8kwdAhJ
teR45rc4SIDMXjGTULpzhTYu0ui5TqkFpXyHec6AerxKuWH6Q0c1n/Bj5UnnF8/fcY0qMR7mOSwC
sv7P8jLR4xau5gUnS9iLVGe0Zcqylur1Hz0M+ZKUduUE6iDZGB7qo3YSaaSfBBzTBLuTHWk4NvqT
FwCoGkF0jDD8opCHRPbKtqja7W9CL6TuPCVNd72MwdnipX2BKPHsk1ktC6s4pr9VTFDQ++sKdFBm
lv6NxpNCrYK/gQ3+65GI2A6g4GXzDGD/IOLW6gTie7pP7UoUTiaOfgCPPFMFgN9WOlRYkD9/yRNM
JqV9QOPeSZTorIeHZWe1kIeQZ224szTANUbkGC0JnGHziC0DGeQSGtDjkOwGy/DmYfNBNA9llwvo
cTX5BaHn4YIn4HNoL1x2aeiOW4tR0RcFxgZAjT+n24YWy5LRhlWcMfaZcS9e+OHZQH4N/aGX8MFS
c8ad9e5ax4FzAw+RsZRiJ3NovpFx6Kc8IguytxyN3q+ziqpeQez/XJdNLQxRs+7KNR3ys/VNcHX0
fVyU5ecYqq76Gqj8VntvVpgl5GLoAHKmqcYppx+TBBTaIZt5WxsPJ1aDpeJuvKKEiwfwNg6IEQ0z
mJJjYaYqF3crh87Va2/jkyhz2FeWsAWZl3QhAaifRfAu4wEBpmzBjVr0nM72VZpMxVhrtNjFM323
GWzbmEFj9O3ZDmDkPnktjDNJ44piIMzgGgRy7Sj53YOx07ErqCum9CY/pMmLR4IVBsQHqWcueaHL
p0BHLWcH7kxGepu/CKQ9pWZ6m5OdMOZNheuj60hzGplaUO5p4WiaAaAxgGNMG9QLZq/DXpEmxl6b
WTXOgyXVqjMxyqMbpkn0oxFQ0M6K6+58gCQT8eHHMgNw6a/rLh6p7AVuh8N5kT2/EXtfjoWZyBZs
grCrkzYjnD4lK6vn/j0xl8g3ATZB3isP9t+oRqpkIs98/z6QZSMSytEWUfS4HeEQIMqfSlIRyXvv
cyq88wxuz3PolDe6m6RqjQ4wfk5mPsURaqS9UStIksLoPN3uNtyUD4ZMV3psD/6RhahafUsb1Wxd
CA1FWzWoBRiGwb8Nle0XJC6Qz2HIpnetlThY+FGFYnCVKrZjicbHGhyJ6/6DPw8I1Oxx45UwVVhX
v1Nb+QOjrW8TXW6oPY3hb102/NrY39iFFwbjsiDZSmy9EzcYKTGAL7uQi7QdLtUf+oLM8DP2ssyT
hqDFrgSN+rj3vZ3d1IxgsagpTdzV9nBEtQja7APm+m6qTLWBedZgnFC6+Fu5bJ6pGadeDC7hwgd8
UX2pbDQBtMAtqDpy2LccVXKThxff/Ft1Qv4vqZ6zpIjRnqdBFD47VHuJjJETn41pVEsCTYYHbiAQ
RAAeiuzKxEN6tWi5wG2+nzUkCjm6SHW0k5OmPY6BVol9TSFGscuurb6ocnC3TMQ7EdobZCiQEvWx
+CvTUwclgdT5bL6O2UcEs83VPPNOdvhyTDBlsnvNMLq16TsvZhHGKMrztHc2Aa9y0+tdPWQA8V4o
l0b1N893XMvM+1xyOB/NhDghSMgvRIr56KU0YRPIkV23Kn4ll/gqMgFzyQfMLShnt9LMq5wGbk7j
N1WBhbr7RheT415oqdl9du1922T84Tb+gXiaC2xAdlVE9tqSIdCXUJp+pIXZKh9JQFIIKQm105aM
vM4bdvv/RDm+IFx3b7mQT0LdWjx1ms4A93maVBPI5ylVzyuHdzgOMN1cuWh63GRMOWeDfJI5r4Mq
I0+1cKJ+XTUF91BP4omx28YuP4+mCZUjPcFbE5wH3NrMkmw1f2YQ78YHN7AHHTMsdrhxcWBSpa2c
Met3LDmRkl86MvZ0ISSCg+2VoaYhS0vapd6tg5CiLOlgrJWw3HGs8hzOo3vmEGzHanbjD9F9dBCe
7GKaQrO4uJOEIcBWeJtbD3xeFIY9pfzU96wDyMFyxmgd4EH0/s7z4uKwH3UomMqx2GbHAvMDdcvV
mAhkImIRvsKUeRk++Yrm4I70jxMEmmfvjqzYodfbOjcKRe++MQ1nbF8MzaOVdmmqgBRCf1mn6GZk
dqCDNHP+tHF4sFtqKAs9FHQsbsEX+K2czmqlFYYVDl/LpyyQeGqa9U35Tdf7PWuFRnf2TBFjmbn8
3J3XbiIN1fktj3HXLp1O9sowlETyog4QJV3hYxhYkjK5uWZ4sXjBjUQJ71yd4M2zWynS72rsYcy0
xrmLWYyf1D3gLSrNEpnpLZoKxK6PJsVZqODEd4ujFdOqrMUMoe3udGi2Jdbq0ElN032EHtGtSe4S
ur44Ymkw1kogugkE/mRiMQbSoSjTo8MoXLJHEk310+UFF3+guRk6EsMhipnfiYXPjj6H4JP85F6P
1fWgmIFi37PFKIln6rS+/b6QBot7uwA1dEumWJq2ji70boLH3JlL6XRAMz6Z1WHTLFvdS3haUm2Q
l3sZFY54P31a1z4y890xh6CL1gY/RINu4rGSR3CM97HHq0t9QaFbRH9Ke4tEjaPpQpFZApkdhn1C
HHFZf8kcl3XpuFjNEN9jDv3hECmI9cZtMlalVgO2FsCthu4JY4Pl96liyISojEg6i9FCHgNk+SbC
0b1dmm7KflxzdSD+AADx6LKV8zjYH1860TF6tc6UueNy7XvBEJ8NYx5glWBN+pXUXGMn1sCVgBfb
nxUfZtnIoJ23HUgM4EGP2orLsy7fW8d0f2uiR2wttnhKbFJ7x1icK73mZdRSBq4YymOQaWZK8amc
OAEw0q0MlcaHiPq+xXasewYqG9iUUlgB8j3CjB3YSans8nV2w+Zi19jeX9q1OzGbfQk5JO4jvfEU
Zy7tChz4J/t07LWy0WCvUjAR/hMAgGBdOC9bcjA6SLcT5MbaKLydr45XlOyUs/2GyISisibVchdK
KneXKeig+RoUM8VU7Rqekv5lFpKQ3U4pNhs5DvbEfPzdHpozrRUk/KM23101kQBl5yWXTF8LeT/U
V0JVJ/CgFFAsIiFUZrSCSf4hlXWk19YpNem16VH6/2di4MuHixyWw0rtLrRP/7PQ8CY+RhgSUXlr
VGr/lBFcayMEm6AWD+BI2vdYW/ioBwjAIRSTKkscFyLHOkMPbWanVIA2LMeQYW9nDXJz/Z6yJZaN
hviyaSA/zixFcekwVokRjGX0Q+WbCLiTMUDvdi/+s1fZd0emuHThZ6Zo90Ao4aFbVqzRLaWBC5RI
0LpVnFG7I37M9FRnFW9VooVFO107HwSn+2x/Z0xiUEc6UAmFt/LNNl8OgkpQ7WgmVnVuHHkk5ZBY
WmRg9fIOYZArlvqIBHYO8Icdw/k5DFutNpPDhjat3JZInHndH+WrBnKibYX4z2i2jfAtqrbnl4zd
33CEzrV+9jQU2ooRRUYdm43DXGK3oW0cvMKl1p3fALcaUsIUKQcG9qwSh1agZMfwxfGfBWAPnaVH
b0yY88W+Cthmw6r461M7MyxqUeRUqjOmsFDUBWgy4IRE38QvFVwZZBgYQVHxgQx6rFIVk6XsN5iF
xb7y4Gdudp5+worVz8QRpBRtTbAxIK51c6NacShymzZECs8r0V/wNVX6is8DBPELd2mY913jNioX
HCySiWxD0cotoqx1R7AJQxe8/6HbgnwVWGsoBJldvVF1BM18aPqJnsXjKXPqUXGk7COCTPY+LP8U
GKzGi868sOPi18ygJJhYuL7/J1zflsZghYYUMiwyNf9b2A2tXISnv2GT1/WQzCoeAgojJv3YODbk
P6K34F4agy0s4ZI8aDTpCNoEpQACbRgBTsfO5GgiL4b88LC7w7JZOLoR/szS8i8qgojm8f64FF8r
U9lpdRxDVsLHfTzx43Mty2rWHrH6cyD75oX50flHf5PJTCaUpwtDmcguWP5+zAno2hoyzc4Z7Ird
/UUXJXE54YxmGNQ6Sk3Cl7FC2Fap/WKucRgu8etq+RIs+upnKDxF9vlJ1FtTmzfVvLx4ceOS60tz
5LDFqFBH5qNiTZhET5NowF85G/GydRg678dIQExNT7l7F5VqKUCzLmRyjcBV84y73/Ut66LBmqYb
AT9R61VjLiYozBv+C3JSOeyMKYmMw3lALTDWNjBqWpqC3NSpYwnTQA8x5/AVMaYZDU5vXvM1qBBH
D/X9lbgBo4cswGi5XKem8vHxU3j18Fme2p3ZVnPM6Cm6TEMVXjdNukFCdw/cf5f0NO6tRDbfPohD
fgZdG9fzojrUvdiQfGqC6XJAH7pPCNkvH8XaWl87ed53BfH2Oj6r3zP33tJkRKCg0xFeom9AReqM
Pp3YgU9+XNDr3UHa1bHZACNr9lhOL1u8ewyIplOWZecSl7TpGukxKu+xEsKIsiPifgP3yBwUFFEQ
L9pT1LkAaCGC2tl8KopBxxX/bIwFggJjEDkp5UX/EtslpWhl3Z+67o1gp/fyh+ZESa3lr9pJgnW+
qYSxI34yNKRWCcEc7BwQ13jPA1Wc4dYM7xRsKmLi8iotgH+bubGk4eBfyke4VvCNpPkItJA4oc7K
I+b1Xp5siLISzASgUH0U0PxLAMdnLIEk2rfLpbPdBTZevryW4GIDPWhYdVud/PuT15VrP61rWk9a
DpBX0rry0VLYF+ib8V5GWB9dxxNwlguupCOtkTJKU7sZg99rUodLdGKVGYebUzyh0pWiOIgP7T05
gxUfEHPpNhDaiw8h5J9TrcXL7Hg8bfwW2fmKFpFeAuXc/SKq6OaEk+RMByLIvFXmFI2cXO9EnfeK
hsc+adJt/bHCpLIqh0xuW89jtVtpwJeej+6qPceT2P3T/E/EkpRTQGxbeEy0rFSDyyeDeVXqhWwr
KcTPSJvTggTSY87qb0UtVlykNs/Kt0eTyFl6x56gHGqBHqAZPW3DKAmyNM0TCwHdVgY1QbTvNjEb
HjDbz22+7YdGrVU72n+Z2Q1W1727f+IX4jRq1/082hxyh/jUnORxSDUTHbW0KpYDbPCTFbDIids6
gS1CeQ5/Fk2qGuwdWpGBh/c4TgBMaTCuShztSQwoN3OW7KsN7gGlr/O80BqiaONNF15lGOdyHyrJ
Md3c/q9hCuFdn8r5ttdNhVgY8cjkQqV6k7LGowdH1CHORFFVEgfvuCy1ig6WdQiwUG0O8tarNQAG
0ObKmeSx3Imv95ls2uqg7RyoW3FZdmB0NRVuuUEYWDiLKvoAimXDr3ZKOzq9OpohAIJJTXuQv/0c
3ppr6xxabEK70R0f9nw43sCMb2+jPGZ1fGejbEoNFTJcbVoYoKRNdjOsw4QnoK0z2X1+9GX1mhGt
UcHM5de84OyRJ5AfLUhmMvgqHo8cDwFfzvPj/HZtZH9TIIArC34eprV5duwTs1nsQeHwWFT40Bih
2Gg9EjwKwu68XyyCWaK/3nTh1o+W2kEYFrTpGEsRJNtwsikDaHO90K2ii0BuPYCTzEa/ZKR5vGEL
IFfY/pr6M1w9jSUx8YOIqwRcUuddAsx7qFZNfgE5rL4pNd/wM6vJ++O6ZXVuIQDbghquOrKsUTK/
9Y4VTZeWICh6BIFFEYMrNBjDoe5Gpr3sWgS44yY4wQdSldtwBt6sbcU0QGcpjufJ/qTl8aCgqeH4
MyBmAgJ82lYkjLr+fE8WoWtoB50cJA0MXHvV066E5bGHiGT8WGBOCaweTPiKjEJLYGIAtBTFiYhU
Ep5wq8xuXeM9nmOjwrfwQIl1G0z4F/sgOF/9nMJucEn4fC5gzormE1zMQgkj1O13MeBBUhNgwFm3
/W5Euzefqqwjr15pWtuANgUvHdmMyns16V0mAj/TJOridHSRwprAQ0xlvMSNZQTlMeqXDXfJVTqK
kG3atdq2RcUbcFPqeY8EZ+mQXl4gv/I1szUTJTwTAKZ8KOcXkt5wAAM5eEPW2lM8RM9acJNL+ps8
qoJrW/PbjO+ciF0w1rO0fuzIkW+J8esQrSiz0xxDHzc5vh/wcSnq1MLwPTrTpj/8JPD6tvNzwE4i
uxOyu9yCbetezNfB3XljCZaIQIroGQUONxdHznFYYl0MRM/618nB/uHzbr+dBB0MbUgBgfPbfg03
V2pDJaJ4b7pdngXcxXaHUX2mEeOKcIyIPiKK+Nhryxkm/e0gbHZsJApZWyYYyq5BukWLxZiM728W
s0faI8i7G+4LjAL9/g3RgC7w/zHZheRGQlGrccAwuP8NLPThSydMzV5ve0JYmule4wR0ocGUM83k
FfubyVqltTWcdnvL1d4CGyFcEsebIgu8jfmNdJztP/iG5kgE+kWEbZjSKNPuLGnnMONn5hZjmXjY
MoLloMQb6K+Fh0wvs0KqSmEpfP+/pyMBV6Cmi6suzx3MsYBYZ32P5sLHjw5fstnb3HMZt3E3+TIK
Ft9EHQdt/AJ70SBzovfeFBrdH/Ht+sa273/iI5xbbRFgkkHEK3zi/HRY7ZeLpRwG/o7sZj1N/awb
QgC9/HFYRmLFpXVkafvGwlnnyrkrJ2GJDeEChUmwt2BSvjD69gYtxnFrRlNfPelNnsA4403Q+me0
rGRYusXrNDRbEbf7EAQH45CDnzPTJOm5DmDWD++0ZSqd5l31BV748zlwowyHUYq7sz09bcnK7hpn
SNsHVEtbpIJMXzXivXp6WWUSMDt/RcpHSelBkzcgBKJLqyAJcE9w1w308fQMq9ptTV6fhlmGPYGi
aVJaOwQmcTXHmjYFHNJQuDuaN4YZ5Yrq2+9P2Tacq0B3ASChipO82nN6aUdz3xN6qlStbwypc62a
ts4ulmW6eKe3kF6M5SXBZ5KamffoUg3L54rRDsblBUSo0cv6PolQ/1s03/GP8qmTP5sVv8uYCarP
yFKzVbI6Qq4ApMEA5RoA7vDOmrUcXNrekFwsVQZTj0jx7Y4t+aWvvGO3fR7an/Z95ef1F9bcVh/L
sld9e5fjdf7FoJdteVYQ6CWy5qg5Y5+QXrdpAowUl+6XM4LIW1FyhU9BqS6l5bE4+EITs51apWQh
Shyi2UjNvvK9adAikZ1ed8UDdARIJFR9SqN98yJauOxSArqrzYgyOEQd2y13tRTmBYrqZnnJr0qe
UQ8rl2jXoF5l39LsBzRBjLDcG5tUlqgVlsQsYu5syYFX+Wq9mPI8xMGxB5CLKq4r42MVK07ApdJe
dEcPJ3Lbb7X5eyFi375+lySf6sU5rOQPLsH1r53JVCKNoyA6xUbbmdpOwAOpnINxpffS8ylZbZx2
pdHhZWhQBTlpDLxMieOiMxRx9GwNXiXiDM0wJjRN8EcfubkJ8U9j/oNGAzmNxXxgPcXuk3+pnGHI
4BiFm4GZMHGWd/Vq7C+nkI1iUUjaYvvoA86QyRjQkVmi9FIbF1i1j+qRTrtxOP6K/mfqvJawXOsk
249UNm9ZOzFtFX6XogcuHTGgHeC6v0zmH0DLw3RWUBwPUoBZMbxmmA5p8260twN9nk0obexGngv/
6C91nlxpHNJyT4RsYlXoFbXmWeX1SX3XwNjjqtf4EQBzR4yu8obF9jEeZqzqGoC5MI0P/T2fUxQx
4nDrkkUGasddd8bgxOqZ0Ar8Dh9ST0dfIa/KXsRq7I3Q5G1KYboCTpa9c0GW90XIiPG5JVaY2xrL
PeqJfScorb/Ji8X6gNHdMqx/UnqMhnexkqT0kDY4bvUDHUAU4wRQFpmp6fnVYmB+Navbb1AD7+yb
A+EcmmHeSTzUcUCD130IK6wg+ib6KQTLZRgve1Vnr+r9gNUWp97E9T2luRBHoaF66NSXOp+rPUX+
GjGNhrTm+DpZenBjFq+eNRfAQDPT+Z5E7liIIKI4zr+w83GU6wuOqlDWxtLT+ZsWPhBEN8d6bLG5
b5aO8SvA1SHcO9ShWQODXiGBqWCivFxQ6cnlVsx5Hfyl2LXBadGNpAORxW/B1AKPC9IqMoYZhjNr
fz/bX6TgiWG/uEs5idoB9nio2ucaVpOmQuuN4uuL6PAH4D74fIfpA8IM7ZW6QhtOr3qQdSZL3mwS
MHSxtXNbBDeUaWZ+Djx1Zvh5vo2aOuFA4n+UePC6UUn0T9LPGl5mu/MqHqMYi9yfPTLfe91Is/Kp
TrkKgJ3oHWWCn6ubCb+WXRwYKqP1sKexRGtrQQHUJ+HA+/KDo2iEz0PuhkYlL9CFy/b889Taw/He
wtBc7j3pQkmcXjprQM7TSS3MinzXqR9N5nkMp6vAX2ERBzhm2w66qa5qyeCc0XhsDzMeH4kWwQS6
9+WGrQXPynRDzGQxwVNijamlWAJ1B2dRsOVmc5iXhM0OWFoLcL2Q7TmAAHUD4en/COVK2NgCuZ35
n0QZOVfaWqRYN66xVf3HBMrOdMcT0nvD+8HNWIDnJ7v1iRrsqm+gWGxkbaEjqIiEwFF//YdIkwIR
i53Qy3xHaNUMaCJJPXoZvo2p3Vj8zxe0SSgmV8r0fnNkYF0f4bFsPov4JMtj2RjY3/kZ9iJ7xsDW
s+H3Y+4BC89z+W7I7rk5YIe0FI8vugaG9Ys+6jF2GvVkdEVvBskdQDQsRFLAp+cr1hALCSC61Lei
Y3P1cZPyHFGi4ZC3CttJ54pe4f4vmqlObRJbC6JhPLgTtRMJGE0+9oDRL1QDeUHuKlDjpddmk2Ii
uEu0BpmKvnk1JGYp00uUoNGVNCU3nU6tHfYm/h8ncr+LcwP3F9IQM3a0SXHlJMUn+MQfPKB7QQ+x
u8bqEZTbji4vJ8qCcjHGcQZkvUVgoTjQoqAF8skb4LU7UZ02H0nMw91lou9l6vuCZ2i/cfywN9rz
AgS4DPffK4e4Fc4+bktpwDJKClOLCYgSQYsQYRYHq8P2QabSd9KwI/tycVy99vIgPc5tgAhM1y8z
jYfZaJChJvNEeBvIi0n6zvhBWRK7YaJQiAscVEEqRTcK4gQ1hzfJa8BDGecnHqGiVC59G6CDRVPv
2Tz3ANpHwKyHIE0DPiYQzql0vIkxP0clHUuaj/V0MmxrLbCJEV9aH7nsfyR1Eit7DYPRTzhB7rnE
iGkc6Bt+aUp8F+pavvs9wRri5q0qIhimzosBc1HQIqD8OItWc/DdaDNQqPtVDjI4yw3F670Jk5zx
uSr0PfCgJ9Kn6rlB15x+7h10srp+2MMDyZgdoYqu9+7BL4Bk3hsLbr7VqWs4rJ5KR0zeIvEJHdN6
6tSp2E2Tzbhp1HaI1JkeWrLe44Dod07kX+koSWsqtSAzCXYwenXnglCB/dZwgYZJf0mghYuPx7xM
7ouPzyf/QnUahVSrpsV7V4Q3WDRkyH24mtQYoiGPvS4w465CL4TcPj5fpD0rbGS92YKIuvB1a9gm
id2L8OCsj88GpnMKZJuyGKMLyFQGQPDDXp0OYIQLSOQ/30I5T067PBpfq0/mfHZzet2xeTeytpOX
jR1elzO/FbpKWidMYQgNK5NiB9yG5RRXGfBZEjfR3g1U+wicNhUPhOGX6wJEjOZenOtEugxIMhAj
3W2KZrKF9tSV+ok2AVg9DZBk81+rwENCvRvbEzNCN7oDlXKFD3+VG+WBQYTGNJ0uQdlqkgs9GS5l
ZLRa5wy5bLbXDJzJDEegvsC3u+uS3wJrjV5pAN/yeaEwCJBtn48xshh/fBal0YlDlB9ZO2cElixO
v/nea4ND35J8fTJWIDMBIWhIighMHMHfMsD0mBH1YENhrtlHCioQuyJAEkERBumZIhalmLdGOfxq
4CPAX9lJDRpdnTq/78A4B3AVlaDJ6iJOMaa5n/bU8X6julb6sfWSyggI7UG0JChgiMAI64qCaF9d
uPDrvVOskVd4NC4AfyiA07h7cQ5vfhUUidJV1uigYjiojBLP0yMk6lE7LXl1MPvElhEsc9qP1AHO
BdGlknRbyK2Qr6BlbNTaBjRM6Ql3vtwTpRWjPB0Quy8R5yGybaGEmYYod23cZdf21C3UDv7WYSqo
zdln2W1JsRv+uYUzCVbE3ToFChbXC6Kah2s/d5DwpCK+GubLoCOtJ8JYYgvuqlT2gwdlnCQ1xUQF
FB2E6D69i2b++hvyN9FgxhlvWxUfsPDKZ/tXCnVbesD4y8NzyMEMDTVF8qePqsShJV1RN0WSSbRp
D/4rbW9yzm8W5z+Tmqkv83ysdMeXbWUr5U1xZkKSyd8KIMj64ZCrAG8oWGmH5juh2w3wYYHnulnM
2kwPnX7/+G63jgDoXRgHTqrZFp9rY7nJt9AyeFJg3Y6pQPIYz0sTYGKbJlLsR0tVt4wSwXAIAl+7
XmIKjrZUZCAyV7ggAwwgakLKyA2yBbIWy/tBxFUtMo6G7e2rmfQm8GZTPTUVnov755OD5OEnH1M8
VwN7SmVNQdx+8gW9jZlOMwUZNrbdi1jtI4zBGr7RLCZSl2xXT6eEoLvxnhJKCx0LuEVVB+ytm3op
1nwKnzBjwHvCspA1yf55MHQgGLA/wZHYWQNZP83arl3ccH2N2g0KRyhmByDyrHiHzxItP0CKhz1v
DE1iJguRBXWq9m2RJO2IPnbFytFjObeSYRICh0n89RLaIO3oVSR9aeDlEbO1n8UbpBuHtxxZiJUh
n/KKJLI9juWjTpmP/F2Ha4Oj8LbyrN8YtoequN51Rw9bGlLfso5t+2uiZo4xCnXzJvIjBdS6fv91
wVpmtWZzxEslNPMeAM3q2C3X0ioeMTE0JOnBaltv7sO/wVU1f+bRf8RgnzMzFySPGimGZJJaqQlh
vQhCV3BUubyioAzIttUi8KJGL0yKeghg3/wBV87bjpbZqRuia/9d9ZjS4YPRSlcAOSv+0t0w/Ohl
hEl34WrU4wH4k1OS7ET0BbjmeejWRfSmSMbZ9N2Glf9ZBKLwUoJNrpD0g3WGmQB6mcCcJJxyrVTi
DP5ata1urgWrNPJIeCAfXvlPnCtYVFj4Pvp/KRkAwOpA/rgy9j3MsCu67M+7t6Bn9Xhic/Z32lJ5
X+l6j5ekmpXDagfbKZ9N0cbWfu7reYS5+au2s3NeeA4Ch8HRgZ05V8zDEjsTLddiT6Q3OEr554q2
Wc2vi8EQccvNLqW5AIMTwN0SIcIYwzPgc8K3XYKze1uTFXraJVoklNEwvF/nxjTD9yKVAgR3uHJJ
9vebs7VwygSyAFMKQ/scomQywI8m2HWCbxtsFU3l0eFv/YN9eAG74naBqBGa0qnttQ20fvZgTASB
WFOfysNnjdN716O7/Jfo0yosX/l81FV03hij21hZ9sl8Sq1ywoav5ukgunnRkX84La1dX7iv2NUn
VlKS+oNTxBu7hEaeTtgOaUeeGFKLhL6uqdGyKk/j19oP8JuhCeTVc2spDyNbJCX/Abx8lk1/+TjK
Oejt2/MF4aVK5mgZ9m+sCDfcatPZTVAKJJV/jg0HJM340dpFaej5qX3qIgOHrMBGOKxeO7wkrKwI
pLMDb7u7SLPC2T+BwbuNfyqKINmSxCdd0D5ERuOqJM+t/mc+076guKMagQnuohiYCCiG/1b17Y7V
fO9KnXNkzb45U0nBFPUU/1fqwYMjxGHySEb0Vsd+pX6TUvfl2QUSlkGzT7TZ7aIIrKpJpFMyzCuj
1tVu4XbFNmAzn4ynC5hN2tujM17T56vvh24jynBMxLOk2PjoijBizFxiEwrCN0k93QY9teAwdPel
/xBCPCC3phzzFwkUwxMjwoas1dT3JGKd1VDFPd2bh+PGC+bX2pi8pIb/QZvUE2m3r7viq8Tmvvc0
IjXRX3Rf65z0q6yisnd5oAhAV5cOslYnTA1TtI4AC24Hn3CGzAMq6ejdbX/e9JaSlhTZqgnWUjxB
mMVVBDkNX17mjr5KO0WGp2qWGvgh1wsJ4sThnJ+1HDGhOI660ghvDaaB66uy/m4eSvgNk3lNe8/2
/1uXobPgV/yiA9QNjDvxhpQ0wnLWvHWkgU+xpCm+okjg88xo4Hjzh6qfjnPKF53ru+LXpZmlRfly
MTtm/pJTU1nEoRF7ionbV0SJhyPZRD74HbBAZCuknBcrUN+7N96uBttNtFCXSdAq8uvzU264pP1P
xHGCkpbW2uu6oBEit3vZBxvP1cgQFFfcHPMBzehrhm0NzQv8pNjnaUYhq/cZQUNIF2gQKWHeDm1j
nT1ajyXs3eV++bitF0FisWhU7y5kQdLFek9kqCz1NZvMKSYjVZWyO/WbOB/mJj/QbPvySDlkYsh0
ZX9Kb/aqvOMlH7bzWRw7XhMwVQceN8qXhvJ/e+TFRCZEs/vEa/kGOtiQCs32CInK7ouZsTCQaSnH
I4ilrcoP3DbgtjtWIJOp5JatGz0l/BSGSNbZfVEjRNkn2noVwedDw2yW75Mts/nGnBQSSnWwKORX
SuuJTXMbcAFVmsEuJ0ahDBbI2svJSBZ1JgG8uFBQubA6dvrvo2K/hyUXX0yUNQl1Hlm2MbLJCSRc
Mqiq4dyMgydAocqdpk6dKegAtlLKEhTe9+jc78/EU01vt7/nNP/j0juu7A+7zycj9RKN8davl3QS
bgMKFRdgBK2XJoNqU5PanT0+kEFkXUxdT531aR0XQzY7u67rNhawsJSitKhoig76hr5lLlmYsD1W
ln0VXFEmf3AzmxPVzI2JfT7uErD5oj7JsgcC9c+oYZRd9qi6s9bL0zb1QQCwNSjZakwddiz/zNKx
ziOLZ+SVlJm6PIO+VDsY0Fd1O/g+hvpMo83M1kajtJnjwUNtMt1iomXzHpHykJUjBB6/a/YbSJNG
14xiOZLUAz1SNqlJV0mcEwZCiYUwZIjHF+ye5Ug30vp+VGHX8bsjN5euzLmu2t2Z8mJl7OYiL7+q
FMuxM7nhMB8rUOeCBPyrExG86UCgJ+dBS6zP6Z+rse39+rsFJmh4Na2I7bjYjTQ+77IiEuDfbWNb
gBZj2IGUTzR+A93n1rd1fWTUUuDuNKsiN6DQqysV/xRqIraqUbi0OUi3RxUvUSStlhJVNPnIS5Ze
ZuQ0UBrN0nFe6XlnFWa3FPQ0zfKWR+NEGHX/kVCir7Yml6XStu2Zc3OM+4EzGoKLacbTkkvry41a
4pzhHJiwY2AkuBzcIALVNYL4478nh7j0Pk8/OAhn7cZS30cFt7jzABgu8+t3HYr0VZLRx+Atf42l
1HIhvEtdJMHZAaR7S9rqkBGjd/5XrgTfB+PKArHAk+fSrrw3QGWfbX+Ckz8mBZ4BwASR2hou8x2Y
aK9mZwpfrhcxgEj/vl6Asz7LwX2q2UCTOMD+tq+IMxjrzU9kkaLjiQnhHb8ltidjKNBBsRCRnoAS
tVxHsDvrOAUWK7yNmVjpNHC958afiqqJVE2pbZRkgUXeVted0dM2iKefxpr3z94g2I+6VxMX/xCC
BIZpgAJUoaQxD664uzNFmiEKi+JOu2cPWI/diJpa1oIQ5xh4RTjsOtIj1ccLrT5ndtQyfgKHJbMq
157rz9UuJYjMEa2oQgis03CUl+8qoq+ZG4XDYn2FWZoTC8vFzXyN9jjTKqILqJqgsS/xP4jO+jeP
ZO5ltm4KwQuBJ9Lkq4RUbCiSRdRw+g5UwrdFpoRp0pbssRGiI4x1KMvZB1+T8zIPgxBGXnmTZ+cB
+YYp+MfHx61gHxm3f+TB3zkK4042eamG2RCgptruRQ36HwGf5gLCHBxskFjFjbRfkGDdvlXqHSSD
5MA7du1aUlVYJ+GKhKA0fdeSXzX/AlmZVTW3w8LdAUVHWrpfxcmip0f++rBHlpXJj5L5SvYIYnPk
z3gdyBnsHHsYZ3OO7iB3nmEl43037VjcfKJZn8/MMLqrqOaKFbMSu8utYlgSqcz4E8O57rLg9Kj4
d5itDA1z1r2UsgTdxUe4R68G7wQ1WuOpOfnP0ZapQOtPWF4YZTcVJwLwZWX54V8+z4lxwrZcElnW
FBBS0Z+YwpTCQKY10QeFthwMNC+WlwWB+C0G4EH+auALfwhCuJU3ZcwB5OGfc/+Rw6ck3IHvxMul
BREWvS9j8TtJHByudEP+oE5Iu4TDkLwtpfczoyxhHoJj1Ug54zNOoXqHd4LBpdOZnpy5DeSZbG1y
1B15B/FyaNVk6hZV6Sgk4n8bmTQHYeMiRXRdvTbCRAejVnkDnZqDhbuvKZnUAF/RQ/DoLrCxFdQ9
hH0Xe/fQZxygSybah/KfL8jC9HewDgQcU8qkPaR+fdCMl+sqCVHrhTxfnSgrjbS64nvfPOosMkOV
xMPZ9mZWm37QPy0bH11J5Og9hFek0kC3kLIdbCrqVXv5yzyGjWp6JAbnPtyPPxhykI/RSnHwVmmm
ihCA+rTqPV4C//fl0BWqU039EhV/MxKqDqzogBrhoHZ70jAqm1my6RpJSefsyFkN7LarDDlekw0b
CARldq8vhqUWgtRWb540WREItpeFySxN+wjGVG8HieCFTeyCjbPtgnvNVFD1valCvxEe/DdMaJOf
LJ7beIxNlYu2sQebm1fEzg4ECIOWPpmU8kHNwKTimJ9lb37UXq/Ol+RLNalgEqfH1R6VkBBPINtq
VSM0V55fYdA0cZvsbJ3E8xlLjN/6yWBi8MqmSQYNtFBdfEtj48iDTZcQC+8TcQQNmjNu4VL2MHx6
qlLAS0K/wzpgTUT1orYpdvnwChrhUKZlVez9xVaWzHOzvyQfdJQ03I4aPzKfq3nC+hgN5pIkf2r0
tWqDJGAMlhgL03bj3XUPmGt/H0k5PeOYnWa8RXh+qyf5gIbE/6trGa4zoQ4k+ilEhVnE2w7D0kC9
FHs0rCI0+qPNLT/WXbsVcKTjLiT5UYyF7ZFvf9jkaMpANmPidoc7Cy546f8jCEyXTUt0MldWVLnQ
mqc/737J1BCPRiUIw/j4GnRqXJASxxWsB7uuR+VJtAEiztuW8lYZN4TKQv1571lp98rsggjwIoZ4
7X7FZKdDtbFpOrykTJtiE7qR8aTVBS3SkpR+aHB60JDISpWWRb7KmXeZEg+IbJpBPTOt3Shst3AY
vcE3JxC7KqRvJpnJmzJ/lvmHEJtyEd4r7R81fCwGYnM8lSKvc5RjW9bUBj38Ppsrd5wW8oMnqAaD
h2dLLbcPI5prf59z1bpBaEhcNOuOdtprQuisDje4hOiTbnAQCl+ztWyGJY+Z3sxVNaBwyagIB03n
Qze9UFcQoPFjE8bbt66O4aqJX/JRFFusJONguasM9tiUjGW29VcDIQC7fznsrXBd5Zuqdy0qNfkN
P1X7/olAShqKgkNoZyo/H9ltxlpX8DniufMyNfujiLj+OeE3OLygQHz3wQZPpv2LOVQJI8h4qFqv
If2pBstYwhzrvEEDjKzegIW6L6yMbfgEIhFJflg/ZsINB/1l4J0PkgpGqVtcAuACFtQFW8YpO76w
aGC3ZCE4fMEyyG6S4Z/0rdDUwS5hSYTi2glAyoi1EVX/lsEoek4uajynKZn2bDZGFa6XoDoRE7V3
4H1gzpl+V5d2SJKvG0wgggIVsb/AJdDvQk0DUFOUiG3L09qp7tsJe2X5C5iNYdeIHlPHnHeURjib
jhR67OZfqsoGkF2NmbTtsB7MeYOXaZqzpgXV9COEwBKWASDOoKP3U1CowYVIW7Mg9bAqRF9twEHo
wudoDjcZFUG/273Lee2zUYMHhvdr4AgvPxVD97Yz95M742zjatoRmxJRkZpVNSuWMQ2DQDqDTU7X
xUoVYAE6MXQQHaTseT6XpSb/C4BL1OiB7LCL0Fg6eND8snQJ0sVmv09CBdK3TYOFux01oq2AvWlZ
FybxgX+71GPNvzJ2UOh2jjK1G4Z2FYeeQWvZBOScd1eLst52Q/g0HsfKmg6kYYTztb0vuXVcZLDy
THPSkBj+uhja3iT8HNYNG5wMC8RbsaNb2T9pPP/0dShgbg9rqBGqnJGgz+d4Uwyx3lQ+f59mRokn
RPX+2+FUkowaEa7rYBe/xv3kk/DBCQuxXwKhpGntJEL1LEPGDYa3OUIutizeQBNDOmubOxoJCT9l
DQ2mob8M4VBRLlYAYuAiew3EXzBINuNXSMVa0iU0CYJgmohy5Oiy2lgI6TFZ9iJsqAwKT8QtCU1N
Vn0pknZi7oaQBEpKQfTrfhEn4DawkxNyBruWisnOvfezzMXZtX8nUAVPMbwg9YKOPLkKCs0NDPcy
5yT8StOkqV8ETdaZOSXXjlRBqW0q1alzpKrQytWtOwR2rGKZSMtnwRmICeTStWiVMTkrJdIYwxVV
vVgKh110s25a0LGeOvlJiWnubK7HYpBYpLN0feXUICNHCq6dh+D2SNlrEho9UjwYtwAiTIYU+v/m
5A/OGD9iQQKt1CZSr00TXSAGJlr1VkvfkESZUPavqt7VncUFF1Moal5YsRRITKm5ph0Ge2tdRE6N
gouczczpS92Tvc2yNRGl5n4lDO9NV6z05syAxI2gWBwaO8LgIjyE5nbv9LS4fLbHpBwTc0bOA644
y4C6oZ7ystuzkgylVjZIEJ2Nwra69S7vxO52EjXWV/Zy7FYZEHmj6e3uTDTjdRajVeqw1cBw1BOw
6lh6Lc5vZYv0r7X7cFyUhoyUV3pkn4NTDfuSZWzathHd3BoXKT+3pLYO38Za6hmN1Rhm7YHyjsVy
yKjIEjEdcjBCEH094RUTSK0oaIdR1mUv1Waq+vi+HwJ95L47YvwfDZYS+LWOwYaBM/+4Abm23BZK
umcvNVoOJPwxT2f1xUsC2K7W8JnHPuQvKvfiG9C5kjIqZOwzp0Wr3D8MkU68J2lnwqbPbpKNzXBn
X9I3gwA6/3m31V8X0TAfmqkOpaiQr4hgTZ+GZc5MVL6eO3tsMYezjlG3j8RgpVcpcbycg8F+GFwQ
j6ElZpMEHS9BCUmMuPpNLOFlRHM/2gsbjENO4LjqAab9KpFyi38MuZM32D+/AdiVHpIQmww7vy3N
S67feDLaUVDeb/r/TzSnB2EmyvTh4qa358BZKVd3UhDboY1paWT2/3wj4snJoQoYeWxopYlFRopc
R1IwdcUVC5KHFRTjLTURt5FeUQBC4nyh/p/D1/3PMwf4YIKfow9NuRRbuusjyjWF2VmF6in3w8em
n9tpFiW9lI5nd7msZReFO7EPMo+L/i3XsMB2V/6PTD5IADIjXTz3r0/E0HHFHCR5anoD1/pvDHRG
txo2bMWqanVKV+WSFXA8N1LyjOzTQJ/03Y20uEP+4/tKnhz/WTq6wQ6dCvhOo18bllYUvh80vIZ0
JPC2kbXSOnxZT60tNC1DEK+VDiqU0ViQfIN0JGfINj660T8C8L8YoetbNqCFXm0cNXVqMjY3pZNL
thKrIo1kN3Xki7buonwDURj51LNy7EQiti63FK1ZY5OzOxU0DEqA/Qg/PKR//P6uLQjfmjrHK5Qf
Hc2UXpDvBecAyzkqk3BmLc801e/tYXMcazUFZy9tNXmmGgmWkw2grbIPhk+RK+SXCn4m/wwuzuNj
wfkIzulo3XnFU4BX/no+EwnMmwPkxhhNk+RO0YFgskoZ7f9powl6+H4r10l2nRpsOJbvnh+c52zP
mK/HR1qoKxmmBDe75aFDCaWdHcFXusjMBnYfX0KJ4UPK+awdSRNHx3GBJQzLTDtpKztyYphv24Ua
+/9fyQaOsL0zvxJbqZP/VdZ6v2CTxafzY0Weedwd0Rj6IKtD8+9afXuDYUbFtBsDLb9OzfGkJfDT
0WYTXAushPM5OCkMjuN82OlnkHPRDPg1HO/KbwbAfH08I12klVDwS6ooYiKHciEq6MrCnJxr2bnn
0v7SmMB/U8msMY7onZvW+v80Q/xzG8DLfkSa7IAgkcfj19IjNEbb/PzqNBXlt3tsZV/zz1yJdbKb
yVjyTYcSwZBeWKMUothUCgjBB0eIl5KwAECAAya73FLimjSwhF/3iipWK6cJIuxSxvh2Q1j8MfJE
43hh2IkpfwIWgf1awMzoMDYAG5c4d2iycv3mhQ8V6bDligAInjIjB4dKicnstDuH5c2QJ1KfNkRj
q2gpWKIV0Mur2rZhoedPRlAMms6aWTX7IHrUT8d16KNiaraeZkWb7olsutzYzSuq2/Zbt3XKb/Zl
A7vH8Ec77q1BfXWNI0b5Q+AVAGveP1AuR6DPTSWH14pWtf2S+TR+sgoqaTCtMSAWUKNYutaL49qK
N+T8hmo+a1JvxXjHywmiw/62JrHpf9KsXcfYBISyc4dbKRH5By7ePui52TOkmYIFDCD5pfZys+Om
lnCoENxeNxkLycj1Nvwmq3a2NxfN9Wab0uNmh43UTUD2HrTKo4blXDd4nf8P/AdxVu1ySY75wocF
lfnQAdYRoi7CDa71OLmYBybyUgjQiRyiQbFlkr3clpSad7Hte7zcIZtMcs4/xYmm7pU5JVl/ecRT
arkwCqh/snbxqY8ogHM7sHwOcYOPWtHdMg+UbYuqqKSQUZrkjFOwh54e+GNJBvV/m8BLssm1/7EK
zNizVUyN1Z6CoD5mLcphUeVrZK8OTGrJFdAWjIa/wQvNAeyO/q8K+2MixxLvYB9Ee1pF/ktj4C1j
7fGtPWp/k95QnHTGW1mQsA+4AVCxwhgRbMEs1vMKvdZzxSYcCzXhUDbFOHgSieQGK1q65syWD7mJ
4juaGmXH2ArSDbdXscQepoKgNZBJPqA0ZLqd1D121JErJfnkLQ6I3v52vTnd++uWhqs4cQqY6WZm
hZfup0pYFKhRuW56YF5BjtXFinuJiAi0dKeV3c62JiXt18t4ERFrwexJKAailC8gnF0FF13OV/DM
bt/k3Exlfw36xBhxxQhHvjvivRCx5q8RTQUz6WkQp9WMqQGoy3kk/2VQxR/t/G9B5jYoZCVa5u1w
cPvRhwxoiqGkkRrWOuwTmczkdDy29fM5KwKm0xSvzCf0plZFXjayDt3qeRxzRXlv5nPksmBkg57u
s1OVzPhrI3ruuXLVbR8JfdIueB2lS8Rx7wL6Ro6ziEUuikHgOfjBXOjx1me3IDab0fPG3SwquJ4J
cg8JnPG8GLpnBVvcbuVe5JSorZa815DtFh8SFyJ2qltxnGIu40ZKFWmr/H391jsih2cqNv+x7UDC
fuEMwlZRIVDB1xdFyOdxtzEWGuTy/gAuzWEw1DRmBvmznXdngm3JiWQEjOwOkaKa9Ie/MfmjR9uK
cAK+qGhQRTZ6HzgVgjY88gGTZtErGha7ojI31n4A97aLSNwzYZdtHOb89PQttCOA4LN5r8sfQiTd
746cTwY4qP2k1rMmo9Oqxs0qX4OSTYvbbytliqIvUMkzFuIpjJXt1baoR7bVv7P7hJ4Zb55nfr3t
guRBbs3TajrtIffj6sm/1q8vDeenT40if8beMVNNw0399RWSm7k6WqdIwn/4oJOUlpPXqOTDYCAb
B9jNVnDQS1HpjYQtcgEPer4OIG/NSDwP/t3x3aSGg8qpSba6hpbvAfqKVKSjDasdw/IXH3/JYOMk
Kx84AN9Gf4epW8xYcy5wwmxBWyvalOBGNI1HRy85lL8VvujjqxYkpydWCxl53k/EVSDi+d/3mwk0
t5J9ozH1sKVyVITFiD6kCxuIKQ5iD1Q8r/sBnnNSVihtWyi9fnK3rRC9zkdHSEJ5mXtj9MhK+CDv
LcC0Ij3UhIqOphZF7Ik/WES/7Okzh6zeajM3Yrz8pqWL0Kq0PPuEo+c3QJD5g0LHsqTBrmMODdAf
751rcQHuoXKuRbVwrs9as8qa8YjBW1+P8IxTZ14nIgB2I96b6+9y3z/gDmkcmiJtE9FURFIKBXjp
GnYP5ruDwETYVZEO6MxnDW8/Q2BrbEy5YILd4UXfFE3UBHG5uDx3FhGSssflYwiYD0kFULYVBR6k
cZNTUhROxW2nga1AVLyJ4YMELqLTtZI5jwDocu/TOXSyfz11VZIh/LcsOecP6Q/NFRSNy3MupSTt
rUEK4c+Nh1vF/OuXwD/6Cp9F7fbpCeJ8alJCuKFSEi99TdysTLXKPylbQgaKScVAOyn15ktucOOw
kqP462LL5XpziOLmlhP43CeQOlPSwn4zTMw6ZtKqqQy9QNOpUkC3e5UlwhJbhra5RxCLiIn6FKIO
xP8Art5Jc/FhbPx11S6CPp5Eq/SPkar2GOvAkHETVCWjpOUZFtWs/AAnmcaXBze0nxBooVR3yWtZ
if2No1RspWWNiK7fCCkrM2/3auirSPirk2pDS/176Kd2BEI2K2IF1cNUBBRw8x2NS6dAW8FKqAbY
0HkxIXiSs8E3+AKC/pHoYEjrcfknV/48Q4EqIaDIvD/qqAiR9ifCRlhLMj13Qj6VgsHgjKG4ip/G
Uv/ijKSwRX1W3hRGyibwjVXMbk35HmqeMRnHJ+FOylb2lgdgGmoT2hXfpxDxQvO+caBROAlc21UG
xqA6XYXE0mGrZJgvhVcVHcgEo/K748FXxgdPMcn2XPbVfCPc1QC8ERjJTtco9BxGUzH//RB3bWgO
ArwI1/sX516euyHRFGvUW3wsnGcNErs4ggS4/sPFT7cxkF97OPnfjfs4EPt4TYHZqEGuts9zu3r0
n9rJcW901DaZjuJVg9sRuKCtyif3BRgr/BeHfwAG5PCzP8qFXz2Y9WnHtwU1U+Dfnns3/bbsMuu+
QAUpyU5BlTVO67jQiF89dwEg6eoX84m5IENgdi1vFf5XyStFKPzNLOcHs6bAMG5s6bqCrWzyKbPb
Hc2gYVGgWfLQ5M1M5VOeeTWgTT/ZTOM/jo0bl96X2UuS9dKv2cmbb/SluYH7n1hnVWZlh3ncg1+5
bf9dmPt6eyjjQLckTbSRS30LN2p54gWE89x8dhUReUQk4NU2rCL/264RuJWALkJELFmykPY2uvGH
Jzx+QdXrZUZ0AeDuyCuaZHQHUtBPjEBNBuIKg9p9QsME4nL3sFg5RwdFDLybv4Fs5T3X9dLwmPyJ
UfOPbxaNXui891PrgHY//O/BRklX8+B/qARNjlRCySmYGelurpmrwjizEGOL7ypaRqRAwsXID54h
QJf9hM0qSrZSZzLjVDvPxJRgGxpw/0mpv5Sy+NMr/1j9HS8VICdtFJWWivj10gi4i7CgnV429g3B
MRR8vFvGRynR6wZ9Ar1bgfTiJ2AbfO3RdcQV55sdSaQ6rzTqVmxod0s0tUPNFOMoKNCSMepWoA0+
hz6xw5vKUJdXqTgNeF7YeGDadudsXhpQrq9DFAhXvVgpzIMO5ugMl1IVZI7iFTmPR0rguKF+0YIY
edtfuovZt5g3PiaB17Wh2/13p1Jdh2/Q4okL3x5laDEy4Z1PVTFqcX7Mxo06O/wPd6jXNbfvoYC/
jbXwMaVhjD7pLN1FRCE0XiICUDlIFAJuEujUlQk81reVwWJXwbJPK8bQsNQTQVWej30U1VITDZQe
vCO0ZfHUPvTqRY/QVoCTSQzAVYRh9TdyJ6kYcwKZt/9AWYx/0km1528PpOVN+sAtUmUyXXBJDNWW
HXlluL/gWWM1CvG75qpHJgSN88bn3bCAFv/E75nhSt6EzaDhTkxLzU41X/bwNnAuydA8SXlZJQ/v
zNhtCHm8xKBdk7Wu+uU3akhgWV9ous4a1kFE7IJdIl8mWpgdRmKc4yNXp4jsrqC8I4G53/usFOUt
N68bWKRHnhft6iWe9fXHlp9ODBZ1jh1VLL8T0CYK4aItxtfW5mfyrP9bLTXkMPoIzq4GoFCdG4z3
5BgP1yQ9fY4WUUt2+ZgdW5eHjbdE7Su3Dl+7pJ8QeEQDr3l9d2uCYn7tmeQQb4mOFYcn+v7d9jRc
tHJn8I+cUNR214mhoOI2ITQypY8w96QdJy4aP9ZVHE11Jfl7TsaI+jh/NmvflhTWVLQCoOe5tqRl
SYl7+1wlAcJ/tpk6EUNUsj/WytNCy8GgUexkQyg0ttFE9hdnpUlFhKZUtyfFZMPUUGWcO9j6tvB3
6CU9BfCwvWtIZltsuJu6I8/6RMWa8g8p5HvTMwjSoeMh/TqpMkTb4jhVCARnIhJmOvhx5vVH2KXW
eZK3UsTY5lkIdSUH8t1E3/ClOIXAKCZl6POTb7sMl5OXjxqA4R0clWy3O0q/bdhrWihup+bZfOfB
k+TGGygUWJFuSiGQKrYqtCn9IXo1Jj7iOip6zNK1VE2YtNqlPzXP881xwyqjxIAIHTeOwSa0ay4C
AXFl2nYwPVm9lf+gmP4LOBXAXvICkIKyx11wuYr6sWRZpnPNav9pkyEm8oQrqAyOscZBLYujoT5s
xKUFA2fGI+m7nUZruWqPSufFHMrMPfq7TLjkzmTZKfkJORQ0CvEw21M7SDI60PyIQOeX7Svvq7w5
6jxxV2c0zIcggaTltyVcBCcySx/MSEz85TPHvr5XTL0BzEcdcu6MbXeSoKOVvdSm134dsTPv7joF
H+lY3cDeSBziuGbeBi6sd74R0Q1vQDMs0A14DV+c9sWuj1FwXlk7z9MmnpH6OK0dZrNFZKZ5MP0X
pRTzrOef9gnN0NtMFGtTd9X7hzL+O0Jo/nQ970rrCbRu1DOhqbXPn2GcIY0DQzybN4/gxwib3B8x
Cb18wKqgO4x1y3+zY/LbP/FK66vKINiQqDmI6efVmiJz+IYRTZ4klylIpyQLL6DXrDLUtcxdkUob
5NrA2T6UGQufUhqJAfcn8uEvmIToFkO2i4ihESO7XBWL7sPg3vbDQBeSMdahUX0EN9P2PUOT/btZ
8veUx/hNuux7jGUx9ywkxanRBJZfm8qdeJkCtt3WzZ3e/91bI5QDdFqFDPQmB7Is6HokKq7h6qnv
MFqzVFRkcmtrQ5TqYDW47wr8+Ha69vs+Q3MPiWIp0C/HRJUYYabanr5hFGtHnIvI4zaZO1fZoY2j
jUVfmcnladVjs7MjLs9NL52I8kF999zi+wHiAM5CgeTNhklTjdKVfcKDx6acmDDxlouNw0LVPJgc
j2SsgEgRxFh8xdnpwjo4Qol0w/OnACYUUmo4/TvaOYiz78rpowhQ49E86vT0QK4wIR7CAQ18ZDu8
xjsbAXMnwkax//u5AgYOWPlHhND7dn1C1PfE4GycnVHl5QthcMDK4VR2PeU7cKfv03v+8x0CNQaB
ciLlUtrvSts5rcNz53nMqjiek5GVuuWjVg8efd27FkcA3dgzcVH0M7SJGHfphdF4V0cQWN3dzTM/
Sl9qdsmFmoCZALNKWemOrkBJqxw3aYOufM8ejxBNjuxR6/zB0liItE4xa+6jAaUd4WpHM98KfsPV
hfiaHdYzgRqEe6QuaNGUqLHC6a3c4eErDCdpAJJsWBp6/xh9jwUVSVaojILhzOYe3DuqPN9UefmR
3LfOAmfP2vlnOwI/Rax2KOovp9pyeFFzXiDRTFGvNsO/cLypV+/5GDdHOyW116sRZxpEL+jqAWlk
sRY7rANdZ5Sk3ia1mgAoJZR6M7BIqsgrwV/nSdnEAtFRT2rirKlvFokCBn11XFPhyUjKNdqmFvxt
nFlc/+96oXbUyEJ219Gm1Rk1fgbh4VpsbeYy72zA/6M8h/e/tn4CH+BQWu4BW7ptC6jgP/lScAdx
MwtOpsAXDagSH44BOUglqBpGADxLLBI0IvV6DmUj8MqUDB+rR6k+4Bf2wdYenQdjkaO4MAzR5xew
pVdaxxAcap1yyyKQvkyScrMSB8tFeJ9MM1wEe1XSw7MrTiTR6mImzhgGAec38vhUqE/uh3r/o/Vt
cASUH2qap2EQovO2qGUJayJzfebf6grc1UUYCwITfEagb18+FskS76dXVLDcDO4wccLsRYR2V8JD
2e3mAyBrN7EFo8WczAUaPMgdpi3hq0tbfug927n4y4XabzoLI0CgNq5iNrCN5xHzfvUjZc5QfT1s
CahmsJ6Cq/hp1AwdnOKdvpXzWUDE0ZkRzWLYBOdIqi1wvyImXoGPZIC41pR3UvtBOeyp0LwLd1JF
I3ERYWLLTRo4lmL/gSADmZSc9Qsgv7jN/0bwLE8dDpeR4nvyCkcyBN702fJKI2JzrnyydKZ5IySZ
MFyUDqiNB3NJW8Mm6YySZHrYoBhL5m1Px4gMikmvwbgluRfRPTQ8Bwp/locm5D/PlFRRzXYPfuVw
4QfuegHQMuB6+WlAZimtTA5dLc8IkXwNHKuzmEA3FfubMXuOo+ozoDwxvArvTgEmBQfaI2tOv9yO
NdxVNCWT4Oo3chTrdJYlqqsTfE+R0X4hl9o6EoQwhOr7BvgDRVMlN5ATIRZ70Ilq80t7n4UJ1JID
UiQb0x/M54KQwpgJJrR+htqOdXYNWBHTmN/UnANN4GI4OosQYDnEfE8ssw7+l7NPMLDLUZwL7HEH
+TFhGGoITTaWxvDCpASDoIMALtuxpFPOlTqpb+PT4g03QLat1BTrKHI5UCIv7rouU57xJULpObr+
rXbiuITpggDtJ9SbsHZFYR4RSEUw0ufCKUy6D2E+V67emgMeG98f6Sonwx7/tVUW6YTC52NiE9p6
lYsxgM4tz2GK3OkgccPFErYymXjmKi5Uo3OAQwD9T6xtSjg547rZUAWxv8qmaFIf7Jz0bKTUToGD
JfGpJZzKSe2MXFk24oFengdtLY5E34ej4OiRATJB4d6EmUG4OBM46SRTE01+PSvT0k5mRutlERG/
KqfQnMsGWMhvSlMHx8bXCvrDcivvAqskW/2w1Cxkmsf/SgrPWW6yL5Rk1bcLGcwfeofO2lG3/7iG
HGqSjuyFcNsAQgge+9gBPIItJ3KHcr0PJc7gptElnbH/UiSIo/yFbRJARE8WqeXLZrpfeFL3FFzt
hqN9c+RWeFKva9Gx/3YP0Hp35BAbwOzW8Vb+2l2EpLW8tknLMSwV7Zqu2l8hH4MmXZmjEykrQkUO
wQyUHRID8cveNGaEgyD0sv/1yA/VQ7NIdiXDV3g87SK8KuCc1ETUdj02u2o3XV9i1GuPPIskH7SN
XpxPhfQ27FjDxGRZM4hzahniPxZlD8ommDE7jd/wv4bw9tefXpCZGBRQHmm5mz3Le6vQHnso+Gg3
kzG30RH399sRwnwnUzYVdby/Jz9w/gjB40VdU6dREXFTbbLG05oULn+HsmSBEO2i18tBUfUAfNRN
hAYXVAnc/J8vDC8TzCoEK85r+iVuqrGs8UEmQlfDo6kg0mhRW4bdQ3YMFMnADbuv6bBFHrcbO/Q/
MQz1wKPh9qqqs4q+gXHRTdl86WhHXeDPL3unBK6YmHDuc6UZBAPHJCnb4+ov2VWne1UEkeYqFn4a
UA9yF2zanJ//MGb3WtVS4vRXbSuKe+C+ORoTEaG9feZuc/nIZgHKLTXPHK0jSixHc7zz8JF52l/6
mCoOemCB8/VMdnKlUCKedBWY3kvG0jxB0u39tXZmEwC8rAdA33PunWoQ2AITrnCj2jd2e3gS6E9E
qPxpfLrAsAKqJfzs7jr6R76di3gOU7XiPawvz7DLNe64AlkyygpnJPkiFrtecJaEZLmQLK8XD8LE
r4sLQoHPPQOnfbc3qKYZxdupV50vEiNXpBs5Uc/YwLA1KfJl8FLrfWD+VLDL7FS8wc0JkNpKogyx
puUXr3qd9aNgEmz8+i8rPtBkli2SP692fRxyZGMZachQBAZOg8GKRbVphYAQJyH/MuJqIjbjKNMo
LfecwolwAQb6CSkzS3tQdi3bUj1rZ6t/5asFtmcIUJOu1pzaBPTfn1LaNFpetN2TEz67RHXDvxPg
6nPE0ZS6Kk4PWH27WDlYEzDZ5BcDpEoWHVtutZukH/j2QLVBMnWOQcS5OFyzgiY4tASPqsSjm4CD
dDUKioWLY8+DBdWDmPoUATu5+HxlPjsOH9/LAXsS8oi4Ni35P8DNQAeItdsHMsHgdfN/whU0PARP
kzMmz7z1t510pRa7R7Xn65QXng4j8ePsF7vYtbA7kCIX4nHI7Jx7c3oMM63xC4LSNchYAjNPl/tp
M7DYF02F0nOs0fQTHSRVVN4MX+f9bx+mKyROu9TeZt2Byb0uPnDL6dXo5kZ2ZXI6wQp2xQivB3x5
UQLpfYyuoVxQWvsuavXQGF0tRpAYrYVK8+z7AjcV6Fh6gmKsRogkxmOxkTDgNrk0bfE8TJ/30h6U
5SOcwCvB9Nq7akptJiLOjXwfmqTsCsFUVNZSYrszo381t0kTlVDLGiugG/Qfw1T1HfLKxt+42aqy
6+Eyy6i621CDa33PtpBwkSBCvq22fj2Ldid8D5oYNRpvqFcQoggCWpplw1o9YJ1Y053xQG2sNbaN
O276TUdznwSqZTLpdU03+vp8aaVlWufY/2YfLPKau7MQeFIU963R/44N4Ao++iN6CI+niVJuzX9R
iysEQqtvL1NEvXR4qmbX0HuxrS2IulJQRZ91uhktEb0C9da7uW4Zv/C+bNHk2AoUEsROGa0WRz8W
ASuENeTG15kPEq0JebZ2hkKApY7CCy2h8+YnG5lr+Phnorcjtwny6MZEk5RDUgD9HDNYmo7vPnWW
ZJZHGInEZbFYlKS0AxEs/1dvGuk2NZ4ssaOcF2teEY+B15zT9Hkfa0TcpuHcE9tkJrXb/DSr1DPC
wCP83Z/sgufoPL1JYQBTZ/6W/nhYjDkltKhtcksQqVmBgyD87l3m7e9GKmGCiHWIb6o6m8L7ps5B
Sm4fmlv5gThizXho2K/pfLxAcfycaMvxvN0fB1tEj8V2MnOJC3fO4TU6KknXJxEIzJrV724opEou
wB9Njtmi9SYOjgG25RGbFYBXJektBBcGC32DxW4a0Sb51OqEusiwHeLk0sZK9QmdS4eIWreFFThY
zaFBb/VNF4KbBnf66CDGuldaG0c0pzg/UgGVGTH57OgHlI/McRfs3sj80w6OyITwBsD0Oc3HpNG/
jAT8BEVXmRXPDsYqr1dmS/p3dLqRn6sasEqmCZG0qGZ7773rSS7DydhP0c6TIlelnJeUoC1VZuSA
/yhWk7KTNPLah0VnJ7dZuJxvlKkTyQgYIc7GbsO4PsblEeZA8LkP3h9JNM+B1z2n3yM/QoyVA1mp
07hjO6HGqK8o0E0bozOaxOAmnajKGL5/ZNEFlYvWFaT/7BzYlSgIG8Hj2WMZB771Yg4SIDP6W1e0
/8DVU7SMAeke8E2ItXJHRCNcS7BM/hru9bKNlY266iWbJM6UYWz/d+lB/AhComYSyICdBK8Y1yJS
tnWTwPY7tAZotdqSQi65V7vNqg4WEmxVkLdggXX49cuHEoZjbLbDSFthH1/heLdMs6wI8MgQAicS
Wa1ZXQSKyiGfqwSbtqAXgd1Z4HYN7Idy4R0uuHlSVqqBAow3rShzTUxdSlWBiy/UmEebVGkVvWsT
DjXjq4J6L0V4AyNsWthD3vWNoIyT5JDn28VSnCUTwctlVzEb0sUDB2WrtKcfRUDYceniJ81REwxG
X94QR0QTQ66s+8VtZ8go73Psuz/kUmRWVVrl57qqTCE2iCNI8q1lIlNKglIuAtEQ6uy0QY5EJ4dp
Yd0/qWjeO1NUZjKV9JSH8A88opvmFaBcGutzOVDifkG2BpqmAVTbO4KcDXQe2AwWZzxD58RvrLce
SgV6J0P61PIR/IP8AuavaM1wRDMwHB+ACVHsmvFEkzAR39lQH4wnvx14OKP48+TSNBKjf3D3DVqv
zxc7Cd9Z7gSbANyJIgweYfoKLFUbgSY3dPTXo5cpPfn4psj7G4wuPfwZJ1uq7L1S09VItzfLFugT
WdIlrjTkdsBUtF7X2+34JyS6kJhu1Dk4q9pG8/PFD8jX/4ctJiAhrnPFMSJpRddeGpfzFSmRicHg
m1vmcLygS0JsYEGgnhdbzdVl9okWnThai7bge4Q1OinI3yiVibgEzM/GWA2Te2rioC5IuTBnLvSF
N+fwWzVNmJ0l+NZH1xt3QxDsZr/SHUV75hNmZkStznip4z8XjEDR4ouy1wvIE7DYouEsua/71SPO
YQHYZHNxWXzQT2++sTeKGs5vtZXwZBuyCMM4+GPtr5NpJD5+pJNSAb/itluXIMFAVeXgabBpwavP
xjKUvKISpAZVWb5+Tj0WDiopHGg9lqS8cioQmY/h/BcCNohOW8h8ce1hsmkP7fWkA51U6w4bOimK
0+41GG3nm1BbcA43c25SMG3A1+V1y6qfLcI3fs/fF2QM49GbragBJZQFir1h0T2GgxBmPbtE6qOf
u0z6nlV7OqmSP0r79ltXmRnHCK+k8iisrjeTLwhEzxmz4NfoA+GqJ+sC0m0/uTF/pvPbqKkKW6k4
udg16ELKig4V1GTkxVVTnlXmYGQU/P3nONlKMNdUli7NCeoM0g5B5XSPmoPR+fFLNMFynfNR70Xp
oS7JGU+zy7Eo7AboQVEGDdBBfaeXy3FAdH0phTj59rI/73wSFn7Ai+7TI9mGngtzzsi33PteOUyd
2uVdUerm28XU1cBi39oNawAFUFfnEiVsddN0tw0UIrDmyMLlN6dDD3zeBWD/0GtJ1Ob5E7auKqCq
Tc2j28eypGZFppVbFKZ5ZrykstfsbIcgXvD+acffoae/0797vaxSwPSgr2aYeSFSMUQtVXaO2Xgf
JdZu2jC25D60ee76YcuUkAGaSEdPHboQJAMYp59HA82avd/soaN6BktCxWp1kmm2fbvVjvmNlFAV
eIUKk/YGZgd8z0DKmUaDt+vYaDHPbg6sVa0S/7qEh9J1DXpf7Bgi1wlvO2BPoHbl1+x1Z3du1HZX
xv7xkBU+SdDVR0i+dwbi/FgFzVS5KjtMrBMNkzaZBmzFs/I5LRrXeWfi/ORQqoNv3qK2aZCUlGdK
lwiBWCrtH3wvKDhUntX1Laa8LZmRhXS9guqY3cJ1PLafKo7VxLXJ0mLl/Id4FRylPN+J9WT0BsLW
qVkDorqY+/FuxPXXG0NhbkWSn/w9FR33QrHRehdD+W7wDMywxkidnCfT+hjmevK4VvRATW8Q9LFI
effh5YW5CdgLLzf3zbPjjEa0IlSZJtAihnx9fa/i0C4Ua3mKQFWU5pEk4ICHj/h1ytXFVpDeI2co
ezFne6prbk4nJm1DOLyDWaU41dBMtPSjQDVC0+FrIvWVDBMvjQ9kjxYiso+TwmCaG8TYJYScWRrm
UIOcC5mw1XzaW9qCXsCFMYVMgDj/0C/xWUZISgpKvwrb7555uzmHuyRjusj9BCfbM1AL4eKUbtYS
IQusN6Thu2EA3mWCvIk7rNqN1qgT+qY7ieTb586ihBGixul5HjWKMcmsdzFRcm8jecknEoRSU7Fj
hibwNFCuM0hj5tuJGre6hfUeI/+9fhxc/j7JN/qvDg9bOApOIMq7L/fm6aXcGf87SCiY0MyMCPr7
qhqwWiL1lNIdYY6v1XKWqin8dFHtmDrFJi+CDF5Gm15rq0plPdpUdw8XL8EMwoN/zBbQWUDKE+/H
QIF4jDj72VCqdBkQvTV6jSsiL0jNhE9Cv9gCOXLZfxlaYOGMQO/dOC1plYprGoS6ejCapatA13JL
fWBjCBBstjHGA2qDJkBnATqkGlnRe8s1SRjnRkPCqfdmqWhdZiGVooihGXo76j5Dt7nI2ipni5iF
A2+PuMEu7n0kgoflIUWxxWUJ2omwcAjekC8yiABTXaNgc13KFrCP5xsrn76LqX249Ft4gO3gPHxe
ts72Ppl3ns2br6MLRwj2t32RPja2Swsv53v39pDPY2RKrakLPg2UbSzBvO/4GafTNY7lkpkadhKz
+x5yXg89Jv/Zv+9G6nlPxXPANlt4IDx2qpbIEXtiEYaWfWwWZEvJpzJwbk6Dd3MYcBUNWuBs+G1g
cy9wKXkaTPVlh+TckXRTxSUCh3WQggQVik8ycI/Ccqh0u9m4LLZiI/t4AVb3IKhDOXvBFKYvJL25
sNZGlImVM/CvI8vk9c7KxaFfg8mulHLkItWdT51F1Pu01TWfxTmphCMZWpjP7Z//3WoomnAGoPOm
So1P0KjicUrSeYDRMJl3zcn644/37fo6+vnvafL94fytDF4DD/GM3RG88/BVEWwrfRRmuHf4tYHs
q9vAItmSje4LmQmhoejVyUQyJBoQ5fRNSexxJoLo4RIp2j9hjAT3F9KFjNfbPZ/mvM2fVzacKwmi
AsFtqofydas0PguA/hWqu1abPNAvaTn9hyKQnBjypJKAWo1oXzfyUEiEh/fumG5vwE+mGisRo39V
++WQR1jewMezbKGvINpO5sxLUi0hiWdOFYc8jWfR6GVnetR11YaLjuJ8T3RRf0gadkCC0r6vbyqu
4RcSMR1zrI6nzv7FCGdf9gZ5m0HZ1KG/qkoZRTiTFqeNUT+NYDmIFDubcQJlAbjIcPTubboHQ/ez
btKZgjYtCL78DP5P+MJc1nXtXuMVlfMCfAShUWt6cQMsMjBEPfGd0Ip3eK1dhylaQj9lsqt6hTiP
awhbkKXLoHYShhV+MFhun6cMVOQcQrbHilSBUGDy8AOSVk/1ZnrzchmxmSkwWBKRjCSruZAH464Y
t5apA4woUxLVmx3vcwJEBvz2OfrQTVt7slh5Z2OAx2muigS/ycS8f+y6cMp1WhH1OPiAe1gClXfa
3lWk3NJTvsZE48BwSb4Rz12Dufi/ailpnJUVY5N7it3bTfRwv335NTB7E0qtA24oOeVdaZdv/iXP
m6NzLmPt2RnnxLJbwq/nyOTxnxsTzZE1LRqvoeGiekBh32eJFcnw4mLhSip2e/L3FMImIfDTYaqO
61oLR8INHycBZSC4bOokCcpyYI7SvMFPWk8R8MwmSnOZZcF8B0J4qKUI+yxX7AXzhXLXQoJ0drGr
PyUaISe+bWwVUF4BpBplGM4zltpzLAsPkQYYtDwH0lkb/XPM5SOMtyCxjJtgTfq1x/Bb3xTdVxk7
72yEU1YcxbX/ysvgFYdMnRWcXgKDoRHHbDiIPCJAaiXhuXg18LAOA7kAMstBbUT8OEbALLGBvfwi
Rofe4uHrNfsftgM7SJrPX265538siACdXQunBOkEYZTxWUhIIAf30qQw+iKgpfD7unLQLoVyeYbY
vm2a3mwibrHk+rgRTF0Dwp3utljDpjykpLDCagg14oMb2+sw7NLam16NtoWbuHAxTsVNzW0ttssj
dDiaRny692LttEPjPN/9yW5slPy0wTVEQx1wWT0IncOgs5ZXqpplz8U/lUugMdBJTI0p3Nv+8PI9
97+GqHIyIO8uuAwYrxzi/XH6rNYlhDSxDfnjqHvGt1vlg9Yr9al90IByZ+t3zfSmsHXMjAjXtpNA
E0G5ub+TZNjT4yGB14gzWzMDvtkmxx2UJqOMD+HSCCUJUh2Aek1R2M/JhzV2htre5WwFfUKvkJGC
DaStN/OqC4Dov96oM8KwBILi5kFwDeOAmea6FqSbS0iwcNsSoFNPx3Ys3Qa/+K9D1M8JMSiGG/ys
vwSDkPceM3Q0lLscI60dxKfhETWCUq4Epil3UU/v7HFv8F8NIGTeSsVWgiS4FFT48h6n+b7C6URa
MWsHEEDTTiUcJNugCKOE6Ld8T5FOJOdGYsKcRQPZ7NbguO5lW0+1l12KYy+4x4hEjUrCmW4Om6rS
SnkF7hsY0e/TX6LvuNbHmQJm+60BbyENKpJPqNe3SQxmW7oen8OZODpDjZPoop+D3gJwel7/UPPd
dKVCyF4dk5sxHujcPff+uYpYEEsczhooMRXAyV/Kxw7Pk+gHSLiqEZD7/o8tRjFMC+kttKAy5i+0
9occU5XDYeoqguULdw/f73NhMd7Cj2aqYIUlLguwnpwyKnfyj6IpUuRUUZnsgHM5EIOzWMUVbsVO
Xr8j9ZuOt8XPlezFGa5zV4URHLPsevTheIwIw/Ux7aI0EK5UCxHMGA7iOgP87c8h2LtUqv1a5OYn
c6gqLG5M4VuteiNoxSC4U7RmEQ0GI/meKNWSRLM+SQ/YpRtNrf5+JPNfiMy4bQ7d4AuUlfWqQODh
pO4EL5HchRoiBgBggjnc5QispFsOpAKZrAwU0HJ13cCZq/94Q+59iRZIP5YG/CLfvY2bJ0pvj74n
26v9OaIEg8byhaR7rEReprDxduPfoATQwHBevKh23Fiw8N1AbVAuuCav29XtswWC4q7JNHzV21GU
rJIisOxpWb8qtX5BiXiP/6dF/iZU4/kjKAJbdUkwD++54UjxDEZssHwjX1OTh/rz3BfK+YQJSHhE
ty2XW1Xk0mocNbJ5zSQtARrU0c1u72eFUzk5744HUTYUSZlm0TsPxkLDnC3pO0Rm5gpWbTD8SlOE
/4RTQ9FdhvNlq+M7FYXroVM1vtx8CciYLqxsZYgY6MTMsRuIWC9OE9+f0byzTU0yuXfWUioTC104
+MK9dijfOyRv0FN6gVJo9R87zdZxS1ZbfMJiiOn1+XyWYdkdUUot6dlVnLfkQP0jFNdjXHZXt+xa
eVIxlUY+SI+gmsbBT7gk/zrmlZ6eLOUUDJTaf0XvJOhKBdliYWVKAM4Z/5w7bElsyxcb4Y5K8yy9
OkmUZMFKXquECNKop7HXHMRmEhiui6Md7LuANFyCPvG8+meZ9C5MW4w+vs84EeiiWJdyD50S5a1u
29ff7OmcGdU1ziSROaQ99qANKrOK/rf+8yAhY959EUOSnhmzsG3DFI19FDW/IpIQI8qayIr+0kmM
c9Y+upLXU3QKFFS6UoEXtCm2ryLPvRKD+lYe+Bsmh0zLJTqZiajhW6BNfB2IRauLy1K+ACfewD04
nSfy4fqlUbWoC1OeMGaRS/ag29QjUFiNPkOM7HfN3rH+ibwD/hngAyRlxgYLXvg2Bg9hrt8wFKsH
fpYRyNDAQGT3PGDERaxjNFfNf4hfgl12rwC/NFzshbLfp7VeaLb0IUu0hSG+ckzwbIAbBM4ppXnd
LjF7BG61z/+OK256gWGL+EtAPBGJo+4WFwWO5m/9/zUcwNj1PLl9Oxjwc+hYoOoxHAB/1sZIp+6n
8QsTAQ6QfzOTukxuoiYiHTTy7/1//azEOwgdOoNSFrr1s8N8K6r4xIqB5PRwRveG0ACBJQDtFTad
p5tg4iIJuPs5gYrbq1KWVVz21tobZSowuqH/HOJWztLcjAh69V11CeBYjZ6M4nT1sG7uqe/XGffI
7jcPSoUNA7XJ7C5CXnNHbAuAhT/oFerXVYen3NKpqgl+e+lfXOnBLh0pIFsrWbPdxvphPiwsuRf7
ZTqwuJ8bkugIoFYVn3xlByIaU92jEYSpk0qNOunF/EhSdM+Cqx22T63PuNg5sx63ToYLfuempyT7
0+GJONPeLKdW2k3mfjQIyHW1PML9ha5mHUW9KfyMWITwC9S81Qm7UlLT/c0IsZmBnxclQl9PovIx
PEto6MfCMNwwJ1rvyjprlcw/sI2Lg3SP/NmY4oq/XrYKgXNiSIgyJ0db04XBqPNYq+bwCxcxT3MR
z7v0gOPwsqKppZRHmWofZjeiccyz9uGbMTDIF1Y8SV8VgzsfB7gCpaFMl+NSwmHWyxuaBHITOL1p
rJ/0RTOUGGKpRbNguSwpg8EK/x0/L7LnwfMJMERfQfDjF0z+aQn3YDvGxN5JK6hKgWhnrvRYh9mi
OkQ8x9Q2ajKXezMVyiChAGacppol20vvj2NMdVNDSPOJrnibHUi7Tkek4G6oAUlV21x1QQtqDI3Z
0IEgHtVEFfrnxMYwfiTWdGhkY9j8AT62GrrINAlnEBj2h/J5jJ7RsyYVhzLllfaLBET/ZRbLl2+7
sX95q1KON0lXubDo4pg+sigw6RrcxlyITtCpFcamo/AD9SJIjnM64cwQ4i6wjAQwqyFaCp2TJpk9
bi8g50pNiFQXQAayH0yxNn0jiqAgwrGIt7rmTIWmkImT/4sFTYIPhYwnWf/UynLxNXYJfmjRmUqN
y87iHnP1q3Z5dkQSzCcpyiBg5BvhLr5cWjocBb4F4hFxsSOkYJJx2XMLDlP3HsKB28PkYN+2rfIs
Nk3CgpDfjmuiI6CYn0hE7p8aWsIV/ah1bSkfN8+1WNfFSFAVPEYCXsz6ZViNrkCPjToiApxPJ4Tx
MQ9uvn2XaywVhGTyGquQqZacRlezkZHcFntceCX6pEqOxo6OdBk6nVSUt+5fGhGW4XMt1PV0+72d
J1Cj1trKSvgDyv4P69OpjUDzY6Dsii88rAtlZpSjOenbnvSlw2Zi8Ak1g+66yPI9A2bNQlzUeHR7
+3B69oxVmZTUuOvcuweWcKK0P+/2SQVpH/QOoqOdtzlKU+ulmZVDiZkXz+wGfOq2HrN5oY/8i6EL
m8O5/5JdaAXXBF2UeYuwfYMyrLU1GV677MJSsZlgUuW8bP0VdpStZOFuGAWeeEUkkR6+PP2FxJT2
Gj7+tQxoXPVRCNQl3R2ybdbR0bWfPzaa52pX9NYQGrPZ5m8yVwV2PXd6rJZNwK9o12fMI4h07pK1
xCC/YQtyK3di8e+2XBUO871WtY1aIPPESo2D2rVgcgm2bMS9Y8+1nMrK15wKRg4D9mvIFJE39Der
1x34AZEHjXQtFydQLcrP6kBZELmUPqpl24TumSClKJtoZifgaqN+3B/9BnHfM5WoZbovubIjslSn
T91+2ZjBrc1MdoMuTaAgMH9vMGAE1HjnWz3bE2Y72N6RppFxtvU/MbiSw8yRCf4UUmsxGBtdsx9l
iG3Y2et534YQwU1IrwDIxPpCGk6sSzxm9PlOkr90NgS8j3Sy9aoNbX0jsLgEFZbBroKMchNdE1V5
NB34tAwiG0tTACFnnG+NBFDHsaL0uMoIVUA5o/e30k4ueAwXUupPphhQNbtqeKQ+awTqY+bgErO8
hLfyT0nuSYt53u6lKYfANNT0IEz20ci8i0e1RFFDwOvNpFF4QT+F7fS6HtF1UdZUfg+czdcRtRGx
HczenIuNjX/1SLS4WZG2DkKeBa5T46B4chdnPBAylyfa4N56YM1NFp+rDAma3iItI5NPgDLJoDgN
Y4XNCDomYzsxbZchd0dhNxDZZYa41wzdD4IwaFqjVu7GtqeL4Nn7BficYr7dV7X+lcDRqB5VXita
17c2tzjRhkr45lK57+0dI5GhuIHC2FmrBlf9KfA0kPY9QN9Go4DVjM4ORna4/3Nq03og5bq7GsU/
nMp5i2o/LlZ3u2NpryBmEXNCK3744hz6l4YltbGNwrYVn5ep32z6vR8gmkPfDF/3xRkWJg7/tOO/
kpFwn8kORNd0xMBiPgq7kyr1iBzhD1IA+gr+V5Zz/66tKHLk51eVMbFHkmN1waREwec7bfHgT9PL
r6+4yeDkPyQzBpMCW8BZW+s7xAqxywfqZju7aVRA8AzJEtslNU/LaautXTttMWrvoaWm7n0UDsGW
LvIX2ymuc+5moGI9Q4RZtLL2SKLK9poLnigZ434Y9Ha6RwHx4KBS9ZNSssMXUaSApRpq+AP7y/DO
tiaqXsIixEiryPNB1oeiRxRTK1El2ZZ0sOPQ9ACSm34vygvJH8jR5npnN38otkIgnZsAWzE4rVM7
XrzoWDZaQb6fuIg4kglbBHg/2s9qDCx+Xvrhos5RwifdklMgb1WGWMsoB++Q1IxeVoj4z/HAM046
c2f33Wm/FSjug+eytD7h3NrXClKu2UnfJEUJcWN7YYHH54kg8RzKoKVxR42TY7PiJKIMDzyrQG+W
tjDml1dN4d9aCFuzbbI8k7zYmMc5L3IE+/maLOlYO8L3/I65odMRLVpcHp9uBZ1pmR/vDmJWOpI+
aeG4kOLCH3KOPnQCX7rcsw8t/WdFrYg3X/94MP0Gz5IXikAWpj2oww0Mr2ooLZj4je1GbxAJAc1g
Px8fjhJHlzrGZ7pE5EZayIOIluMAfP8Gln+z05i4QQF4zTTvdqNEDmigULvFPKEUX10P51wpupd/
FhM+Tw+KT+1lajHkZ3Xx8tIW6Q76SH9kFxb0KuQ/1u0m//+vmKk8G47ZH99Y6hJa+ILEauzNmKWm
olpAWNfgSvENGrq5eWh2imZzP/UXazz7yfGNxaEhOaYszQ8ENacjnB6DtF4bt0Vg6NfHMImlD0Sl
GTLXtvgBqM9rjOOFCLxp6LVa737NFHEr5d9psT2B2911FfzbuRxnbKeuQoaWkiNDzzJ2h/u10VBX
H+fMas6WH9ermos36FXQ6KkhuhdWqU3UtKCSoGeSaWgrADhHyIduHH911x0PjLEDXfus02ZrllJW
0LZrQBtAwrZujJiMG+QzL6ekbgRtzuoaOj6FXkvUwpF2dGPRcduywvyA30TH/C9m65xK/jJ66+2Y
LLe8mTQ2u/1r/RuaFKDirAu2jS5AFIQtGGLC3KVH5c7g6odfviqf7xprRowPO1pu08w2pQy8CHqW
G4BRYo7Aqb5Y243oth5g7CQSjyLXeLqBICbOx0q5gs+Psi3oc2mzRFR6JPHiGTW924keYTVHSYMB
myvG8yPWdpE5EhVz+wUL7oBWL+HLsaBAagA7iPAGR3QTPnH4DY2EXpEcIZEwPPyK28sYEsVSNXsh
oI/3NAnNuyAkeq3yjv2R8NTDu4U32mwTWOfbYompODabJEL227I6AJyRJW6p7eZYSuL9KgPEJTmC
ErojJdQ4jX8w1ZV+EokivOmOWyztgnb0f2eIaoW0/rn/4r5uAPaI1qpsh1nUZj3Sw3CYarZQaeFE
HVxVx0WYKXPefLmvYxRHSb9wcrNmVxk+sPm4KlWNRmwpUac6RtpIXWlGyO+9X9RcxdP7M8DlhqFi
CoaOIFOc9w2qrfw9fZx1zWgFvP+g3QgaL2voTiwJLIxv7rEQzqho/DVVsp6T/L0t1SNhv1mkn6u8
vski3KadjrOq0e8l030kaALQwvNPdQUHlqWO69p7J0LTcxSzEArMK4hrIN5nKLoKz+AHVS5KF+uv
ZIQxdnUaeu8nUBQp35IJPuvBhRFSgZ3o6xVLjTUxWQk5b2dd9kXR/CWndIueW5f9P0BdfxKYX7qE
nhD1dmvHpvbB5wOrzYS8EQ424P86qDODjp5CIhDGT6M8bKHlJxWZlLon30SJu1OMJZISX7gYPQYm
M5abfjIbxRJVBKFUQZRbvI5eAmhMH5P7yKuMierzNZO+ca9liOKtHqEnY7SuxjzNv1DTtaJXumGS
VCnwt0K6ZkoGYT/LumRixyaWGelro5MfSfisscgBZkSAAlDkpsPiMJjhh1ZO/d+MLq1+kJsLaFGC
/fmElsIB0UXB84gJ5d5/hxvAvMoKancWp6Ji/vOqI3+3cV+eNFjlkfPFw+9VezMWD6mKpeZSUV74
Ls0VfoEKxC+u3S6hxuprBGbkeFM8r6nQO1leBqfArgBRvVxYG/05sR7TwtECE+mr0gQJynrcOkIZ
cXzMO5rkG/kFTAj9htjRwD1h0P/R6l5UABM7ro6e91BFwNt5EXQsoFy5wY+eJcLnb1XmXtM30LbT
tKao5SdmFmCe8FuHpluZO/SZ+4StGYAe+2Uos3yfMeYa3/900BC80hNO5JS7Qz3smxa7ocwIeWFg
D8jOq3rmsjT0WV0qL5x6dkc3VwxOmRK7R7aTchY4jH170s4OIYRyE9GFTOndWjBliGra183seApW
Q8/dD+rx1WrcgbqW+Ldxyc7B9cSjolJ1oWxlcV9s2uinJLpl2qAOYr4nyB2m3olM7ANajdPsDfyB
iB6NdPwRZz+hkciyS+MOshwyeqAGVHPUWY8T3I3GqRv6myJCRTrM3vN3fshglyOdyQXKX9E7y6sn
/JpUQNrYa8RBi8WJCqo4nzO9sGX7V6TU8fqXvQ4MEbCCdiio1TDvCdY214gPvmBFK86T0/J4s7EQ
RDKr829Jhu6g52PxDbRbSZXDZwKNQu7CA2xl9QRPBti3mkyQCoh8oAm2BN46zSwN8Jgpb8/s3X0P
WDSZXcFe/9taTjcAxT1f7awZ4kAryYlirPPXOCdOfNXRQEUXZXC4Pt+8xvM/aThn00a2emWEU8Mg
lYg5WaEjBUQYcVcPkSd769Zga8NNEUA/CucKX0ShKTFboXoLX8HthvJHHmdISrOWsBGo1E5DsF0J
nKvf00DDx2pdxG4E7oyJ4XWB6cYT02hdqMmrRlye0gwPc9GTjOJ5A8VPYc2we6aF9WixCw53TOUY
WkrNTnNYW1AhRY3C+pd5Jz8A3aOHIrfWJzmpCecJXZtvZ61UfY4Y9/JIT8lFgucrs4A3urLogBUF
MOcHX2CLcABjFDxguZ64F4lvFJ1CsMQYaG8bivF2bInsxmqYvF2aU5BF9XnQ/JW4NPvDln4gSF4x
+RdGgjR/I6DGxLYC4j1Zk+aghuimERhfDmiM/8d/kFb05Q1hXInDnqzLmdvskUtZQiZkYhLStFoG
shqkTHHg58R+t0vm0SaBeaM0oaxmoWtQ0hdW7+qOhRtFcxlgbPuaHRc5qUxGMkVX6K91kF4UgBP2
XJU/2IxfuHZn68+1jJvv/RC9Rb5MBSEWuHVsToMsmjxKyMJTTXC/nYFuPQBgPi4rXcF74UskRw3+
0+S71qvWGEmAToo++Laxn5ILkAKxD0XvV0n+1MtiW/u3jyxoZNR/sjSITxqTPMPQB3go12ZpOO4g
24w+ChoeGnN+hLRyYHsWoFeIkaaYyyyEAK/eAHuD7ZHZMdxCn2i5+zlJx9saq+41xnfo2EZhLoX2
Hw8vrQ9qvUfIZI2bpgehe2m6CV9frW6iPJNZSdex8PeEHLH+8NvZw/zxCQp1iH4K7Bd4CNaQJ/Zk
2xqcZl6PPdgO3jX+l3kiLt0NhiIg0mWYQocjDA6/JtVxCzUk0ZGPxueQhbupC4lu7kW99btBFO28
zHV9Oe1DIUYci9puG57HsKgL6viLxf6xLFnUXeibIbAZ7dUThZAZreGFOuafbcWaboyM+S6NiYOw
S51S7B6whGHrbT993/itWcY2DyHcljGe7jCM/xcjdGLx3PIWzxhX/PXrw9b4n0ckAZUlFot64JdP
qo/Lwf2rPUZiD3LXr0Cmz1pRnrrSl/XPnTV6Wuw1NxLxWZ1+r2sculBwrbDgl/Lm9sB6wWdec11w
C73xI/mo+rg5Ft36oRhlb5FSGcVp4LX/7K1JMuDnSDFNXKlejPmyY75EkNTknix3WgQHhR7SBtre
tiV+5rvlyDGRreoSmZKTwAd7BWVFsewSv5/InuxLfCgwU0Gd6RGgrANx6hH+vgyBQUqXoFmBueBu
6Nhef1fjH2s44AZLtoy98DrJEeBkGeXXHXcm3KXW8mKfOjiWsYa/VpJplBae9Ao59UK20C7QMTsk
xqLnBafXLpz4+2doc0K5/dYvkQOrETV3c8oMDuVNRHbeDwBxDoi7qdA/Cy0xMvhEVKkHCE6pKxGu
cizZGSldH0+0krCy2fkA74Fn/2LaJzoQlgxrBIYTlgWX/yu36mQx87NlYc6BxZUZ2/TfwlbL44th
MoU9CXERBKM0NKZxMmxUP8SBPDbaFlWd2RoFSgCWxpcuwZ6uO6Ujl6EiQYaPKRoWovStA69MrPUg
rheUsCfZlRnQf5YuB5gVNK4ooKskSGFtSOZU4zcXr0tEcVvcBf9vExXL4SCpNAZ5xLeibgX0rhuB
0vG1y4AzLS/xM6g2iJpCdOBiDBWaXHSpHntyef19F9Rt5JbWS9h2t+EiphckQmROLih0LR38E9Hj
7PIj9D+YRES819uZJb2jRfQyRNB6aOuoW7wV07TEST2WqWbwdlN9oqhie5IulaJlUMmHSshpl8Bh
bzDQ/uWDUZ+kvKfrONnoqEVKw5orHifpb2OmCNhqxCOUHeCeKr8nOwVYeuEkJtOmhkGSQttuPiYm
Gk6PM5D/aRWZryjUtjpnv+Qp6c7KDzn5OuvLl5ZMh/s2Q3CmQNgzjjHq4F6NLlthVw8IsZC6FKMD
iyPvcYtR9eDWJLhK58mW+XWYt54/s/SYlKSxduOLP/Rsw0KnMvnJWZwPIYWPwchJDlDWoLiSYjnE
H5woqJVnH16GrsDl+aKPlNsMLJ+wEjG7dfB07cfsTij/VjXJeBUcSnZjcD9QT1D8kx5MTRQpc00n
PjTggnli0igoYtdNvZn5vaEgBm3fzOVEkfNf4nDxIzp9F7vmwTBCaocmhE/i8Mc9ki4XKZt8KjgS
B8G+EiTvgVf0oKXkEVE2zsWWdo6gy1u/yv/4KlzlTm50wG4i0PVYMyFtnsDINSHB7sBUwuK9OGDB
MxQ5SRKUr9h0/wTqaV2Szwkyp7Vb+9Icwvc27YVPkmpqkXhGjFbPP5dvwOt3uYS+YRoqXKpb7p1R
/m3LG9QK3eayxMSFneBIpUGs6nUk4JqLaHx9U0cx8l2FOe9ewVaiv5WFMBYEcshkYbpWuCRGU5sw
3FxzcJaGcOfNpxGFCSkZr//7mg8Gp3ae+VMTJ0tkk255q9Nbfy316AlSb0mCJauH/hVtZzLLD+/b
GLKEA2FmLlpWLiIJZOo3PT03nlBTMDSPS3njP2189HPcVirDA6oDGq3vHXVfvZq8Bxax+VsRZrTW
gGQDKJfQCLZBe75FNLkujYOZA5iI5U/7SyIxbfTtz1PvYLr0HBTt/Fyrp5IcmPLzs2qRg1zLd9TH
anaROykZr9RSabZEO6cY33CptrNEIKlANh8rZR1ywhDwCoDpsC4i1Q5taORT6Eo4Sa7YjUyfDk9Y
gCZsmn8ax6B4QVdwXRRV9YBqOfa3kSlsBbnG9z7rzIdYVVQ5L/zpSgj+P5CZPfOZTmL8YLus5L+t
oAp3UmUe5E3tOTuIl4uGGIoJMQxmHbUfKISgNoMW8UnWIZ743TGWN7YX2Jat509UMn1vMPh7rhcz
S0XmMvwjv0sbCOByW2wvq4pR7Ir885nq2c1R6XQt4+YTG9z9/P2mOGnsLY+1VBYT7JjpD6VM8HHj
1pAq2aCVxS2FT3yGeGkZ0aLqJG9foaUjIDjeI5QF4XcnSraMKqrG8saAHys98GWwYsVXyFN2/h1W
CXN5QYv7/chETlxnrADNm5TSbLq5S+1yhjVSuaHMGI+k0Lr0ShylHik/oYRWEdcuG8HRYWMqj70t
4eFLfpgxrzF1WCPUHuKUqtaCAmb2+liMw9LK+BqqvIE0Np0fh7Awzj8YoXf6cCNvz6iQ5z9GaINf
804uW4lSZFhfjUlinZ330vRP1FmwwYDO0Dshor8VWmSY1prZDMqMTYs00BLvFUD3ChowI9G9gi7k
J6QvysLMxWxeMqwmJJRevK68pj+rDVL/qYUzDoPuh7jRlZP2oLuj5bi0fcp5qAgyYe/Ksh6RjS7u
uLiklvq39x2tkAsTnfNraFL8L4QqYoZIPdFeh+PWCgCiVlGWwLrItr1UBhtQh1O4JEcDdwDctaNv
hCyBTbUOjZvWRrDV45fljLwIvQa0PTdjz3kkXl+QZrMJjMY0MIR35sQ1FiDSAZ9A2WLGkklcKc8O
DfrudU93ncf6YiyRS1SAsL8rNN2L0qVmeRoLG/zCOKVjvaoAR9u8jMGY9fkPo29KFNn/2VidYkGd
6TZr9P5H9zy6pHv4o4kuZFRuv8uRPpR4IsVOFTOMdwNWZk6q0UaMATLH7bH8uCcu2EV6vjyC+WN3
4/zLtgJuCUdXgyoriV8LT3eUYrhc42a8fagWB/kHI9zlU5MYXkZMiFeuSxFATtlFQdObBmTIcTiZ
etgbtotZFlC0sLUufXmDmjET2/l5UL3jwJv72WgMwJ67riHF+X82yJl8GuSjm77wprKj1xEOYV4F
ReH38ecsVoLNiZRQdDB8zLuxgj2mrn6du/OKbxK/7c4XnJx0vOlPaaGBvyAc2wSAj1QIvEH3MgK2
k4a9fbI51OuQr7qWagiqwAqlYR6Q+DV6MJam88sULpWZXaIpzlMgOX4PGJxHA5sh63+7Fs9lWtII
NuBySgDi9OvZ1Wd7f3JY6STq34QHF1kd5RtNOZMe9gQoBcuDa/P6hxVXscNIMzDeEB0GTj5lcDfr
Ha9CIO7/PkQUgJynqctH2rD/Ho16TsoUvwG3N1oGYDzaOw+mjZuT2zjN4cFhdL0GrQJx/rx/+O45
FhBCcdoh8wOQMKQXbyB5g4EeWkrpbgUNY4KZijepZh8IPPI7bZ+ltc6gSoLG/9siRGpUlLQOmo0K
GpRGsmmKXy6qa2wbLCyYlyg1Ws/kKqa3zz5NuCg4O1LqjU3iBw3C2BmB9H6EbZK7KF45GFfI+sF5
tyrEc1Fd0UEhMkAw3nc9FJG9VDoU5s8EYDwaIMBEEWqb8qDGw3iAF1Vyp9ltYIWe/NgiPxMTVbdI
PqOb8/UpoXm1i+jfDNRYduzUlP8mQnq1+iix8IHXEffoWjfiev3aKVxNkYntOAMVPtGjFJRz66s9
/x7+YbbPMpyzxQF7/3/WAidYVwUv+yGd1tNq/DeHiNga+AUneGqrZoL2E4AShocK0ZiATp9qOaSW
mc+rJZ2+Zjrhz6W18EYqvtSnFiJXBk1BeQor57BtU0LtjerjvUO39V0noKQL06KWnZqArgbAMdAX
znkxWoSDYkyolyHELe2foP9GY9fd8YAG4ZMzlL+DizhxpmZ3R6rlb7ABcSWaC4+jmC/thztEm1vv
VGE8MQnjO48Wi5QdN2ot25mgCi1H/Jwf2gjtXLPEows+ZxWUjIdXoG+5sZcnkbzph9fq+5An5PiN
8lCczLEEP6P9EknEYe1SW5y3WqfWJD4ia19bQOmKkNOc6ocXbviCJmkuBAUGgqY13pnFkDugNMPj
3vKNNgZRcXv3nDq9L6/qLPuVPW0ni0WIsttxbEG43VuAhHWGGUlVOaJSlV0HTGRqu/TYMZl0jM+M
Bzyq7N2fvdUHfGFNIheD0EXQWTEPzEd20uxiJsKiKvbNAOpSw2kb1VOaJUyShdOd0jHDopIldi8e
6WzOe7q+BN2bku+yPA8YYnUjawmZiNj7x3qEx0WoD+3/YMWQ4aN7rH69MN0llUBYxKq71nKClKQP
eCtK3jHzVhnVFcTEF0O6psQSfKLD7emYzBqa3kkD8Mw/SD/MedZdLlJ71stl/6ltShjzieNqfV4i
DskCowFq7JqFZcPEB4uzJbgFB5wmSbaaBU34CtrlWFSH6pgJV6QcIRnex2puWnM+t5wBBmXgLsmn
tJj+0Hzk/ozBDpqkhWjC2uBDL7hNupePwNVb/JuSA9fhWWeE1jLKEwfIpu48Sh5RzAaO3KWYnSpn
ggAs1+lqRiK96SVRXB/eS6jchRewkG4q1BhCOtptBGEqWOWeJLT6qUDGv3J+CDh/KTMCJXisgRji
ycME51n8aRPM83/iReWNDl7EKEVLwfE1BaOFhi8NIevNTdu0H6wlg0CXVVp/OlfsPcr7667Vm2nB
SsMtefLiAtSii2Wy4JWJxdFtJ+RVF09XdhiRkTbqFX35lT//zrN7SCx7q1lqVXpN1BGwjd7bi2mc
ovUHHpaHi6ZKwXeaCb8HV8MlH9qMmFluUkiPQrNk/iss5FWRIuC/gUpzvLxiFzOH3DsjSnAyxmzW
Pe7iMOyTaXaKQNAicw9Useg+N1+QAu3LwdD1MkwXiwG6gg41lvk1mzfEZi+ii9TXPn1q+QT2VGOa
NyYwPHPRHULe5tx7G0TjSR82Apv8i28Ey49i1d02VF9tqUuslOxykRnHMBXHgX8gTHsDiQnIae7R
zXgvsFRYlr67xyH5gVWto6XEJ7TX9sA6N+gi6A+wd0vC1L240TNk9o+yxjflktBF66HV6LOykDMK
MLh/3k2Oy6te5rJrjncusqXtae84NiRmIBq08iB9KJKSPoxM0okoPh5G5CYGpUIZ/3CUFKrAzGVe
osq+Y8iLgk6XCkcUXl01gfobBrQd07nHLPsc9uMGqsPWWdMHUcDm5HEBDxLWcs8d0TOmG671KbO3
QLescWyGHFw7hr0h5jjP3YX6EmL3o+lH4KAmEWv4zb0tUjNIMuU5CIVjJLLB3n/gcsWkgCL5VmFX
ytTeIAMo92KBkON5tT9Or5wGvVio4vlDgjPx/1zTe+eJrm97cdUA0nLu0VE5t/0ZnDM0srasD6aK
ipK0hO9liYZFiaH+QowWgW5KU7Y/JivYuTqqgT94hqYGETjrsLXEE9sCEy30jAKCV5coxRybfY61
Bl+Qtczx615n63L61A5fa6um+qr+8J/sNv0EepAhEpGJJ9JkOGH9XlXjnMd55WuweStG2uffLo/7
x0Jx+eQ65xy8YurjS4bwludAJC4+SDM+twwiUwB5bPbBbr4Q9yyBZu/POK1MQQgkfpuQaBraJcdw
tOy7HASYauuj2WBOedrTsjw15gE0XSZrGCEe6Ww7eZef2n0oxhimO0wzxgPBwBSAO5+MA3QWyLlt
VU4kjPPOLUWkNEqvIPIKnzNl5Sx4TZZddY5nQeryo5OOIFCgnPy1p7BwTMUm2SLaDacpQiFaK2se
4qZ/klteLfEoiADe0m8KTMngKQfy4zjPq/0bzdPnBWlQQ/0sSsl4PUWA9KSYEVoDdKVcjzMthc7V
e4bx0uUI23IdzWTEnjYbJqyxac18DfF2GJD3oH1k1tq9yeOCRe94qTQ86oWDcNvhc1ltVTLNtCot
r/O26ale0saHL7nlOmQHhciFNdRmWs7wgf65+7HiF0qWnqsCrI6T//W5MG2AClzB0l56ctScAny+
yEDgzcBwuXBr1+5w8I8k7/+myDMoWdlIb2kmYV7GLt1nIo84u75SdR1pNlw2ndWmxvNS8aowGsWq
7q+/ECpKsJsN0a8T61LxEeSJFRKOLaSTUUTPfm0n+8nIPPqKAB3DJLviRnBEQf59i8cLB/oFmHE5
pjUIWwRq34IHRyDI2juX3OqZ2h13rJosZUT1hXCi8jsdC2VOkPUwQ/MWNYQzMUkDk2cQQFyfM7+7
B2cnLUw2oN/hNJkbQYn9JPWtG8r2mzqmwM2Jo48rdRJNQV+cXllDTIOvf57oI3J6zDhrUfxNCWPA
oqx0yTq7Qclv3M2pSh7P++HDLzxw5ueIZGHw2fu0OQoBCE4zTc572MZlUHupnUeeT3ijwuiAljbH
xWtq3yQUhtW9afk3l9lPOElsaOsrqm+QAfPP2d+WbFQUTWXe0GM1whFUoZ/YMt+SQ96jFCfKZy+U
/+ODnbKT8/fzobERD+FHsJ7JVfAiLSC75L9i5Y9eTaoA0v9ufMZRE4ohxyDOm4vgG0uqTSLt7F1X
q7QXfpbkQtaHRr656FQ4ZXSnrefbHUnKRkr9Ml4QbtnarSr7wM7IXjLXYfZedKeiTxWo2YMx1CKQ
O3V0IWjWE9IZG+LoyeAQeQoFR8rxLnopB9Ky5MUaM+pPGslIziRv6jv2yjidgW3ldFH8XbmuwGoa
xl5ODlQG5EAYkPEG4Dh6vF3oANxtpaRCXbHTTAif53Yxjvp9xL2FYYWUeBQoa/S8puUVgaf9muHK
5QUHaMrR4OxyHwlL+Bk7FckIMB40TeeNmabZ+ouLTrb3pt97SjXy4RFx3A5LxoTzfscbsdf4zQh0
8jRKXfCSiAPAy94JHyb/5rHyxJfNeuDNPDq96SvaWMEdG3U+3Wbu2QhdYQRIap4FpAyx0/E/zG1S
oZFSe/bSRhGcFfu1f2BoZdnsISyGlUbrdlatu28NwtIhXOKvCTk6w+yI5BXOiU3N3GSV2CeGX8mI
eRw8yh8YTKRIMnN90A5oOsiHY4A6CDCtgCmu41QL2BKhamtUurQEf0+8fFdGxTXH9n+WAVhgGzr7
4ksg/sEnWX7VG2MolpkDxooi5enKvHJqNZerHCz2CwTEbAlynkdTkslY/GC3EILuDvyHxFNTFCcB
kLf1Bp+OQlkjaRtKZk0EeZtzTaE8QHiWzvAyddiEJmFcxBdP48JPw6zcs1jVblbPZDD03zPExbTQ
VmZk5mpnkFJDP9776LHatiMfOA5Fi2BXb3/mPhrvTGsmd2DnvGLfwwBAJvQQmtQ5weM4f/+N54EV
8j9blF7ya4XL9uVu9ExEFcJZpLTYc2/udebgYEu6j0q5/PPBslrAJqR3+9apf6tRN9BDBnBockA1
OPxq/Mw2h/buCrwXhVpWyzpGl+cA9CpOmtIFzmucBgGKRxojeN1ipa7kO+5e7FOGZTrmqfBu31Qu
PtYQHH1hw7tjDaA4Sa/S6LMpcBSpEpAgTc7aPk+EdWOc0KofhqPXBYhW8+MBRlC2zJ8XVoj+gbto
MeV/ayVP3zHs48NZuRN/Pg/ELcLDcDRIzGcME45PqA1a8ChYX5KzlLfG9IWnrpThfSlQJ6+Vi0Ya
mohhRukEieMrltFhl0MU2rpn3PTAnfeUm//+UzDUdW50PmpvI+UtxYQok9+KVBPpjNpBN6ztF1kX
lUbY7fylJqtaYkKvSY3bzECDSeBD8ikWphrnYcgysl9uT2Uc55weL9I3tLmyc2m1t8fYFkfIOsbn
Aao7/87CmVy4o2r6qooygo410YLsn/1qf33X4t9xiIptE77KhaQ49fFXBkdbbtAE+oF0Yc8Rdh+v
IhoXHsOkR40wpsaaM9kWz0eP/uzDhTs79jT52LSBooQDkDzhX1SqKfU4/a6p1x3FuzcpKjG2Hplh
Is/S6wfHavECl0DPyCb8HZlCoKFb4sfF8W/HhAL5dj/KWKAurWVmCWqaRyTMArB7E7rXe9oxCVoq
3O2Gnko9po9VqVe98goLV/EeOjYbyZUwNo2q81X3dYaZ17jQ1eIryqLlk96LiOiJmXfgEtzUFB1b
wXRjZGDLFQsj44bCskIhHIswQ+8LFJi+WnD/RhTgnhRc3Tx+UcC6ssmp0EsXENw1y3XUWqkL0L1n
K6eFETfbvMJDD1odmJJrNqF+HcgvylS/w4fSdNPzrzQ8siMHfQvpdQwH1jmlYQbBCeOjXTxzL2Zf
K+FeOaDExO16T2RMJz1G5ekO4wxomOyJ5ti2oxeHutTgljd5osZpXs0uh6lCpyme7DxCSKZbO+Ev
p2uCmOBO3oKjbMn+yYGbemh1dgPOFoZTVhRG8NCwY6GLgtG7DpSZ8ERZsgQQICeqvHBz1tOumAsZ
ZcT0dl7mOWRSq8swrpOrfgaTObvaBefQJtghHfEXd3VGqw6PIlttA1W8ObTi4+Se9xWPbeCQGZJJ
p2FA8z/MkgzqIjtQJQaODhF949UgcVAURBKyxE9E0Z0tHeHkm6lUEMYM+3zNVoM/1qrSeCrQH/c0
U8eblAO28AeR4OHY82vEaI2khanEzHfCy04P4rGWhp3HYZ5vqX9YLUAUydyqLRG7gbmq4tT7MdwC
3Gm/L6JU2TUL8X/bQNiRIKN+H0dB3E6Z4z6nnYxGhOcRXKIh0wH8Ob0IbR/UetKeURR1l5XNmJCB
kUfMlbu+32VOjpVAJHha4AloFvLbhwxif617iSS3LTHaCGqnDBU1rzzZKSxuvZ60rdNbJpD7fIbq
E47q07lM0i8y8n0p3odYNPQ6VfuYAGzGrHJkiohloINNrCyzT4XQO3E8/V/MpgzySQwn9h+1Ntl3
cMdvFF9FLBH++9AQ65PogzjjkzR97oahGXObV7z983ejRmiZfdXIG9lFvXfdcMn3rADPm2JXdrDx
6ZFFffpU8UEjxl8Ipt4q/W2XOnrbD931VaMD0MyLfLmKY33754239szUbGHxqEYe5LF/yErXdrRT
FcOpncCc+YWU04+s/hkJe3+QmlYE+nAmEu2RS4w2zjsPhsDSi7e8tMQvmYZgG3YQ7TXDd2UdxBPp
1PBgekpYvkLVHx8dbegcEhqbE4agoWP4Epw9s9kqEdCjBt5Y92Z6l6vDle4AhWoGF3x4gxOsddYp
A6+Rh2saROnCT4R/8V9zTymYwtRwFn5YaBcJGA6l9mYAXt3nZOu46GWDQZrCuJeLzBbXLfRxpUkB
GxLL24rXRqVrVqdN4zKSZ51X2kslIf458vr6fIEeQG0bZfZTxat+Su6PUp9ot4ppXeRyBUC1e53e
sv45HiUszHpveXMKTqUSvS8kN3DJtiwmWkd/eiH9SCB1b2C5HpkyW7IQjpp6SX4NUpU1/wIZgc0V
0LVPWT3Cu7TYuPjFNjqIBLOnArs8rKun8EczHD/fyCBLTESippROC/rk01MtGQ4a/WuK6gw99ubp
gjgB9/qSVB59w7PGV3HN29yOjL9K6DmsGFBgB6ZXwaXKoJylc/ApHiOAm0KwEb/2r9HIueyQH9rN
B8Nb9n8k7kAV43jZjyVQMCsI/eGONXQfPyjrFUFHlUibY2jAVXpXbPQ2i8qeeVGhTIS40fP3a2rg
yTFLovXtV58oPavDdVZ7a6F01cNy/bicjZzLGF76hwF7P7yAo+MGYkubdKKN5vEywj0Q8b1aTkS3
xhVYx8LN6paTFXbTxRrZMVo19vCwqxw/2ReZnbLYX8uhHQPhLWqEJivrEr8/swecL5R7CLQjc+a7
oQrqw7pbJdDOBqeMBo6mhw/LETnm+xGPgss0FYk2jH+NH11dAaPpdpmtSHzt1+b+cKMj9EC/lVj1
3bju+NnutI5UQqD02al3bGiGSY74xfLdErtl/0xCYBFcNzolcBIFIHRnQhO2jaT6xIl4JwKazXkh
H54zRtHadV220aW2OlNw1CK5X7FnFPAV+YbjqaR2dliMlrDrKHqAXVgJEkmVA+be8iQIZMs7b29R
phV26Fk4zgNXIkzdcNwrHB1i6iZzuP1vHQBK2a54IF0bH2o+qiqEh55Cz2jDa4g8kJJJ2rcfTZ4K
J3Y3rlMgIsgctEIw04+5K1AYJ5AXUb8jlcov3/pbksrd2XBO5zHKs31KJFjeMdzBZpPZxK2lRSrj
JkpI3rHflI5wTmh7gl/dnZ0kLjIvEeYZ+Us5bNSouvHdCEteX4RP/oXkRSxGwBMx79MjcSS3MvSz
Vudj9wFWLbxPc9Fa6bL8w4c7z242Wc0U48TZqmXaatrVMkcDV6rylweMkJCMBUeEvchPViCQvCaF
2ZcipOlh/SKs5K18RbbFtfEkb0K/0Sptbz7NQ3Ir+EuEWLGIerP3McS8Rs9udK/j7q/bKvVC14w7
GSiSa9v6Kdy4DzeO1DjN71/5Jhoygk8UouJjF/lptddx4wNRGZnvUm5jn7eC/fPbnKcgLXsiz9ZI
64nkAyB8mCmQoCuzrfV2YLQzpkvH+iIpGQbdokHW/gyPVeZNBQs75Azcu6bP/4KL2QncrROQeGR2
TI+lClGS4ISoESBUB1MCM2f2P4/hqB+9GT3PRC+S4bL/yChcszRe+zSqu3d12a0RghTwZJTSkiVh
FPnGE39BQ3/d9EzSddVc0l9hKkvS3Avn+2ksr4irlehZSoLxmiJrh0VMbTbGZx68BtcpM7rgoL3k
233vkhuyLG0zsFBj2y55XKxqiFsoyAGYi3+h8pSEUZZsTYt94OBa+/m27ODffpAqlie6Nu6gjdJW
2CmBaV3jxTclrqe6dAeX6rKiHww7+plAVqXo2LYFuT4JJyqcs71rMVEbt2fe2DMlilcbt55dhlnr
1Gyw6WBPwhzEXKU2MoFnNais+d41S8/x77Ku0picd6Aq0emyKe8SteSA++M8NFsC1t2nzz/Ao+Sk
vY74PpUwklCLK5nqeMA9Ci3k53jEIDS4TZaOXolHqU5fG/Sd+sWqdHQh5SiSoEdiYkY0XbZylD1A
Lh6YYZixNP6KwhoydZMfjoh9QnihJKGryxT98rfCv0crlp7SLBIthwqfN1qnzDLtzJLkhpPOSSaE
O6pZ4WTiKC6ieywS4Ty3tjgJVfP0xWvMF/8qmtK1y72sEtnfeg5fXmh1IS6PxL6/YLBZHLiKXubR
97fFb7CeqmHMEPlF6OaQUOH/pG9k73Ac4mH3/r5sBj5+CSeBxJSycCx6B3PY485F74rFmfDgRTED
H9O/UCXaJJyyvpZU3u9bllLZwb085DcuHf7hPVCcUMVxv+yXzFnVmjhmsUySDUDfVFbn7zmTOvJp
4Rm6VduzKjZIJWc7ypzeHUy1kQXeAPd0UQwdXcpAX4D3Z5+8TlNWHraWYdNFBx+4mVdvioeC0Lpi
mNo+38UkiF6a6wR0voHi/+RO14R+c8zyxv3yd5bSRXXP7iaNErfMBr05IXVuEeZWDE2zYgLdMD+R
fHYS8EkgZyxvdyDKoFxgwwP7gBgisFVrDRC0F1UOedn6SnI8iBGi0ga1rS1ehPRBX5Z9H3E/nn7Z
6Lyhk0LBsIBWCwMK4VmXp08kluq0o6XWYzG/NAoQB6GtE6vG1pvnZeJTltTMKSQlzbZbElJ54nLa
MYXHFzzDsWx0F+GIyWqAUTu0XplWdvqIDJ62DkUmftxAb3fMYcJmmbfwLrEXK8ketiBSUnKGjqoK
nuefR+vPj6aOSy6Km3nQr76ziaNDxCbhjJfL9Le1cI7kHFIq+7fP5kWL+oX0DdX5YTk/w+/gVEVY
xGMwG7Q8ycQpaVVNzIZfoWCBJXNVM0kk/gHuc+rsoLUc0SkQcSQLP9WDAS3gBOd9/ks+7ujvuPRJ
TV2kmVsVGawkB1bzkBptPSgloPHlcGzAs7YukpJdbS7Aeyclj+bIO8bxFf2tfUL2FArAPB2wtLMT
v3o0HOFOwtKRZ1D1AI2ANz/4DID7RmqA6LsXivn3hsk3QC7ygGxbNSFsaTc+s7KoTsrywK5fRQ7O
qKdKljk5c1B1REytzFZjInvkYIO6izPhKY04wiAPaWlUNNjY8PGALYw9PaIlxva3elCGOf4mqMCP
Su8YKvOY3fZv5ESRZDjCJNBm0P2e2alWNIoqBsd4oedkfsKOC6ozjexCvKw5u1brqBTBWdKRERX/
AfNb1iCa9Son27p6dS4EFgrfgBYfSX3PV44i4pE+wJYp3+qtA+9pnyCwkyxI10qqmRdwhM/0qNNk
aO9BsdImCp3XxYQc1BxUhWsEYqKfjgyD29nONB9OdJuylsdOwMX9dYIugcN6tQwt8j7ph0+ETcgv
4PInzj55WE+Gx2HVvtF2JPHeFH+fFMUc2b3xbgXLo9zHOwduiO7o4F/LuGfpHljEf+7VInCaAa4t
9foq9ST0Yr556EUjQI/rDz2n7ZzLUei2AYX/6ex9Pb6Dcnpv/Kj5nyWDI873gWnYtq7AqLeTsWDl
DAf2pbyJjkQML3NVemcH5tYv0ER5e+v+uP67+lVgUb26uH17LC7Gt4HdD/CseRSdLYNoMyYzBUBc
mhks6Tz7WYFf5xU0YHaq+471y4Urr3mNSVdnFP3z9WLFpZrsopASpCbGVB8iv2BKAzv2DaXurbpu
vvi3B+VYmJfQF0wKtVbQlcqLUJK8fbbV0CUjXxhTlc+ik75guFubGaKDC3ydbIAUR60BtmAQAT0z
fu4VIFLWMi1YBNVoVnpr8l8wfWByJeTGYNz4NQLygNSvhrN/u7eFXuwqPc67F9qeUtt2DaTP0UT/
fI41fBCoguIekB1JxI68kbtx0+eJoTFrCyqLLme3LcWFisGj0IY+vgpwoWtpzcu8tO18MAYeRDqC
2bxGSlTf2X7zBQAA3asid+VzvUdzq71vkjrlF/C6BNMMLQGq6cUoRXuThEh/Psr4LY1D1BgSGk8X
W8INyBVAJOu/AjUETfjDmv6vfEuRKKvTvBknq2an1MmgVjiECgjDwl+KxcN4Y371E/U4oxDWqAay
whB4HU7ItZIz38Go9fRjejoOFhSjykIhTCNhzFyxrLCHtLfARPR4Ab8+srOK8YY1h+nTya2KqS5v
tBMT2YxfVjTU5RpJEbUTunTocUjbqoAPkxjFL8n4RjVh5o8SuKqsXyxJYqbqzh4KFP47rSkl+tbc
hhTetAxmBss3JcizWZ/vJ38NWmZkMo9qlWrG2tK+E2wLiQzOVOCXIMTVaWABCqx93jDbWX+kQPs8
nRKl1xDW6CcUeZhbiEUAXlF8QGdwKh7DwJwIlXnAF7gEBFAXYN9RatXs1jh055RIO6BPMNbUAit2
P3z248UD6QFkjwTArnG95ovBrRq2+WSkcS/pwtkFfJxM7k4oWmbkp88D5+889AzMsrwSDRB11qf7
h9NTOLdvE+Bqyny4Ef42N4rbgpmMmSFHwl+Mzs7gwDI+mZS5qlo9NEzx/FAI9m6xQqVrXCqrfo+k
/mptvwrw4iKiUMOgktiI53Ubg3w6j0YjogzxVem+yrp/Ps0YruYmFY9ONXy0K553cKZt5jKWjrtC
84s6H3YssOHiKnZ0Z3B4QjEp60cskRBwgWoTzoQkz4p1EvET24YYs6FT0v++0kgthE1Xio5JiZe5
ObRPpRmD3WQoPliAheJuDxFYd4PB8ElBep/QBAwh1lIBUzU0rx/V+1HOgZ3hTlZW+Rj9+Yyn6/R6
aCAef15Z9Pitndd2BynFBfJn4mltNuxVjiO6CuUSwlwI3FLjb+Hm1EkIUzvLrfnUGXT/FqS0xdqa
jSIeEiQ4nLZef6m19yq8jrmW4WCMBKMqi3lO+3n6AsanAzN/aD5xRRedvugzM5p/pncaOoINEUHW
H7gPLqwXsjU0/p9naeMg5lWPaf+SsXMwKZxNk5E3pQmgxYzjwcB3XYtIz/fDKd0r+42ocYNcB4N4
QmdfeOpKIXbDAm5JdraHttgwb6GPdVAlFm0yAE800B8iN2fcEcntfT9gaq4pOjyRbfBSKhU3yaSa
eD3fi0eYLZw7qO+XiMfRFEuh5eFW+praKkFW8P8IeaQT8eHxQiocRGPV7lkSQ+V5ZCyO+R0NA6vv
wP5sQieYqDI+O0IqAjKpPsmgAMhkMAiqYFTtjU0hymg8SMw5Eg+g9kCtLGyWpoFxb1hrz0LiL/cH
hvzRtI0DSS0S5ijqilFK4+LUUoyPY1j4W3H3Engf4XR4q6Wk7UmWVgQBNKvGTxHKqolNBoH9lgvb
M77ERcueLW8ac89lBMkogtfpz/+g2J3QIfn3nz1Zu7fJM3IWefGo+WXErE23TfpCvlcSU64RIFNv
6PHRkii5PD42bRrUmVFnXEC4pk7Ao+xq7nupprNLN0elwZ8L9P0WtvzI8ob+Socg/T10AjdTRd3b
vNM91B7NwL79egj0RfYXmdioB/tdaqRK7RvhMhPDkBcEUDHyxCZtrrUasu3OV63RHYLUQjT5JgGD
NvJl+QO+KNO7DS7YIQ15Zy2jEHBXk5/aTpIsaoWRdyW3Hi7Aj5rs1coK954aSAjbS+O05EK19ODW
bhjpUlxE8jJKMElI2N6KwJdz5yHBuKQrsfgn+ygSt9HNSQwuxsloIqEAe29itxfv2Yqg4eQeSKhu
NMh/JRf6lnXO3nULKK5hLF5SZCbLyaLC3D7J2c+JnF6i2oDHIoFE2Az2/U5r+aGne2GMPJKU24sh
4qRioNjB3nmCs9tTFaRE8Xvl9D66GQyFvxrPFibDcPFWKjEyNGPv41/6r/Paaepd/sU7GWaThqe9
gyMSZ5geqwUL7Y2mM3aaReHuj7teG3i/zNirh8246cuJkZCUzW4Iyq5tFjFe+92K3N+mdFQJdSsm
gTY9sVkHVuiogBI2NtlZa5RpCkc95KmL9EDuWlYiPUkS21EuqJMIxAjpqG+DTxmZdyGfp8EIvUhi
qDzI44J6JQRzgsCmoo6/Vae3xntzwpL8IGHXporwFqORebJFS5VIZUeLsQqpfDQLdzz3KxPgJu4a
9b2OahZ4LHE7CY2F1jAk8RsihlCgeInPmAh4zAYR0IOGyQAf9UzlQ/3DIL8nrJdLTLt/NKhmUPPE
W5/LSvhw7+h0wi8BK/nXsC7JYJcBbU1FnqqE1qO5Jci540WhRpe2ncI18eWVwR4qJ7W0gFlHT1t7
H/TPGCsWVSyW6D500ER/BAuZw04h5putfLSgcWS8AUPxTRPgnRPIS5u6orTyg8GSDEYJz+dX5RLX
HWWp3O/QcXrW1wwM1Vk+p4uCcxa7szlGH9AW3lYpSOitD+I0p7I/b1mH1DURbBpihcMe1NDwoxFJ
kGU+4THKQxbSjZ2UwfQSofsMbkHeN4VXVKRAZA0LFKm3O3ZB0Xdko7w/RQ13gijhCSUHRgY/Z+gA
JYLn5rZtD255lH3pj8WxAYbPh2mFV7TZcL5hEgTEZOgTv4/0Z23pBRJkjRQv0iHny9+0VOa2XQIA
44poG+R+3e5SS7CT4a0cViqqrLltZVP4OEJ4H3fHKMcU4cDvCC1w+kfCGJMhWhBDCXaMlivBGz5M
YNC0vnX5lRYKA5KwOXQARTx+L1cltA4Iz+3iZObNJqeo+aBreo6WfOabikh/AGS1T7viJbPFQ9f5
sKHz98M8b/t1GRMPaqSjms67/2O+e9zxfxnBCAqlL/BSS3H6J3sTVXpfABS3xp1JMvMfwnlNwmI4
QMTomEQbXtKgc2LeFcNtcfps1ZGD0NKRJ3GlBriJCSf2jsZEZkjrM/QlXDEoliEvuOdUT8SwfW5Q
DfoDflOh+e0KS5at8gnv9HoO2evjPL/H7Pe8i9baYTR8DcV9Qtoaa+77Rzgs8TuCwuJ73dAI8sCh
GC3hs2rEvjwMrrrZNI1Clc7ssBHdko3F0nn1Yk5QVZBQHspQTAL+asox/7qD7qiUIdZCpMNjYk0b
I6N1s3C1ldyffSXFTz5y99Q574wwxU/xrCfQJVmK4U58t3JxRbioXo3CWcVtnPxOZtw1ixtVmH/f
rd+OCwQ13/IBk2OAYDLipIGfbvxRKJwPc8BjDBJXMfulDyU+5W8df3jxnshOakEEMLd9rX/4JfkE
EK4nMz0zu68xKCEhRUVsQMlXcxECoE1j2p+Dd5ALMA7R50/o8r297xu5AGfPu9UqNbQrupZy5zhC
J+GLgz27ybEOMZCOlZ0W7nLz4cAA4vXsGaiJX4BiJrDcrfxWw1LGpK1NQGXiJ3beSVngT7ftFlcW
xqZlQVvpOtgfUYYOvcujaEqzap+ddNOe9FffSVpG5bGLeoVKmTtgqYXT4+LdLwXyHRu9i1koPQTW
uiz67hc1ihC25o9GEpo8aEaL0I36xIIJE05F2OFdjJNe+PmafM4omjUgEXrZQFdRkFzW4qdq36w/
4Toc+8+CLiAkKdxvCJ0E4VKXJz+jsrLw0lqDnnTIXamJFmwfQWyqQpYiv8sgW0TMVDbdWkxQJDX7
oMzt9JhrQgA7OscWPct3D/qtUl2bpwPQRRwKlFeztpeJebybTmbd/sxUpM0+ZvsOsONL3lVQ744k
mybQU+QQwMuEYRqi049BXrIXQETkeuOtzXovohIX4wrpfzLOvp3s9neo8F9LLdPYqlf5INaF9aOw
rTJnq7q4SYj0loJCKjHpHjbZwwhbFeA7syIdN158HxWuLRYJ8NZpTYsnkIhSTSeBmZqKOiQegSl/
RIjteGK9wM4yBQFvfC8g4vzOakdMtBjL+t9XGFlUFRdVZ6Wdeyw6p8bktdQo62GNv1dbebU2G5e4
amLthXk18lrRUjVDQ/TD2umSNG2+2L8Fgqd2TzUu4HCF/Gnry4cGacxj/1Iv4RzRM/v4nQqwgqFM
jr0MiXAc8pDi1uGWPZBJY6w4GC1qp1m5uAgSDbGoDwwuFdalr7QP4Ve3i4WY29LikwHeFHHn5Prf
xvT9tHN2FofBBFPVyTSKJklPwoOV7zYUhoxDXfvLUI2Hw30vFGL5EsQYHC7mrYRULWo6iCWanjGa
x4WqmUXfGf0BGHA2GlJt299krf8FZBy8j4CjHTuFTNGIeTU/rBKX7XZjGz/UJN1sRgZfSLWkUFaA
Ub4owEZ+AV9oJZqYFGLUJJJZ51miKULxpvqUfoclbB4/IWNa4j2iCXgWRdS3TernLim68p9dS+FY
aZ+XPcWUZvDmvNLR5QkzRMB5SztF2QLi9Rfc8EDnN3FOGEUnyZuQBlULxmMLDlAV77kUF77fbCEO
Cz4stSdDILEx3hRZemyu8MYJFUQCeBln2of6xYh5HrLM194oXxUydD5JVK/Swr5H4j32PtTdh96t
PkNVJ02es11nR4trZgAw0oR68QGFY0EVaYlspME7GJSK289EgFlpIe4Yx8erHryiPzsLva2QQjjV
mYTWSM6YfcnsmI5k+S4FYHDXDyLewhDilYTrAI5a/mGL1Ac+sF3IMnfRGjmOS086TjjPQBLO9ebk
GSHt8dHBd17AZGPUwygiaFzpYOMb7ZPFAGhqcF3KhZDgwd2w58AT7jNd5PS9mGZRmZ2MtYSUiCe4
WeKbGuwgA+ofr+VJN3MyLSJJc2sAwW55qb9SdCYAJrpBiBwjXSPfsfdoIqDRzcQJ8dSM58d095wq
IGRoMCclq7ESWPhuG/aDSYhNEvPDRc+QVA1PiKKZ5VWTjzTZZlgcg2aL9RgaV4FnTIzHJ2guhWYO
C5416DzIhGbAN3rzO+BIOAAWnC9IkHy+xP6ikdrLXSD2x3Epec8YH9gDc1cMgpx8hDJ8bv0+S3/T
B3rZK57y2EuiAy4/oXDd49wozXDvflSFi8Swi6/j/pDNJqJAXobZWNe77h4pPlTT3Q9+yo+Wpq2l
R8T2Tj2tQ0//HUQ6NL6Nk9zzLtIP2+Ad8rpzj32pLp3e9jtvsKNDKxX2givGjGQJ2kf6QPsM9BLD
Paz9Pu4AfnXnNG9i1YfiU2FJm3ZKhimB27xZrN1dWfsLKoL+kOMe+iwYMe/7ERVhAs74fRZ9xEby
v77caOG4I73/RVw5oStxzUqoOXEIp7f938WIr6ti0f6VbaaOWu8CpXRy3wJGJNvmE5TitabW0CBm
1X1kbDsLE4AD6ecHVW/y5KZITGO18H2bAtzFW6Mf4kAON4UJnXPiVIMV5nLDu+dWOejntNhEhw7A
Mdrr7vB1f7yTP0Vj3YjgjEGWwb7WWARr0yCqGG5nmSqpbLKNPM1BpFSbe2W2qcFDJ7Bqd3v+EfLh
Dg1jA7Ob3x8PVxSAcZoURM5YWgmk0TFLpl9TuEU+VkDb8ULZizlLHYeZLK0UDX/WOus1qQVaMFZV
otNk1uqsLwtz8E0X8KMsresFcRP824e0LHSl8rGZPZaaGSNHfzqUZ/up/ICZU25FhzrF/84Tjxcu
VOqKrZ+cmW4JUe0tjB/n/2g+geXqnqpYCUOXKeQ8f2dZ/G4k+Ifdxw+ac4RmIRd0ItmeXjSYTPPe
VGnL/krcttnecibXClVhx/PU4n05Ge2Zn0hPmEh6j53kffWA46p4Vf/o+fYIksT71E4gC10T3rcG
B4XiMwWR4ZNhQ/wCelo3GZKskXAfzf9nBQ+ydkCHroIrJIgyJDbyv7XgMGI6Is6kqgDaD8u9+hA2
1zdnx1xBjOEeNFufT3OKLSeOr+dfQog1wmuO0LnJ0BFz7Xyop3YVj1ylwT++Qa5N419oofDneiGs
9fubyCh5PzFxbyUVPGfM7qWPg4OgTpaoMQUNIXn9Sk4l+1q9W5RVJJOmEJBjJZdTyP4tKJ7/ZGUj
qY/nGO5HqflMHeQdrSBETWPZpASi9pLUrX/YM68TWaAv7ld5bqpjVNpOSyEMyWOu/oA2mwkFAvb+
1KkTa3wWs4rOB79qoTzfki9g2cLeYENggYvJwY1TuhQPodEBnPTmMIDosskK2IdFCCFoswF5cYLY
aySkRGZ4Y9dZxUbTcTdMjF15GRvR6s3sjSHf3tZL9X5Ck5WtxB669lLZCYspADgpoedhxgCy4jeH
W1xQwVUJ9DFjxJvhvMFZ3oBW0k4y51UCROAqJSdelEiukHpodBkCf7StGkfjYce3MVe8zq7bBXqR
sOjAeOe3vq6OZUg3ufj6GJnxIVeWd06zOpFZ8QJB1U7e3VTpYs0Egd8KBA+UiVA8gAyfo1pDqwOP
RZV18P34IJpe8pc/QO2aMl11H0AYrKRMyoTID9rqsBbtjPbCVRGVdzxAcqsgkDraoOrYCQZutNOM
Nek953jrYfJ07yzB/jNbTOerpUjAM7Mwat1kbpVlugBrrwi2Ypt1Tp3ZV1tTayE+1e6o4FHKdf/o
zV4bNmU8TJb1zzw9HLRaWu2x/fwcQXVNA7D6CR6/A1r1ZQt787VXDgrV8xHbcyLgqc4PQ/Hcksvh
dFv+XtAx5oDpOYMNkEDBzHjiJsQcYuXb3xCWJU2OFcROXEkU3FPN7tkjb0b+oJ/gCUTYp0YM0Rt+
3M0S5yBErp+zRWsFwXrTTKQLpeDAOSI15/VxKYFN1a2vSbwUk4sMidjAedBb+jtVgTjX6M9q4BnD
OAgum2UN0fa5k1z7XER5OMMW/xw/z1os31NylE3e40JoRhUjkFUtsOZcveiwdVb5VW4TFkadAxGh
vmz6AitizI/jfFjfpwHXH0OGjwTMyVnieWX0OwzPGRBXhwoCcmXMnrFjszQDZ/iPpB4wKC2yDZU2
n2EaPdDNUiciZkm1pmnLpxrbxx/6oQ/M9sXdfwbNxPXwAYAd4vboLdZfnb73+OAxCU8uJsSKl/1B
Ecni8Od2ABVaSHGKq+aJaZ7PyW4lVM/+mFKOs5c4xRKgCadCgd21hx7S7li9q5JmdbNQTNABt8zV
pGjOFgvfT5/JVw0mH2cixy7ifSByJ2a4FcWs7b2QQCCc1nfi8v/QPOS5OWuZEhzpYEc8pbYk39IL
+Ty2GGdy6pHOKV2JHrspq+Cx/2pfX9glY+Wcum6nxMsAnDIv1a/OM+syrvIEx3in9B24Cye8Fxqx
Mp3K9c8WXbD6+y2aHZt3NxDU0ST6tZR0HqIChjVrOP8m+SkdOz1jD2OTXxJ7P2sOTukK7tP4L1N7
C7+iZICBNEWmFIhUXnI+dJVXTmnWfi5sCCGzmp0tNq4TbyHZ4Ll64yZtE/ylmEjlpfSj9GBpYkgM
HnKHI5iJBcYB+KeJ1EWrjDbgv2EsHh4ep1i+8IjqhUVu8nb5g5f6afH/xFeOQQ+MTXSOVv859om5
GCGhHbrL32u8BqFXK5YtWt6DaH4M8mIwhVvXvf9/y4IE6Zqu6ADW6Wn0Hkz/9oIjx++QMja4cZJJ
zamv9CsQLS+Ot6T0TeYXPId4qeK9/OH7TMgdKK6S5SPnbX6r9zKRGKgC6Iln94L2mdE1eiZqraxJ
h+BWtC4Qje9pn0F8WFXIxexrLaAtF0CNiwd8pRAmtM0hlJy/08olTP6AVh6GYRQVWm2n+3g0bKvp
m8rbsARARmIvcZARFWzQ8qZy1pohW9v4s2RTeWJabFdzxHlpU50ycDjzV0a6P7z08hxukpjmBOV7
DTAxVOxi+vVBkImQf//hsZXvoeNmVTjAFoVrfaVjeXe7o46XqcjSL4y3U5UNSbFmZRKL9Fqofal5
XCDb22wUMsaW60Vdqpa91ITjHSN0U0AG2H6oSS1wUjA8zae4yOEB6cfnEb6SZyp7UrwBhtb7ejbU
xqeFsQmZfcp5lbwbVnpApqn5bPkhj4rXghFhJVdLnGlYy0ZY3O+f+Rb/Ras7hD9P31HcVHN02+HJ
RNoZ/Xcx6zuZqUCj7oAKxoCv1Xo6zCymB3cEdtTtwbviHGK4bth+1FJDsiB1pFBRuHcgCpsGbtON
n554hk4GWWlb1RmFWNKPz4H/1r+VErPT9/uHW9eToeZ+kbhXI2vxBk/cXw8cOus5yWHg/DQSOb90
Zj8kbK2j94/hsGVlW5Eo/iLOXhlewlbU/qPhTcIcpS/Ge65NmJiy8WEX5BC4tnvF/b/h9qlmEDmm
9VWRVAEXOjJQeM6MjqAjysimxVe2ByfTf8Ll2o1JmK2kDF0Et3Kxh47p/ZtGNa0/wHLjwka3EJoa
liZxRzUldwCiGcN9oqEn1TVGyt86mBJHi3eN/MvcmHZohjx14NwtcxNVDzLLiesEJcKhJISnGMZV
9w9+AJdfyNe1ScAcZWZZzNhNbU9AKwnLP/SgoS4S1A755kOXe9MUqm7EhAU1F0YjgnZygqMb1Nit
dG9EBnq19aTvH5qVSQgVaqOxM7ygWrd4Qzx8k1bYZ2yrfFZLAzdd1OPgzUMKzAkgs12mt79YbmLd
sV4ze0lDGsN7snexGywqz5I/CYp7lUCSlKfY0Ke3xxh2GinSuEzYY+TfpnEuRDtSdaceZYxpEgYE
JyVdnYwRIV301jT3UFgSNVZWEA0WiZ79hA3qiADxdfl/mYNHreAWblyr48d6GxxGs0OHLh83BMt4
WrvGd9xFRkRhhHLaz/pwBThlXQKI8iTXJr1LJwNCibuqZEvvFs4ibiSqFhnwaSMjCZu6K6T2WsEs
8FLFBUlI1lQtTbrVb/6AYkV8/YW624+ohyLNzVc7+S4misnAZATq4e5HOOWgSbG3OD2gCghk6pL1
THxT658rg33QJ4qIwaVScCRvAvcObYuaJKBPxpc3FtXitFV+sotBUVrLSe8ggknHIyylutnvYqxb
K5dJlyP1OK3zTfFVGM/6BAyRVkjgwbB478Qp7FVIrHl75akz1wRziJgeDpE7sOQJQQvXynBUGPTG
iCEo3tsqlkV+rHxy+4EJKd0Jt08We9OZOFFdk2n/dk4jTXI6k4ZRrvCSyNNh2KkFZamfjKGFX/a7
REzpOBTNx4vEffxOQa74nllCYzoyZJd+kR8MT1s7FwTgpvgr0//SKW3qr/RaTrasu5CnIXVqdy9h
56fSdyPvZA5Vd0X9XwD1v47I3NolOJL0rnn+V29L5/Guit64n0OZnpiAGcaIvElWTkrjVzQS/+b+
1j98VB6/ulPZOgLTbQR0ykbJ9ZRbLjhZZlY6NmNeL4nE77tmieQeuMle0VISdfXxyOHkTQ3raQcr
J0vI1X2qJrsJxodpA7/IpmEVhWMjhaGy5l005nAr91U7bmP+bfCg2x0u+msQfr9u5AecBYRig2N+
xy512LTs23Qv7yA4JnYxOunMPTg5mNyAU7KeJ5KuzlZLlThuCuScXJH1VcH+0YcJ3G/hOLD4YNnX
vRnTGyXPhmxEVr9SUXeI5v4m3lUb9RCl+0v96WT6U37ztwzdACDBRW5JPtFvoBxY2y0khoIVJ8NA
2ajAaBu9mtFQJyIcgyRz0oNO/4gT1101HyXaZtxf+6Rw9o6aNOnDHWEO3TqabTQ52bPW79fT9gu7
ETgjak0Fxgc+BXwEyzvJ0IBei4Q+PmzU2LW5wNABZHBbh7dMH28z4p9wx5UCSLD+2oowYVl+wcEX
4L7uN1BqwHDDGvs0G1sr0kVnwG+VIU+jjaAMPq/CVHMg57WMi94QaLONxJO4UaapTxLBtrwLf2y1
DZYynSHElqz6ymyFMfq8Q3D2rFlwaE486vsxwpuSyIr2zoLEvkSlyOQpKFPQt2FMTAJAoF7Ji9zv
Rl4ijROS27ptjlcU4rdZwbENIDW6zlYHZJ/kjnHAGHJPnmIlX2duvKYHeLVJNPyu4uKHekqC+Jxq
V5EMxA2huXTEn/9cm+gM2QLHveFhBR4eX/lNwMa05Fo3dSN4RMIzD7fZhLs4CizLsLLgA5T3TTiN
2csh5AldeIJCCvOyDC4X1l0laDymA+j8A2zYcQqcCuBCK4qfFYhlAogbfRfL6+yBGYYAyL/JxKan
p6twlDHk/KDWJPbFdOvNygU/rGI+UtqlYfxea3L1XB3DCzsQxBYoxSiU7/RFVwhZFSNu7Vs5LGXd
7rUCU4fJrH1/ZZhLBHs6Ll8dPTaB71IcqEfXT7H44+t1KTuxYel4S0k/A4Nnvxz2Vh9noMZ9ii5P
crd8eMpCDSZo/SLvGBLLUcdn9PjwlYx3tswuMPVTand0/+WKamsKLyp/Ky2OASwjvnMRb7YBq9L5
OzisC3h5BjxrSFCZFIaHkgTLeVrW8fw8hxFpb1Ud1His9t5RNQwBAXdGSWImY2BjwQPG2aMTlAFO
Vk0Qo5Rh5JU7wPgA7ON3k45A3TvOUlCYWRXABukIFuwdOrUj4BV4f0w5zfkfAfDlFRFUSy163RQr
/LFG6P7kMZtuIWlAn9xfYFDLvnQeENiIu65ZO05wU7vtNzd63JU3oV3IFKA2Y2iapEGD0NR+B27t
5uHMrW0Pwuevu41dmcz/v3YCHxcgslBKP3vgfDJKZ8S9UUd2hZ0CGrqIUeib0bSOOcL0fdYEhnQm
Lc/CV8r38Lm4+vtSZzCxJNcU5FzjRl5BvlPHXarGOgwYCTSES0ON/fnfqIh/32gFHMjEJHTmQRoI
g1gx5582F/3zBUrrL5iaeq2BR2A9rppzlR6qHZXLaBxfadbYoIegXQ92xtjq0NhxgQlfrYcNOtmR
0a3hJLtcXfAvxqg5/y+4RjC69RqiT7YiHYZwECASVF9U1BAqbDNKnwWU0rzrcsdHPBWYUmprgkpV
KKnUY7BZeV4p0Yk3riQHMLT95HoaD9tIyKhcEe4wHCAY8Ur5Nya+MTQOG9klxnsfSaXN15pGTZi6
/aThpAKiDPSDawoEusIIr/Q0ZbZ/Flcnoj+Atyp3/MS4hrT6VLGMk1AYNZFUb4ThLBXI92n1U8yR
66ZXEsbj6Cx37UJUQSHoTgZlVfrwsaSP01FLWAA09mOzOXI+Ij3uie6+79rv9Y90I4lfW9cqSqx1
9cYqdLD8HFBwrtxxiJxR6UkySHjhT8M1j2jLvPT4jgCgI2kxNNcrRzaji+IVY1RPq5YWeJKCNqud
diD+cb3eMqeOziJ3XmE2q2XNTzOylvVbwf6ky29Cz1sdVIOvqmobEsdu9vOob91ggPAd/wRk6btf
+z5yhEc7Rk8yPMWTeGuU3xw8Nm9iiC1yPVU4Q7OGJn33N88tLElgeU9r1vS0lBd9Uzt/VlN9IqBJ
Jrft+w91ciudVNQPaxdAXhkpEyNrdI/uYjtUk7VKDfVF36Nbx+odqZIpl9VB+sHLOGK6lFw0Q3GQ
/ekZvw6bEaEnrnJcZOZod888LCmKpZuZf4N5xv66n5vxMqh5qZMLxR/d5Aj8pYy9IAi6BhXQ3cZY
K+DsDnmUTyShKDYeS7iN+W/N5LIEGJqYLnzGXtu+hFIJvPpEfQpiAwJgkqD9Hdl2nN5LFFJIpME0
BWGxAcnuYGxEvd5iMs07J1+x7dDzYUlwHscdTZ8vX1k8FaGxWRrhGzxudU067vVjumOT86Mga7Ss
2gtWmk3nhju8w/oHhf+Sc7VUxER5QcHjedRoC/kwEsXr8iSdJ5pZc5EJIFdF8qtZIMWkhD3LjZQ1
kkMqPcDBZqmwOBvXin7T6MjupGHn9v8ZtYIGIKj9LCowrIGw24sQnrd3PmpBzvyYZhoYC5lBnGtc
zXYeSn2uvnjgPRAzRYNdPO76KEudmPU7fY/Jb3ZXxX806KkNfIqjNDVpkSDD2UVHsBTxajxP3GmD
nr0+eqXQBKetIxyfZPbjyJxF01wlJYyjv/jLzW++zsJUdT882TvcoreoP4fjTVb6Noei4jJ4QVTz
TtfiUvXOv9GvuVF4fdnUY9/fnbzPBSRQEdpNIhsco6+HeULW6Ux32VoWZb9Ggx/en2rbJFAf+7Jo
CFMmRJSYv5t3U7eK0gAsXgIbxG+XWBrjaOPQK5XhosdXyF4vhKIrJFoIYHjdjG6biU8rZC2ZphUU
syKFrgq589Ul+DqVZ3Yz5ZZ+nkM5J9v9UPB53t6X7KgpFDxMJ0ISY2HJ0yZ32FjNsDzW4UyB72VB
Q3gQ8vLAYcFzvwSGtudnxnRmoulQ6BaaGhYDJPMIwHJDEBwV3w+ULdXnzkKy/Ax6J/hTcoUT3gmq
AD1470+TLIBVh5IeC6OgLUlmc68wNVTZmuSGVNnuvv09XHFwvmwAw5nfqJWKoh1wNtsDF8gWOODS
GzBJoCCiaO0hZfndK5oM651Lrj9qoFsOajBqOdLbEQ0hhqSAkSa9JGMd8G9L3MCLA+0u26vvfqmw
YPXpeQEOivFPVXBZpjHM7ocvyg68p6e0egAVW6wiS9TpnwbNe5Z7qgHrPvkLSO09bPogMIbPqPTs
plBQgIFbCv5h6pAnBMLWpiwYSpgVAEB1GPExAICR/CBDOqZDuUaVhKvznYDIIoX+Y5VnSeAxe5j+
mGOFWGTNMl1iEPGREgoz59YUiWlSP+nnY03+nKfQbK9mqFMP6EPfBRJ0obZwJyoeWEHGqIafHtga
PaX9SOAgsW0AlCoftQyhs4arybRCMRj9s2XjImyorC7/BIWAQCXazKHYo4j+dNs3ae/HWRWUXT86
8Qv8C4pzeL0cFs0E5ckXQH+ncQCGdBJ8DIhCRRX8h4z9bd9TQ5M0XLGQ6wvKztttLBcAC3AA4RpN
z+YW4pSKfMOSXRNiRt9a8Ma0JQUJsMOc9NhuElD9CQnfe42EDcDYHzdjAbR4Em1OHM6rJUXnxya4
sl4stoxF/OTpiDcF9HMXYryRCZXtpoeXIgR1NaKpiScTw2DLTP8WxvtgLnk2id8+4ubZBq3WXHIM
9jiG/yPhiQ5iYKtUvnhLQhSWZoqAT8UjYED7yvKUJi5hKrdXWbrCEz5Y16IcHkJwK3YhphXMC3at
FTZ1u9X4cnLD2XLPdQXixG1ej8XItqHHoFnWBfCt9nHpsIXY5zM2n28dk5fef2zcmoO0w4HxVbhD
+xP22flx8+mXCgaCHgODbvAOSVrC2gFsTomAO3eidkXWyjcdRxyYuF3V1zzKZVTFBkucwVep7q4y
aajZMz2DgCAPP3F8AWP6jh0i4fKsKy/B8BHds6JzKzZzvUe1v/H4cRrR9cMxr8yZQzJw71MMJpq2
emZ2d9poDIZ02No/s00S5j8x8YfsifU2hZO/UemX07alOqcbPZj6wT7pGTdLsc/rUdy1RvuaqfzN
P60AuNPU/Pf8KaGFcPPAIyueXI7gyijZk9qVJbjbnbyG7nz9RY2s87VeWaE+7i1kTVLnRTC6nNss
bkRw+3aj6fyIWkfMoU1igrSgSylfDyxVkV45p/mTVfXhGX7IArRM4DWP96RMZbnfLNdDnPlsDjpd
mDoFlwC6DzgG1cezwkVsMPwwPmtsd7u0a3CvF6jEb7opTP8J9d2/6adf8ulfko77zCkym3LsZESo
/tTTRW3vlq0JoC7ziNeVAUT9upypFsyOEDzZRWHzmJcqbWW+wfodYUgIFjB1qKD+ukF2DacVYvD0
TWI2iBVwtNVDwLTNZIPt7VX4YQNNS2tCJ1JSOdbwPsrzOcXuI1m9EkW5kb5bvcvAQ/hFoedChg/a
rriFMuIAJlNSJMjk2SQhA9WSuSuIKptZleHbAa/0NKuURiwM2wqllHtPshHnH4/3eYlNhLEnD8sS
xM7D0UcayA+9f9vLBV/U+PJxiBnADdOjk6v9m+wJDWbhmGyQI2k2r5Qhuley0fsmQBk/LurvsXhY
eM4jdgoNKAsYrHNfT4mwT6hTQn875lTYgIbt52V5sMB8ohec+6bVhlYA3qEk6Z71jPn2wYy1aAGW
uV2AFJlx4Yn5tlGWxGhG8vydymiJ2j1+T83wuaCjm/XUeAFodNfnLr1giTu5ehEkpbLDgmP8OWn+
3E/MBwWcoM2qfcUS6hjrt3JPV5rKqy4qoJ9nDt/oFtwLMrSINhnIpyE3RQP8YS7GH/QXrGlhou1w
srs/RpAwqaiU+R4GMGNx/L5izKoVDhumeYKa6vmCnjbixfCmyTAUHhtGHoqR0F1YPgjEk+sVjutB
QL451YXhQvtd31iblkawe3fb+e5wQk1bfBUJ6Fz8JfAHId8wvIpmzZCDyUue3ZKQZtm4vn2kIss4
kgl7m9wZPveYvnnE42afzjFImjPzt4TxPXM07plxXPYVDA9gO/ZOtg/yNeQbqCht7ApJzGuOK5cU
0QHXALXLmmwO1/i8eB+mA9RDVPBIeyyzdLssRPVdspHHvQ+ZMAwWXrXAdgFsuep3ee1yUnDfRrzo
UnyHxZdVdY3lz98zfMRnb04iePyoSBqwFLDj1tLhFydN02pwksR34rHPx3oE0S4aedV/27NrBDJb
rwi3cHgS2R8m1pfXGUqEr/fEvnKD3m9Xc9x0dOPZsPO/Jf4ROPB9zgmNsBvyoKM1b2S7nO5uYHmV
HveDmpis5zNTMrHjfwsBkJgjMfh9QQ4QWdM+VA0suU1Vb3AUdVo30FWxsgXzGKz2PEtBtyQ+nN6b
h2ZfpUc/nvBs+xqIQAkSxls4M7ZIH3q0JcWgNa0YYNn6L5/zD7bSOr4fyY7I0yFPeQSd5oKNZibd
DwAzDNB343ec+060vOMgY6XD2KDdlor99H3d+exd56vRFN6ybmepE/uqMuM6MyMmPuRxBlycC05j
/liFLNgVNo9dXbnOw3vh/ic/JO4p83NCmRr18+JzFYm/cOezNph5ac6gUus9d+KeMLroMkNIMu7M
6tmOcooxSyTV6QMR5qYaSm6dU4xunAknua42ciX01FextFnKEpk67LiARKE9kOcNUMUlY5fyICmA
VciR2rWfPoSVMP39rTKQlfwVMj9M5L9qo8NN94ClImrZV7NLa0C+U4dudY5nLbFI/S8tGmJ/SLbb
7s00j1UbpDHX/b/PTEFytwoLodhzPF0s7cx8gQbyq9XJNy+gqTBbNfQfqvcx2tRaTiTOL6bJCUX+
95zRvTf7j7wtlpCz1UYhW0faw1xUkTOttiSd2A3hG9QXptKtmzlOmXHCIx7jdeTI7MmzfA0txZ5Z
yoMlplVnwVIi48t0XNjuehMt0WD24YauKJegJsssk8FvwpAnvUXemu+w3DHTUjbKkcNovGMi8jX8
3NN5S9J421ayMHvKRkfL1ftGFXMkrx+5dq2Bv9k9z3/FI3SExFoQpM+p0+LiPNUSYABtU4RnCF4f
hoBMIIIbRcHdrmKTwG4zfvDUZd/1AJkgwCD5uTINN2M4HFXrFu7q9gpaJWv/Q7TrihqwGl3KypYM
tWWcJTtP8EySVOQ9Fdlvi86bgdXngLDXFOco5x7Et7twUnkY5PTJ6w+5vR4y8ncXdhzHchvwXWaf
Bhqmdr+1K8XwYIt+EMS2NehBcP0L9bhPF4PYELOHLFcM7fQ2mCLfsuKbENE8vAi0QbpFP83kudSL
vwWE0ijeN0ghYGhkVFMIjoJPEYhTgC43IZ82rvr9F0PD1TtIDHbrrl2cp8el5G/V1aXqZzHmEHaV
Z8fGyXiHoqZYtWH6bZ099RoEMKx5gamiEZHC20LFvt1XQsSxTEFjmHRj6E8p4ujjizg4N+d5NEsW
C8SXYbjfIccOjQlGQeeIRA12oId+KkYGlKqJFFMRC01VtDUjGs9LSECWDUjYwvPr148cJV1QE+Th
nSK/O2AZAvDNIfwUcwHpkXDR3JX71Jp6J6bAGERqhNcnUIAw1JG0A4aFAn9JFF2FTRm91iu/BH0L
chlAsd2rC19HH2SQiKHU7kYORUrPIasnffKsk/aZNTjGtpyQEzB0q0HyWbf1Ld7u2oIGeJ8Qc5p5
vN7w6vL2lo/CXgl5H0rvyi/p5sN5yWqzH0dfZrWaVQ7ZBLV336K72wZ9jVjJ+WvXcXx0NQeVJmn5
2+y/W12khlBp1gOerNa4+/r7VnUh4UgWYj1+TYbMwZL4omtNK9qNm+FLYG2epJpWolHAIdeOpfbd
zIsrq+ZqC5GVncSMdDUAISn+D1Po7zVAJMgHlPqUTFDtxNOtCFOHc+LxpidYW2R+wAMWzBJQjql4
gfvqr6kVtNGqORIrHKb+zzpRVYmyx5s7CerY8CTDweOSjwUQXXvTF/ni7HfpN4cgsDoIB5sNxips
YiRwrtmlJ41kW+YQ3nxxM9FFlWHiPnPRG5feBxkQP3K8ECdZ/oOGXoLR9I6GNCq/OKsY1L8bbplc
yAV0Gxg8iyqCLJ+7nelyN6WkBkV6axer41l33Zq+iy4GkpghNsy477/UZ1fRZyZZ+BwHq+Oau+ob
pOQXookbBHUImQqR6PdMDcvbDtzIlEW1fVEIsO/gURgWRl1sWXHn06lISNh57AgkqPR0VHGm5Xih
QWm/EEkHvOkeqUCiis6JiJCZQbi7W+57LwS3S/U0cT4OlC7L0C521G+Anq6S/nuVyYvMkKnU6Ppw
UmaUU/ejOxAPmx2bM+H2m+i5BllqYQS8dwcuEu2bdf8tjsv2w2GqCdHV7xiJvjwsDuws082I7s1Z
nHUoFoRI2sHquNHZtpwhz0f6Lds4/ZoMkUS/BFzCir7yupl5U9A8DUheodWh5Hi8GPo/m4jfmwyc
oIyHTW8NjP0NTm6B1yGNx0ncUJOR5q09BTdJXfkMYSvbWUj1aMHIt6CL9z0fSoa9+aDk9ASyyajK
7Ie9QIGa1BeqUt5/VasmoK6yUIfds4hCA5FjkNd/WiGG4982rZj+294ja+7QVHx5omqUqB3Huha1
NYpqYLUz9frHZ+sRDFqXI0zGXLrAnQ8cSLfOo4ZFInhhUxhUb22St3Yh35gfI/m+9GEe24vo0YB1
R85e3ZUlvNXrUKD69ffrbBqJ4X4o/R+BBTHnbu6es6uV3wVrqkvz0d7mJAKyTnLD9SjsqJy1d6OJ
4gmyKi2Np18zgin78QM/NAv/RHgSVafbS/44lvYcEE0v58/EuSfpLjhTbsckuzkWdnup4YFBhvzS
lJk7rcN18DQINHapQTjplX682r4PtVTcaAdeiJ5TCdJMfOEWDOwnRD8ChMCnL43MqwzCzWJodQBR
UDUTnf6L2FlvCCvk9WifvbAdzySHNXijZ06lV9eaSmuXszmLbcYou/TM2Im+4ovW98/IfOE0b+CV
aLWlV/+3kfwSpWrXqMG8oAB0D88uKL/L2FnaRiTspQeTG1YtKPSyiHHB8w0VoUU9pW0bh5gpaZ2C
+s10/e+r6RLxCwRjnFGd2zUuxP1zDuZkHuJlk/FLVKK7P4lVe3hsyW7Xhp6qKU+be9b72BvEsaLZ
cuM1acgN3hFg9WEw9jsyN4YPyNakYdaKyiGrDe/txXOkzGg8BoXLjcHE2WlRKlOudcFqeFBemucW
wXxELvtZuZmVLmP0MSO33ySzrPKenR88VT1ArWHwLlgP+xY6NKm4/AeyWhxDAwNEZ2eF6hip7udl
y+DiOMpmtTnKGhaEwqWKeVwmNbN2Ja+UblVeHBxgPnJ3bfah7VS+CntXNDAZXJ0DzJksioWBCySB
URGYcyw0PybX1Xw6U1ezXSccxqWdtvbrmFgE0GQHWCr+8/Zzkvoug6RcHwbZzcHhNhxWj5udAtEf
r64aZAMhtLFiCd+v5gQx6RRtLUm2/zjv5GtUzXxyOj1lDx0czCeCACz4TzULE/uAm7ifm0b+9m/L
P7YqzRE3SC3xyu1NVL50cC9W9/1egQNyej3MKfQfZdY5mCT6dDuWf/tQQuLKL0liQRJymSG55MsU
6Tu8VOy+Hwn1OU6X0fQcgEp1ik9LE/7ZBXcJ2xrgReoZPsqgMglAWKDZmRWWN+58A7yZ81gMCCxX
KWJ9HhGE5YEbRhySsbIbs/X+FIiAp9K/D1jDIoWmrGYyqETTnCiQKp9yC75aLysKLCXGGPvTyMwT
c+tP6IO3zEB7XpWskttxQ111v3hzraqDapoAn3P4uZuow1UCSEupatdhrrQzRaQK5oxYPu3oza4l
ZK4kkqqhHQGJa2gSMXmgouVCPJUntqcT/lyn3jUNFsiP3Nl0r/gyaWWQKjRTBD9LxNTQvBtWMbbm
otFFZ/NdBdQz3KnuZyZ7kYxOaSy7nvILVy/d/0XymjV/z846lEO49l0uHyUh+BjjduM+lM603Esk
6Llz5SfEOMcU8I4umfFO4nm2cGanfJXLh5yl6LZmuP2Rfs+CRAoYt2xtLMHSgYIkOL+w/2YiqRmM
aOjs4Uxn2SJ+v1zv+JvsCZRunhhGBGcYa7MH/dRQm/r7i0ifEa7uvmDZu6HzwnHKKaG4CpM1PrLD
qXycDMaZb9G20x4mZCQQ4HlO7nM4lFEhQkWE8AqkbrmL9yb3xp094Kt5YHVAOMWLfgnDx1xH/OT6
QVIvoySWBn3QZMxOXhq2yI9j0TTZQA7+RElAYg9NVJ9CW3qETV5s2qaG/9+lq+s/XqMAlX9OaD2+
jK36TdAfKUUKRtDaXiNUEIwB45tBjPiov0mtGuN5t1p1g+2fYvHbWbf9EaEif8MZ9S3i+9i5kAAQ
fCBN0lyNU4Q4ses8ROVBm8eO4TCfW7Qh8rDrWToMNXZN0h2+RqgZQ1fsp9oo1Ud/R/1Ath3R1oEl
0qns7Ji7L5jyR1DbOHR7/LidS6+hPjKYUOFCkz/c7VymvN4cf8+ful8WPfY6i6lvCY4DIvqNXDVY
gBoUpMT97XHwYcFHTdVzC5btfYaFY2hx3CmFAMv1SNmjpWcMQnDsu0rKXsr4l5UCS1Ib8FFeQ/bd
9qQOGt2o1kRqIcRdKwjKmVYS/MrwaRvEWB1CqOUVwPYRx+LYh+F8NVYo1bB2SmzDR7K7ubkn1Lle
e59MFH8brX9HZfWB6+6Bst+jTg+Ym5weIPzQTFuxu9U2gcM9yhmTEYZt8T/CNOzqUM8+T5Th4f5p
IgAFhgY0mlbzhALSKns7f0dvXQJNQd15Co9tW1uMOmBZ8s4psnWydvpe7B3/7tCqwT2Rt6DYMfFT
3DyE4gkqkaaYPXhlukB8leGnuIlaoKMZkk1/9fic4MEbQOcTcqyfx5wRcWBcbjQmSQoSgOFRX+17
Oc/lukUQxyTYXBEs0KySkL9RuuE6Kj8GQ2qPJn/khtxDhhSoCriKmBbykL1+SeT00nehD/kZtTZJ
0URAtrYW+pycmW5lOhQHIvdCapzwa3pZDHvZkrmXr3HuB3xxrf1wDf1wM5i5PLx9gBzmMfkJwxvz
68F6g7MFLlt3qYSsdsNpIqLjDzoJEoWZT0XdFzlCbcxSLJtnxLutAWyKZKURJoeoLJmHCF+oPNlf
18acfyraAowiWhSRptlG5CF9pkSQrfguuDkT33nRdMsKat1NRAM26hmBk5hyR1KX6UD1Tw38Aq65
+P7/gOJQzyUAozcsNSKIFRFAhdoOTPNvcOqWYeLhF5+1Rh8oAi9xPYUeC7Z13jRzAyWK5vr//TbV
28uNmPObFUYFZmI3VsegG/CUvheCUISU6I74WLTm3bs4XzhH81Rthj+vHaeKnQJQVAJls7ETqIMi
XwfNKUBKCENWE/oDnYNwXvUmtkRi8CAPHU4kFb1DQ0g+pxDPs3lEv6DNPG1dIEcfc6R4WNeq+lVD
0WOE1N7DubTe5PA7R9fDYC0R4iblVwCEvYjFyVLmKzRZflZgm68+B1SB+kxPoTgkcYG+8pf0QKwz
irmk8G2Rk0q4EIr9+w5rGaMcJwcfXmTb53SYcmiSiZ5um0eJSO8oo1rSYjdiLFKjJvEUuIQBE+LK
5PJpKBE+H6q5auJs8v/3QcDV5oJcaSa5q55DZavTZLOyiBPd5Tls6xt5koOPggKEVujV3bedCOQe
lVtXryXSVcbRkjSZkZ0xBf8yjXfHU4CfDW/mCa8r0inwzBC1kx7usX7axv701ZunmC69visY2P4t
8OF52KqUg6DqMtqau/hS5jCFHeXw56XXzB8yhCIPC0unzf9wpmUXnm83F6ETaUTrDE8fhmAOfMCD
057CmitEsWjI5yGZA5wFmV14knhxLYXcpgDtEECdG10FOQwl+0Od5IY8P+vTGahQxsqDmPv380xH
qUV1IwkVcBqzjxiTPWudWacWe79/v7pL5Oviz8yTT8LWuln6rZzLMbWBPWAH7df8lvUEcmxT3VMk
SvY86uVxZ8MYc1PNlUU6OgdV03y6yDdb3Km+XrFHMbx4bR6A5QwDiTtPcuhbFR0ZsmMTRQ/czejc
EFRBvS5Fs2slXHJAdf1LoozWJWl7azVusCAEUlAmuNTaiKqP79q9QlBy/zDl1FL9qFLzt6UOJRxD
0u7KfCMYpbiitleKUzfOIefFLSSlib9+x11g4GWiRuvyc8UFyN0VZrtCyBxoczvjHH9UlEFlh2LG
H253Jo2yCov6YJ32p5A+teeKDdw21s9ajQi1+1XjoMpvTvtc8Z5AT8ZuJmBtId9uPVb0ubSP9MrC
B12QSw+wt4NFUrKH3Ns5KI2m8T825Lr3xv/nBC4qLbm9whOgqn+wXYxEzAh1aENO8SCtjb3Mv7nw
V+nW9p0zeAnfykg0cy/zcaT5iU5rnVtBMwLgsHPjpf95mJomUJc6I0uq4CAEvawybTCbqO+vga2s
022YFsJtpZlnwoZygphGkNPrAS37RF75NUe4eqb/xbVep5RvqSuXVbL4tENpZAnkkJxaWykaT2i8
mYa9WTRY6o9gdUd2/x5nUrc6rPziPw0bIcAzuYkBl5O798qCWR8zKjKIWJOgpo8ounUnbq/9kq8C
Pn6QSEjoO5VFkllWc7YH2ym6WSMsuCU5wIBezlwq69dCyOzEz1kSYkQ3W6245KzxedcVdtqkA+Be
phtgADLRhwsyMpabphJahdoG9B7Q2C9YxGG0xxXU7s9SHF+0ESmMD6uMVQN2suBUEZaSSDyDzXjH
oHoitXwTVCevyl592s8geGKPx+ihhUU8uBw/BP+pQodmG4kvw1UMFnrHwEtFmIgPFCaQaDI7D2mM
5zOMgTgTvopjVGjEN2TkQZXwpJAMcaddLm6O3Nrl+GdcbieTNMnY7xEKbj4yAsm4eia79o1CUFiK
RiTvinhom8RCjy8k1At0Hb2utEiFrZw3kx8XMThxsSma0+2ctcFtCJq+hsYi3nChldz/K8X5uMoJ
wb92wu2kfNaMrtODCr/A1LzP1ICE7i7f+wfpYIZSMyEjgGq4a6+RHCrQey36gbq15DpGj3HzpYMk
2i58D9vhuoc+eZkydlGV5tBlHj1UtLvgkbqpzRSaAfsaVcCnvAF05NIu0sTfjM11v3gJP4HB0QN8
bie0y0UvqGtQbgccNGVUFqa8fAKuRQXW0Yx5E+SvuH8XzVf1xd7hFg6tzGDwAKc2iGPqXlrMoHQk
VP52Mbd46Cg87kw7q7auYFoyVg0exSXzW62dTe6+2yi+JHqtkVLrNjDOA1doMfLixM2UebkCidM5
2xBY1Sr96uYAbbzY03afTmPD1RJ7phuo1yjOVyaMakTEA75cbqzvnXHfo/BkV3RmcrReS69BYz4b
HKEhA5J92cBOkF/pIeASI39gW9qQIkEcJR720txgfMbquPznWcWwNRdfJKrWGfi0SQgSqMVPtX+d
ModEiJFJfdc5N4K4UMX4EVcIBRTt7UfprTA1Le4OMRYjUEI6pRg3Wn3C65DW0Sj+Eeh6T1iM6Z5E
5pG2vbuNuQr0vUyYlJktDuE6wm0Tr8bKgtOJ1fhqAAWdCbsQoTIGwxzQvMcTEeBzsHZcRinhdYnz
TE5jDzHAihN+fYdlYVL75XdOICPA97rauV2eT8sABCbvlmeqTnFbZPwpgxPHZWw+fyaqLAk0KRZ8
DDf/4Jp28l+KaeZeVl7d5iJA6YhNLynhT1QjOIvD7FtRFMQJDAc42DXux/ZgxUCoFsOkxlpIKm3V
fUbbkRfk4reJI7jrLc/9/qxbhC8glLVhmopO5EqWDrF9VUJSy6YQk0Hd5jrVAXZjyvc1OnVUymaa
dXFC7znvMPjPx2oWUPqnBCP+jQC5rpbc7OjLHDPNmoujaGYwl/wcZqkluHuDBNA2B4KYDnCR/F75
a7WD5/7IDCb8G8b22RQyLQguogr6uoZV8pO5SRJYFXfbPpplA57orgw/ULrmd/fmgpy0j6bJGHag
jF4UjYAuzEOiwqjkSJKTgrcg7lib55j7TqLI+wannRLgcPNTOwuVm4oiwQ1dPSs1I0TNyFAhEjZO
bGa7E2A6ROROcgYoNcAWInz8oGbt83mzYOdFHMo8JSDAKpUzFCKkpEA4rmN9NKJlzFw2Tb2oOCrN
exkiQs4mrnDhnbyRASpzWbhFw2ozkd11bbTI/BxQulz6ZQhmN0tZw4HK07r/q2kLlvIImboWL2qf
YnnT3IzAZ1jLolSaq8ja22zLr3rLe5vesIQ4RCO+MUYU71bzzK1nNfPKpS9FIE3ebvACvQJ0OjXX
k2JhoDWyIUxqze6i1TCGSO4FIqvAb5MklZtSLH9Ti4SA8kEbcx/vNEIbRjGHGw5r4vK4WSRJpCF4
we/lladAwHCO1v0vzUiyJ2SgdKtMaRj7WJLsROXng8Fvt3YBAQpuDkZD7LcAXgba3a9k6OelAyVw
r5Q8OgLA8M+JmJF1Pu3Yy8h9yD91M9w+4mH5XgT7DJJyhcykr019QCGu9Oz7advIsuRW+EzyPQ+I
6rOMUXXIg0HQNQxLHsl3PxgKS0vj/euHjVKmt5KNiz/V/eFPReIpa28EsNs/Wta8ojDv8O6VqnPd
WEPhpK2YQ/TgWwalmIRX2DEIKAUG0inWnPP0rMHxRstJa74E8apOvvYC8Vwl+7VrJliC4MQOPiWb
U0x4CQGI+DfLxL/L2JT9Vp1cYTyUDY6MqXMXsp2KXQ1vs2Tl7nuemBEOwK5p615emv/TbXa9/iBT
YxYYJri0amSzQUbHV3RYIPGcYTg7EVdCeMPjlxU2R1DiTJDoO3roiM6Urh2Uc/MYFLptml2JqM74
GqC7OaZqoy2UPdGfsq4S9mqiytriPbNKc4aNnQPYgY5bycH2UIGAVODGVs0HdPrZlSYyzeMmVdtI
Sb2koc+tQQoVVzH5CPYE4YaB++kUjJW+vNpSQnD6zd6sKfrg2xMYOaXApqC8qz1JXWNoixYb/H3D
cxZ//6IgBumP5DJojz0TAbXDiydv/e3J7e+MWH9QMyUndpsS4yvPSmdDg306FdOApOZTnU0a90tR
ShgTrzjhOM2F37rcWSAcz78aRyOKk9MHmk5LyRMoxUlzSO3++wjAUpwetJVX+pBHoEJFSEcGwtrh
Jv8jXtPB7LdeBUyw1CxjzXXpbfDYrWNcQ5rvQHzX5jM5PRwLDT29Y+3lj541TQwwmUElyZ4rfrdN
Bv2kNjbUrvDIBUucXoeJvs9FMYyEf/AUepE3vnQuw0TAZhOthS3ioiKS1jm4qRMj+wg7+xLSX6NO
44pL789I5Kr30FzwyZbgmdQ3SmY0vlKq17u5HKpU5LSBu7kbl9R09OjKFpgdQrzWzmrTyal8k/zC
LL+6HDkbAvnS4Zl9HMORrMVQZ5+tnkwRA2moLcNHud/mv+Q45Q26gy8FCP+jakLuUMq4Cdo0V1lc
BclwezAwtRslgOEC76e3KUG6stgEt+OBWAjHjwyMHGhovOvWNGpqRiwhz4IrPCmf2S81z7260oEx
2srj+COLUcdie962nvHco9ya95i/V9pgUFZZNM5WFxKTZQnbYlULF1UPpTGER8fu/mzF96cmFdHc
0Pmgl2d2ngJdxSiZ3xCycOa7bKapjLL1eE3Bn8Jqz42W5HwkEdYMiZtPaZb3vS/Qh2jp0lUMyOhp
JeGdCcSACcFIfMMgSxJOdR+Ki1JGiyPaQASKhCoOLLb2SfFNJlDux5gN0ir+uDKPXBenW1d7PzTE
MN5Nhy9iDKZM8uLt2GEk9ujHNhNASPv/kxiB9Y1a9oD9R9TCsomXZO/SxQl1r5FHCJoD80kCBUxa
vm4EFU1fXZ5KpH7a00AE6Jc3rZxmFeOwuPCoQ9cixdhuk6FrrZo+NjZEPFfKYSoOTdylbr/SrLEy
iKrVfencrVOluS2qQaUVTT85mWb4lK/AB37dR179aPPUm1F6wEfA48tttE1ogTvOGxnd1YWvx9he
APruuLMr8jqOlqb4lKuGr7ZnfGoHiZpqrwk2pgaD0ylCHJi2yswUe93NRoNjdzhBZULE87AMWoFg
l2PJMKd0uy67QexzjyjWP1RqYAxi6ruWfFI853LpqPrTc6h2vv1uEc+PuhZA057zLyEADEu5YwcH
X1sMA+IzFz7/2ozMnhYvpeeKHdxaFI07N2N48MF5wpL6PMwn+ZMExaICvy8hl4Z0AIESYWzYRZ+d
RTJsT2bV3kHH0CWs6+EjYFPP/4aCFUZ3QcCMOzjEAx4NC9+wBNq0WJ9jvpRyI+zlsHZ54gX67y8a
HEaa/q1rFmuxDB5swLn1N4XZ51Jh4zHOB51rDJDcaGax8QTDyIlR4T75Oq30wt2kpdBUE6owktxH
dbPJzGpojm4zFAiQyO0/Hp1wCTta2XE4X6cYqxjeil142sRJVAE9vtU6355vBAsUfobeL1v2s7/M
tNFOuTmBTJY0AFyBzdkNK9i0o0rrxuuNnB8Cnd+K1GmVq0zcoiH6i1xNJ4Zees1mVhQZx08Ya8uN
qLXUbQ9LIj0YmvkjdpCZvI1cb84Y7y7uM9hu2GQHYmtMXOiuslsAgtrhI27dJRuj1jOmMUkD5d84
/OQ8HM3uTd97YF/NZlPYNtMzXZmg8PLJ1t0ppDq6gFWp4cvHp2ngiIXmRPs0c31N8vTp9fY1Yr0N
yfsD0+XoIyG7FriST0kHnHsgP+63LVFDwcQFqTBYUZKpTm9h++GSscS4RXG0WLvrNU55Cl6L7O9d
voFEDD5uv2cLrgF8wq5TRA5BI8sg+GPHZxLZMqa0cjaJt8MK7Va1yycQHzXp5LgR4mwaRezhZdOy
S5QAvhj/QPUK7vxkxO7MuCzlgVKfdYt6KaDuuFC8D8grzPG2DuAsRRPG8aoiglxF5ZHXuB6rcImB
Tg+heSRtWc6eNfIqy3EQ+qeW1GQgQKyYcPiT2eS+uyMdvxmT7PN6TjN6U8BkqNIeN5xbL9cd2tSa
sQb9JhXTfQwMJ1QLpy4uw6nPBgE9BRm/4jvlT6uDqj7zixfKD2g1RrZBaAtCkF7Y/4ZBKme+0L9Z
cdJrOwS94Opn2pJZcgEz1BleNfryIFwHuRMxCCLbFVKUrKYc8H7q+mzYNims1npwc0MX4zoXXgJW
CoXbuYHtV4wnfxl+SzW521gqo7h3PCmGned7NGRIa/OausuT4T5bqgJvbrmQzQ8TchwA8k+sJ55J
chUNQZ5Ybs8dXjTlQidLTc4eME9oS2k7/72O2Rlon73NIUmnMMCqcFDYr9DQaCtr99npJWEyqVlk
PJqLPbX5ea6m5G9KS4PXrCkjRj33198yhUKqHtMWVYulL7OtcHcsMpuNSjbmSotnq/ExEaUzJ/HV
uff20qc8byqoLuVUhyRdxC0UlQqfsUGaXbEmCgblH06trNLuhm0g1uVEerwIh1rkc+JTrHl2XcJW
eJloJSibyaEQdvWpB7q8ze6kvvMBXhWJ+CfDjBi9tjx4od3aiFVnYfBdvn3eaKRvidRCuhnzVS6c
mJL/MSLI5azQ/yBPBEPh+xSH+BRwBqOrbzx+qh/aS374kcbGuOZYHv3+Lz2Q8ZEOY8ra02Lta9ee
d4ZAvtEG6kmJ6RSaGrTtXvSTBmj7dLaU7PxTU+4/D/eXkq07dm4pa7POCeOXHjLtCeZU5PK6qfGm
X0M2ziad6mNhOvJIiIOHOycJIzhXnZ/41jWlbrVbnuW+TychfOMNSNg1R2BCQocdsS/O7HfKAdXC
Bdw6NCvfDGVHWA03DLOASR0wFb2wyoaGmnb5uECojgQfvyjhT58uDoboL2nGFUCY4WZ2NbjtyvJ4
4wlULVYD7+gOKOpuckxwwIfcpKsUwYTVt6kaUazmZ4dhU0xchR8LsgPWh/NKQohmTsiqjBcoXmvT
vDEhSchwcsb3Wt6lzt0OS1mAyxBa0yEsmjOrjZvFvEvVP6gBL2DEbBue0sHtTRelX6bQEkBKjyAp
wSHAIoQ6iTIp1w/5hmiUBx2ixFjmvyFl32DdjDadxSgU45hkOzDwm+i3S/o1SgPVNmp/VJ+GmkdA
/UrCC8qADliYWC9zrw+31rq0UCxSGgPcwz31Yc9cLBn+aEFeTLEBknY4mwa4/+hLCpP996V9sxFn
93nvVyAmL3Nv4mbjIsStbolOXQSgtw3JCqf16JsqqxYGsjY+vG3D5QF94rpdhen6SNVm726d7tHY
FfrX11u0NOSwDqUSVR5k/LLQdDGtbA+Dj6W/P1diP5DlxUlSu99T3s50S/+qAN51iohEwpE3BVpa
IpdFvm0igGKlFDMpw0iLl65IyrNZI7uDrEnC+JM6DJwHXVd1Tp8yxQwj+lPsYdULGtz1U0GNWFrm
l1DbClRRJ4WMndMm2JNgCy8kYPAwuIpjO4iAqMPVXPueIX7ITe62+rry8biWqQsNhZ4HA3wo0Kni
4dvdBHrD9Q8gUPUeNwjLKRtqoIsRdajn45/2vZYws1xOpGm5e56xTtD2uiBkqWr2kYNuvK3ieJ+a
W0asfuD0SlYxcQzW0yH4bO1JcRO8NjnXXqHBq1jG1e3HMtjcGvPGY2p47oDYzv2pupoQ4gi3ZyUG
dyuvU+ln3nAeU4MUfML2T+2mYzerqPhS6gAI1PiwMUxulF4R17GNBHPG3vsMfcIuHE/VMuBr8wMg
IENxTXs9L0ZyWZkndoV8XkQ+buVDWpQs4Ij5wapj18W5SMUq0dzqMg8r9no3FKmn2wdI+LyKFy3e
bCoj1XNhdtC3sWO45/0lRH4ijVEVDT/Ti0NqHGgT8AwdWe9XMrjNLZtT553Rjnc0S5RruaF3e8R4
bJpFHk11goCN+JB7ILdbvuJOGr78AQKx6MQ2lGcsA83Bop5yvaw90AQ685blP7DsDLTt6uKaI3Z6
vtnmJZ31gygLt8iBt33A9pmuVhxw4470nZAh2Z14GY2kbEBm9236TSDPR6CxEZaXOIn/rRT/GLz4
Qw3bgPyNM7LToxewttRcw6+ZKrfD2fMBVehOsoeEyp5y3szqK0F/dbbwRDj/ucKJ9paKSq4et4tR
dHdCtZmHfbNQEuEHyuBcCHKfoBq7D8D97DreGN4uYwX4z3YUW/brlHYxl9EbB7mCVuLuGy/ed78S
Uk6PWHqB1MsmuOxu7upJAWdPXMl7gEer/OdjG97eQK0JIGp/oA+fbRx+rQguKXQE6/lpuGCRAPl9
iXDFMTFQxVuPDlVQKmaehJz2echBQ2j94BzX3eBwDo9H+1yt4fhs00X9tmsEv+D1nkMwoBG/ANG4
yIp5ZeTmPYcXkgoKRWwxV76aDg28Kwbo7MnO9e3eh3nyv8k5uMhyrkeN9vPQx6oagLGp1Wok3Kuz
OTy3J1Nz8TzC1ZmHbK4KV9UcP154qCkn8brx82tBalTfH5dBYvtp/i+iI+JYD1vMkMn/1p851Us7
UKmESv1e6AlfcMaP5skx5wD0eBKFN2ER4SSlRpwGQ0zWOSaDvMYR63inj8rm6dFTMtxtJfZtSmIr
vN7aPAqnyP0fH/yPz/9CfJSz81XoT0Vwpnuu+QtT01Xra8ZEg6++F7q0gz1x1UYe7FsAKsRNn0xT
FC6odOS3lSkRKqW1Gzmt5qkO2w+jPCwMm2XzCSZU0CYgP7Ub0BImUFAZjOwrXwJC7KCxyKcBaL4s
3ujO0FeHKXOLcfA+/VgCVwxcIzFwcu30AcT1U4MBaISNaY8pRzl5B5ZhbEGu9E98F3CloMzLvJe6
0jw76UeWp3KzgefsrIiBLCylvWDrixLBRWPFgx4GmYVYgpneQvgQva5HQdsZDwtE856P7IOGtKyI
hurG+k3AqYd+tRE4E5a72maTUqkaQU3didX8qoPl46HmkWXiDtUs8u2NaCBtYhN1TWnwFXmI5dCV
DOLVnThQcowYwkgsV6p/Ud3CcpHCq0PTkQ1naXaL2NjMFHjfaJHF8m4+vMzbj6+AoM+SE+zLfwbL
L3be+rQyZEEYoUoXpIPXuYHfEr2nrIyRhAUywsArwTv6Bb1r8/4uf7YhXYYtUBeChL0FDVoC6qOt
MFBmaTLQpmLb11B4WE2S60kh/ew4oP+ot1U8NqzElyT2SdFAICdMKWJGhvN1k3fW9PCdR7dRuSpm
Bn0NsugFYzvZd8DDrmUizfUM/R8EdAG9AzjYFzG1TJp4iqPmSu1aHLdXG22PCqSyQ+EogJPCdwhd
9aumwvywvM1N9XPMD+cuM/0qol7Xq0MgPdOjKFO90AFkc72fn+fvAS5K+kuBzmhXifVCOjX83AlN
VNjCvz0s41UvmWDgN74GozZMT18N4nm+vkXNARDkk/GgTOKcOGTTNANAMXad10fRkHU9AWI773He
NJxavGUOjm7UVDTtwBrhg4ovzjbqXlYIZmJW2CGnB4Haq+k8C3mhbicMFCac/q6JDafRuq0HXCmd
56BA3gR9ZGqAqUqRpvipOH0R8Bv7lsFAk1FVfAUknP1EVpFPL+oJ/49Pp2GOuYeab8fT49MC38mP
5cDR58Z0tGFoWiGP9sY1Bin9roRdcqMaTxdjzoqr+uMl1U0YhMFrBEac4R5RVh231wOSO0gJVYNU
2Lr9UCmM/P1UH9vSLbgA5DDimX26IRRbRA/iJaqPE1mryaffNHXU/WVACOY1qusyY82923bo7Gjv
Sj/sR3D8OoRPoEHS0str8OUNV8LwBMfTe57fhb66HaMoVXamIGpfeO3mxhOf3nfIu0OaDY+tOyuK
peYxDL7nb3fYqMHz2fenhznXyKYV8thN8qlfGK9HH8M3frGrv11INKWE+tUUBrcZS8DdBqFDRSDX
K2F6EmDcdAFokqtrgwtPPGjTrxG0o97n6ma4xDoLT8Ym1IY8chxVRjbTKaDAHNSUIlIVwkPiUXEA
HunAf2oyoBQG0+MkGsT3qIoo7iuhuBznENtO9Wc29jFmrp11vvHdod4DSURL8caxM5oUGL9J5t/V
HjxwBpLkEJjS12O8JDzElSeI3exQbSYs9amyyvhZfqKn8d1n/QshsGpXMh55KgLUy9OMo0nhGtRM
r3+YW4zpMdkhKGwcinHrjuDm1EJlDIbqU+Mwi1b27y9rGZehv+iz9BsZae6s3wiQq7mu3IYXqYP4
7jvozVGEfSFEbfH9dNGS+/1n9gJsIT43Pk5BT+1aOch+3dp/xZ90uOGbzTOBrK3kJYpbbt0G/HMx
LFXrntkIUFJbMA+g5iC5T2UY5qmXedAMkpRYa73bSLwQcmueYLPQ4Rgw0cbTRGp1GG6RYy+67uT5
r7boC7aeEHvFC3pHHdE2P7IZbFEll0p5YP8LOmy2l3y5l4RALA5FM5jmvFQ7cHPpHc0lHW1ZHEHy
FvKsQMVZnYCLW2kRJm12Kfs5Eq5/Xvsf0yZm56DWFDAKwCi5JS5rKgB3/zZqLx8gXfZLk50D08Qt
pN7NWbwJy349KKx1SkbnzmTs7vELjLUP18LajP3bVGapdQ4eo63q07vltyRs948ZPA5Uox0jsTBl
ErBMpC9NIE3Z5gBeeQ2TNQVl1PdluuGJFTQXrY0Y8zFRBb0KGX6svaYVhc96dMfIg4BrQAyGMbKy
FC3j/kiWPQ+wWz420Teb61VfxQ88mWQlqF2qvgw2FdxPBkPClcdrvkMxlmTR5e20VtSGROgPX1o5
lrm0Nvtrqt8siulUk7kZgQwC7MNnRFPdY73O0j8QEmnk7V6px4dO+YZD6rhsO4qFmVQAEQek8d+R
6d/oQPuZ56pnVaikpGSBKknI5SwsLqyDR5HDdP9gSs9SvTHnT36oNwUVq54KWOYHztHElQzduVfe
6xwSzHulJOtDIcyYzoiJfTulEsVcO/gMHklDfcvT5ZYfvB/YmK2ALrSLJ0/cTsPqoNsYJNxPolS0
BjWN+iwbn32vzNWnq6vrvHcRGmdcRHPjj0O96oMq/PLTm8r9+lR5KjZxTyumxmisVOjAEooxP57T
GkR24MD1R6riV5+FsQmKmesANli3+7TvWm3EkKBguVHNY5baISRLqasRfjgTOGIvN1MPl+eJzjAK
qrv7v3K+CLJe408ZHGCFk0eQTGOtThholL4tFuVmbwkfNVLq1s6DxCY9gBImKSi1hlrSG2+9d/bz
fZs9EpMeD8HaxcHOHoJN3blrCzD81rlUnfd4jtxRSuBPvzckyo5IC2yW6ZQtVLV4NmdXRhEf846R
YxjddjB0IPG2oRu3YFE3iaNpUXL8FkN4yocD2XZE17R3vS3BYMWZVJjCbpyG79nJ/NWmgGpzdkmj
xwwornkPMHMAtfqhW+wF/94EYqeaRKXrs3Js2ZlSVvj5OnnF/1NxGuSVbJwFdo3NgUU3iqyHeSXB
yS8d6Nql8i6K/aOBU/hU3TCy1r68odtks0CIzAplHXOlO1OjLOKHTn0/RVkaB4SKcCFEFwmd0v7b
3OPqaaQmweehPM2RdR34uiwyXQ9KkZ1vYgh+R3JEKf9indF/JIr5dKnlHpQ9udwRl3D1bDkN5IKU
uzT2gtKTSbW3RvBaVY6DP0U08QGfJqrw28t2gaI4/xfVJQejqKwlGfDoBitxkH77H3l7poXC8WoB
jYb9VecOIl/cHcSZPxWX0QQ4jJ3HTKyYaTnxKT8bzT/CbTRTcPcmyhjUU2HBFIls1ND43d8fhwbZ
b1kZ8nAnaV6inwWZSXGcNX4OfK7IDaQgKy/vFxODooFP0/P0rXiwplJDWWVXg+jkhoE5rYggX6ad
Kgs5uovZjUMo/Ej0FBbuEw9vjnTPLXH0kzgDtVq/C+TCah/pSR8gICoYmuk4uOogYhq7cK949hHj
WtUtI5gJsSlNEKP+VxzhOrxfq9z/HV022cuVKacVU+IYGMYSW8Zk1cwu7PM86IUs95goW9Lwrc9u
eGjndfKFjAJo1SxQWsIGwMyNODhOGYqWgr1i/EbQRBywuIycewtXB1+nihPa75nEsTsdG9An4CeI
VN5GV0kuVrz6sV42uFJtHzkbLgOauAfvG2TtnBuqeGEJ7z0EYDmps3+vjWecDcBQceOCgJQc+eX4
0hdf5lI1J+iUkJClAlnW6k0HtiEoN12zyZcBiLSE1S0tWBzmiD3xpqNJG6mFtE3MmQy9iCJDm9sB
EnsA02KEMD8IxuaqnEfY2cuQYz3YUnk6eNZBkR07cUiMBeRIDjvms9/BmMN+1nao2JXCWbc/YFiC
YWUlQoiP0lxEiS1ofh5ixMazzG+xKxf1UaPtPsWTwQzQ+VzOMTadIV9gzgMHvji8ggToTAIVhKqT
MZXvyh1CJfx412swgHSCU7vnj7zAvaFBDnvlx03Ddn0sgWcaSaSrg4j/TyKH9Qr4yQnljs0xWcwZ
LEX0+FdeSqtKFvGvcTUIudIyzoiHPX4JoPtE1ctpJVJr5Kzd/JaRysSQ6AdRCcl+Gcneg329S7H2
vdauFDC54cylDTxrNNO0/KjE0/kcwpaBx8JfZfnIAQM6E5gmcjD668H6S+iRW8jX8v2PZ9eLdFUu
IrZmiowojB/lyJwkSsd9M7xnEWTOEfW2uPBFgKTHpG7E313lDUaXwZG2YfnQnOzEv3f8xdC9+pTe
51KvOSmrNn+Tr3pFcxYR2UKLI4Ig/8A6T36Jmo8F7Pzoy/xomD0P03Vn2BLn86mp3YLInt1N7j1I
E/Rk3dXyI6xUtL5u9dC9/3BII74VOavtCXJyt4uKJQbahNpT/bqmCfxBgH3Wab+CeOGlh1/lHpSL
BbxpIHNKLlIBhq+djedGrgiSZtfb10hf9lQChZy8R6BKuuJs8GYdpueBxRn6gu2ahvSGuMPCrWpg
71UzeF+5A1fW9gfNSjz580OzYdevoyVxL94lkrUAhbFzw3xURcsJk7iFt5RRjn14AR3l8w9c6NYN
DGdj7pASmt4gilwPcg4msgQ3w7Ve1aExo7TVovwxp0WRYpdnx5sBl9f2pyt2pcJPUVD/FZ/M+J6K
aPzXo6Pg0RXHZN4W9H3/Y+roP5sd2Lgh8D+TlR6rOagsGBz/pzozM42ABS8TcW14mUM9P2xED0u8
+puSERBpHzNlGz5rr2+eJ4BNgjSVOjcmwu3W4tegoZN96iTMEoPb9TBZeJ4y34Xx8TJRkcehgQNt
cxcerGJ+AL/X33f+CqE/5eSOlkaGGcebDX/de7PvkpdDvfckNjiihXN0NojlZ0ob8aGadbUPwvTa
SF6XRGngt0A4ZuF8NYHLagvEjP/twuRQqHKyC70uK7xZiULwLNUQCiGzMathZ44pev4i6ChMSkGW
OS+AYQK1zMhymMFamlsmAPiyUk/Wakq0hA2PRE2TAAcEN157eDDK00zmGaE64YHdj6GYCvijIFBi
sU54Vw0klMxftcw+4SyP9wgNienm5NwqY6BE1n71RBMTd6FPSIFL65JK877e5EDBzH7nwcB+NdGH
GyaOGM1ZpKG7FaIyR1/GmpkTARnH59wHuJ6KcWASGEcRCcB7BDmjHTV7OC0IKLXfXdQAeQeXD8fx
3LeU51LCaKfAZ7LQi9GrFO4Z7orwskTUYcW7fOWU100OnDzghSklRMk6/+KlFcuMjO4LBjpFgW0G
zvsNq38sDXo1zYs+OGO5ZIuSOJOhzSagcZqcW37F6Bd+9RHy63sOb0F/VtUiMqaHDQn2YkiWdvZr
nu2e3C25tciMztYBsTsRWgLzW1Eo7uccot92Ilu2s1Zn4PqZzY/bj+8RbXboOQhM4fwBSdjxLamJ
Ppy7ZCboobC1qcaby7HfGHl20p83qxMO5ZMq31LHNq6cNCDlJ+Ir4ZC5R70wv0YEA0iPTYrTIaTa
WBS2/VdJnTtTtto4ppcR3i4NXvnTd9+dZwmxTfmesK479PQuFLUfBiFly7iqk69HyBdmjz4In4WL
OcLJkorPUdO8tEhfSYisRhLX15IM743VKejHJm7AnIKW1XrOmcVaJReO541pfDx/B77sKakD4S0Y
5DMPz8CepkuF358XjVQANUGXyo6ORmj6eI+fBSCR8STaCCx7Kw4/PxJ4tqgg71YsxZay156hvpDj
RElYO9BZeZ4g+3MEbtQi1ZJikVBtTfDgk5f/yL17Mfbps1OIX7EPzpWW99toEuoxOzuv9kMiPZH9
x6/dZqKfOxAhadDZUoE3m1XFwWBnY4dumqe/wp4m2oIuQyUOi4c3TD0WLdH5wMBpTBo2srcv4kjy
qzrcc43+FOzhZpyslgL9I/8CeGqOxcCQAZ2I85LDJpLNONK7uJ6xw4o3pV0h3wqluNODmpbRo7Ej
0h5hH4l4As+80jhoQzL6IEuHyUghNGPRLOlCIIAXAtJD2Hpgs8iD6v0ZjfKnJ0Xoty1FXwNhf4jo
9iGtDQGCaioRLSi8cDzv75Bpp9xLpn5+1UKBpOxDLtmCwGV8pysbVmBtW3Kv5xq5j1bC4zz7GTxp
BL8lajIBdmXoBLEmE6HG0DP2f5IOIemAxvZ+wIAWa2j2e92XoedhFHiTZ+T2ggcL3AzzsS/Q34Ch
x/D68Cqz+xbjgmPjSiNYxFOwsg57j7VT73ctXOKWuXar3V8eB6fjmL/WI5mu5XTkZKcWLTaxPVVq
MlEE2Q9TDmxGWe1ME7+BJp6l7P/rn+QY7NkWUKxPO8br7bPqhn13QqxGtdsRPszGlhyGvE2mN/J4
suDeRjayYj3RL967SNTG2f31mG0WFWTAxeF2L02Ayt9KuFv17pXsVHtOetq9yfYPUp9KrvAbLB68
n2ikSjI9nxvWv4a9L/59NHJpG+Y6eFzgcGZBrieVQWRy05AOicuzg1kS58Yy2PLKMbgFLvGCWOeX
k8jww5iZMQye1HWsGcZxzrY1q2DGfkWTeZNbIP5G7FTULKJIuoOx4e9Ghf4RVNj+7AZQUzYO/+tU
x1L/1WDsxai9SgeiQA/s1yrl4VcWCO0PKHP93JAh97E1tfQlW/8KGs/KNPQpCMcbFcJMsblbTnh1
x/BWC4/iybeKHb9rO5c+Ie6k7GijtUDCuW3uC+PiaYXGyLBHOyCd5sr14874gR+MU/3ad84JPCS8
YpT5vVnYYTmNFzlKvR5x0XUkbC+qZCll7Il5BiEuxW7rM/5Z+9QXa7a70JoPkSb78EMhYmgDLu3f
P7jjGoIEIGktaQ7rp77amRXvT4s0QEKJ1c8+wWLXWZ+R2/wYWXe4Iis5MUHrIXE9b50g9dLmmEBN
LC3wd30/UFYm7nESP1aUmVikzRZfWYzzGFXlPMLx9yHu3CPNxoz0P5M3s9/LHMdJH4zfUhlwCcVX
0/KSbpQ01hr/EK4l/OCEy9TP6iDUjdw/Iu1Eu23sfP84Pc2BEM2HwwO1TE/z/h1rGEyCXwXRLQDz
9Ehi3kXJqIVmXyHUOCAWGGnyJj8vGCmbvlk+ofvETp9lbKe/jAEfG3Y1aMTWs7AVqcDqDRK6QTGH
0ye2r/JqPxrdGr4qATZSIXbxwbULEBZSofL+AqKwqGpouOJ4dx5V3x+CVk8FlgVc/s9RVCZyLIJF
l8OnmrEKVvTk1stIjDOe9y7WVr2lJvQA9tpd4+nwXdr0BGfvtPk14Ype/CmxXIuDpwf0dZK9dTmU
ge7Dd0k5/lQYblXpHZNgI85UqfsOatXIE36+A8NSGSNRnWG2Ngy7zcSEeJmwKZ2uabW4bI6UOswS
oVAkaD2krJiU7tt87vk3fv6tMbQidVA+TXE5dxU/R5BjqSqFBjTYZnmYYP/PQ8IyDh3G15ekFvob
w1ysBMNF+qKexc6I07a+Lml6GRSVFwe/avsliSlbHS7DS+cmGokY9/q01QRIAx8ry+Qc90KDBWRk
Uwboofq//uG1OZhSiWwcizfzA7Bci9Rio8spdh2o9GkyLcm+iLaLyhPYnGfLb2QY1q6ZBUggUaxZ
9z936ayBNJIeEB2ZH85302w9Io+9IdMj8Ljqw1U2FI9jAOvoRYYqrpY7tgjlKv6EymJ3zPeAbYd+
V6WV1zjrg+kJKpydrAm4aXL7zVhG4ABiFrsHzQX2ZH3j42t0lhMkHJC0+L2G3wRMmev2/X3VU5l3
FHC6guKl5JacZ+sG+XpLAd9LsYBR97vNpoPvGBxgk4QPhw1W+cXj1M/rg4K7+zByUIs3uEZ8+UIx
hcdoU33dqnzjPtPP4T4TDz5zMrJPHZUc0ywWWJpnVDhyUgf8OXBQokLAXPtv85jpNUo9OxX5XwNg
x3WNgZv4JCiM+r07lqcfXDUmLLpFp98M9qee/gJzWQtDOw9GJ7eXLcsw+fFjTwMUx3EldFbBh15G
VNtJyrXwF9PYF12LAnuS7l9cTjhvPYLpv/FCYS7ZhbR8LNFBQU2luYcKo0g+m26G9W4WkQDl4h0J
O9pfGPr/7qatMOZjdJhxH3Nc9oI5iCmPV9xVUEeYCjEjs4AA1I1SPCsXwSZTURCkiMhkNpjHzpbx
SsN6PRRD41jinvWITnhxftzN/Ysovzn6XEs4O5gSSaTugXGcI7HlQKWoVv+UMwirV8FU9V/lat+o
zd9Odqsv+ItbwIpl5wH+beISnM5wcu/Qh/QtiNhGcQcLr7dx8XwL09OuzCUPeDBnwE97w6Y1wn82
DJZ1X2umh5L5PwpKbQPJSzZOU+OaDgWFUYKppWv/ugcLkd2QUPFlbTq2VduEdZn/+ZrbeExtxbVw
5b6GxTccJdc+Ia129bHXlNEI1ztC78+WerV4doJvt592zWGaROzrZoQ9MUKUekxFgoV4JTXpmsiy
mWRCSQV+5kPkMMc63D4JPk0uAATuYNfPreXi4PgrYybzVvKas6AyQC4Fjo5SF/IQ3Mz8yK7ZcNbw
PaNBinA/yXGZTrwpDi1/QDHWixvQc5gjRAPINBUmrsifIs8EUvJZwqgpDPoUUOYaDDSvt5m8VAhB
WX7Fe5AgGD9gp75wcT5DHxxStRwr9ntoaWKG+iIk0yvqIScVO6AnQFrfBN2MulyJnV1ocIygYl+h
za0oaQN9xqMSQN/8R6TVjSCmUPjTpAADM7dcqeuJHK8zGIBsx17cAPBzDUkkw+4vQqz6NOtgDArG
iwom02cj88jTNFAvQqSDLRWmJjC0qgyPuExC0GFaXk63g1JIxxWJekr+RDpC30C0ea4+rGWWUd9x
u8O9RYvtTlMzmDkKW9XzhiA9Iuk/E7cAaGg1MebmxIbal8+vvrj8RsKq77U4MpcP6REgJIxLDg+p
vze1BiP+lWGUx21Jg1SrhH7s2F4XFH0/2b69UxbOS1oUuwgdRFewtyz5jayHoCTHySeBnhuqZwIg
+eyrsN2GGjEl7DztHTpTkq7Y0+hRcDz4DpMhweuNAepymoLLRc81LEy73mftxJvAxeeHl4q24A1F
7rTsII0ZHer+5N2rEeFkRSO03NzcVQf/gJIAttRW+YIfEZ65eCrSKc4JK1P4TKuFse6UYL7HdVOx
T7rUnVPwAAnkrI3PowrFBbD70KOlbO1RArHbDo04MBN6UJE+mqgepV4LtcIibJ1yjqTvI+qIS9ds
ZptG6v4EF1Qk2T3cPsdowHkeANjH+Cnhr+5C7IUy0mVs2uYvdQmy+fER7yuECgHjO2G25dyKbc60
jUSKQ28a2EdkRjtjTtyiQNlNBxjJfjjYfwkuCvAkjHDEk4BWkcSfC3SsEJn3TjfKB45+JuX+AvZv
3vqzuExsCcDF63lZXn2UjFuA7EYxXcLcDyHmtIorbY/pW9kimtOE2+FgcR7vy6tCulV2HeTc0UdP
RQER7KiTItTQ+0Az1zQSl826Pl/SpicgNDmoCE+LWNDxG3NlgmrWMJx4kp/6OOnVe9AOyOIWsa4z
8i6E1Mt4aqZAqWh7vPJ0LfsNsVEzzv45+Hd+5H4NNFjILNLvdE55KeYD3AYz7PuwPypltn5QB0Hr
GLVqcheNRToFrcCl3x11GwZAT/qs8ik52usxEsKtwnj00Jg0jynfYI5CN19floDAoi6a3vhf/GzT
BILpa/UJI1estD7+WoE0jktxp0FMf4NEEn/UrR5iTggw0HILi1z3toZgvcqXztkdi93sXbX8XQrw
2hClJ0GLxfMR1O0kkZ0nCFaOANuVtrMTWGFuyE44jvstBwI7uVrzy7CeXUjvWEJnqd9K1NnavUMV
/DJxJ9pDdKmXbVIhtJritN90WG56GRGQA6jElRwD4qWWChRe982QjllEJ44nN6hLazKUuF04elzP
zgokyqiIJgu7uKHhRpWTcMzl4GRQgAVmj7YvNrmkcwxSRWfl6eKE63CsbMWFOrQ9uHxGO9/oEKVk
vkzHGR9e2EoyeZNNvs+lQ9P5kJn83XMCffHpOj6iLCiFjzoEWX2bCku7XyVRQEL8uMpf3ud46NWS
NA8In7hCdyA8evtm7DxYZZaFKEo+Xtp3/EDq5zWV15zI5xZniifXxfkLH8GPs4jW8S8vTZNDISK/
n6I5WVKzxkGL7pncYUMpELyC1Ge/ASusmsImYYRHJdXMZ0MYyN339R2YAVnN7YwJa9r+7SOKV/NR
Cv3qrWmNjpq5ghnsTudxODtn+OPUWGzmyl1UzBEffF4HwexziR6GBUUEJX6ismD4NHYawJAJ94q6
StFYliLxDnK8WjOF219JxR59ZU+L3QszxcP4WUw9g7QuOalxAe6nCEav7fpJwzhLgm4p8HiMM3bD
JjkLu4lHATquXTiRPdpcfXn3Mz5gkgx1TrLF1b5ErNtctoGQ6VGAsF4TiV4HhuitF8a2DKR0UYch
W1TYsiyg5UZSKTb9rTIxKDalF16Ggjy57lVBx6jKon9+jHHY1qmL4PJDxhWv+jjWqTyaydHhhUci
0J6ls/N36loyx90ApCT+qYLu4PUyTpCSkTdsKB8Vjd1HnXp7XRM+7ILoeNu7WnrpfALplSVbwQdA
Dt6SEBfhsrSliVeE2k0nb///inwWTTx0OnN48QpV62Z+6vhGeynfXcxsVHtE5jhNimX3OLQDHgHn
Ho4umYhhibTTS+UrQTCsc39nlUhzetq2IQFgggKVyQZVZdG/g1pNWgQ1bgNdhUstELMsOWD+e0Iu
EDJPVtdtxLhT9uAP4FbBLOsMWkvO0JZ1NPsNr9gaz7MtqpY7BVpKmfzFInzs7dlh2UM6RFsf9Nzv
6/HeZAbGoCxhR4fLpeB2LMfzLxQnWEr7yL3nhBnQhY/yeNVjeK7vgX7n/ae+25dyYkKTP9AJjh/g
Nn0aMrVPD5P+0/hlRkFP7XbxGhrwgMFQkXy54NptN2YooMlr5jigbFCm0uzBRTf2HOAq2AMnUkm+
BdK5yEgTaSB8IXZmEbks0w8BWI5jwiABr4tsh8wPjoiLOJBdO/giFxeH5sjB9SqAoa0IVWEH9/uB
g1oqVZozVrkKkoJV1jHPzUxVQyogOsr7DztfOLJGOw33xIv5Zr2Wy0e+cpd3x4Fgfzc5vZ6ihsXG
xtx8O1KQnBB06hGIgnB9Aa7EDkLvzt2Y4iyPoNVmapsFwjQy5XkNhA7mmMTU4G4Ynu3SHA6ZG/lr
gfQBWaFCemRF22CDWOQLuCMzV+HC+YN5Jn0TITvvswvyo+2wfXPzEpa5pPD9Tl+z2APnU5UIh1tB
37KHOfnNv0hl5SRTkx65mMDRlcKeiwht/fZ9Xg5s1L+HpHJiphONBEFvSlAJ2659/+6jxQfeOnTY
YBqPMkIrqzl71weZnDPm/+KfQX1Ze+fERfpC2k/RkxwrqL9DmKkP8uepIj41Gh2Mv4n7xm1aCBg2
MuuJS1l6ZH51piHMwmZ2eVIz4/9u9ArxMaBFobX2yUmcUtGUTd06FoO8jqB+qZzY9+3XsXA6o608
scCxNp8mDwroeEjyS1e4zKsb5mR3yrEucCMxXa5ZbfQGC4bx1pletCBoEdef+V5SHUXenqomAAba
b6hCvHN9S1sM71IheApWQSYSY3IFdpVEzMb6Xqou/L/qbcVfz5dxeBSsYADgdmvxFJY339H3zCYc
gfhK3U5hUP3pNidRpYeAvNsBYjn8KPooFTZY4kZUrXQ+opS5ppN153yT7lFmLqtmBGapduW5hTC9
dt168ncDsmCntBEBCl4DsXUlrlSkWupKfX1priCkYqJ3mGRrYVZeCmZ8jhqfShN/94mY80f2B3jo
ad2VvitnVri62y77YfAUJCrkOYul5yufKTXC5rmUixGEmplh798Jy1Arz4tOSYK9qEh8Cnb1IGxe
WPUZ0FWRzYC2PM6DoPnBLXcOyIN98hdnk4Mqp7+5G/3VQia06HvErdg0dH29g8X4cUlIjIeOTguk
WXnwyFF2EUeZlw7kP6Y2K9+0l9u+G9NHcXNK5p3PX41XGu3Kv9mMMOgUuIBKVA2Qh/2A5dK0zYsl
TSQoBsPMp+OuYITOicev2SAIg34lQXkhKlDDdEu1KSbbImrXHIGBSbl1mYrhS0Hg4D1wQsMPNfEX
45N99T+4sSXg4k0O1kJYIedwjtEcOkFTP8FthAkeufnyR+XgtncX2MwEa/V0QPbIenHYG14VqJUj
XhCIrJbc74Kl38TRsrqxE17iynAMDzPeCc81rOF5I7zu/3ZfElyf/L10IicohOxpOUQ4UO3ekbPV
yjzwqIIrA/o8V94FOH7vnw2nhN69gnFahqGG9cYymni8agBt3yoK1iJSWQ2LOmH+tvz5DAu8BgRJ
jvqSoyU8V/P6xWx9KUa3gpMISeOuMU6beRG3AHV1n8N9Z75HZTsFqMrni+/0NuuIE9ahOrOGhGGX
Kaw1yltq6n/VgdV7YDN/JBizNuUbBJkNb62u5OyQjcPl6T4CDZYjSRvXvSGpK2PRA2u9Kvm2Qehn
adkgxrTvL/rC12tcdwJQs9141EMyYlXFhUcHKuEapU3WgUdsZuiyU1sJHKHjybz33amgOPvDXbk2
Z+PGeRPp+SOGp90Q+07zq2pLNOz4WEbTh9mbkDF457574hSG+hIP6rpnIq9xPMJx73cPzZqXEv+I
ux6te1lEMf2Y7RkDnZvEjvw8lFvEuONQ6zpwPtl5A/M5ifE+6PRCYonGVgZ0I2q3OcLSlRGK3rKt
IurSQchcJi37T5EkyNdMJVb8UhDHgitVx9KtLNBRRBPauTSxe6RR8LO2LHSLORNZ1kxaEjMUq0Mn
VFxY/Z0K58sc9XVu/cWJ9gjpr7wcVa3RWL473vMBFlf/cDEtDwJ0Pvd1ckMbyaLIW4BlkMObBzxv
OJ7KC1rMOiG618ypbSST5xhpuX/0KgJJcux/1ogS+aW+K3/+olduX8TqzqZQZ+NHrOBlcRlksOfa
dnwTetjJ83nzhl9+/QeCmcHNn7iRG7cT1sYjoBf6dcYVJtqYkqDx92tMIOt8AqH5y78x5Baz1X7O
MGQOIw/Lgs3d2D3ZmdZjsoRG3AWYOhs1ON5bkoEwC++AiVSr9dQvl6REFSqCuR/mDqKKNYdqXX98
pi4z+Ms6MDPLUkTLho/sQ9Be+OWudcQO9qHJqOGKDiKDEUddOT2xGgDxn1tvqeytQUscBK2t2veo
uOJkhC+4LewWkxV7ltv8GjEd21foxNTHIxgLQAd4e5Sq8Ay8oHWpudevSs8LWa+PUgjC8TAeISd0
KbUvE2LhPWS/TElFnc3an5wXrWSbkAdCUGDxgMtgWxGq3wYWZjzhy2Awo6cDyym9C8RxFbqIadGH
mqK3loXy5XxBBXmJ9jd+ItOJu2Ri39Ke27XvSrxpWvWtL7q7k765enNRAKF5rLSZ2qglO8/plGSj
MEJ7Fwthe4BpAdyoucV0LF1unRGNRhuOL6xg5RIPrdaYOhuMnPQHHWiDNkiLQ+pfdA5suI9V+Yfp
OGKPh3aZ9RCaFY1KkTf3JvJUL0tfEqWAvm8VViDCImuaPTDRuZSAe0JQXKxpaQ6pLF2mKctxkVgt
p3geKLA9PJZyDGfplr3vmivBAvsF3c4b0hZe3u6axKn4rTxb4d68ldxwS6M1XfBVV7NmrKdbT5bP
s+V0D/QnBVip5QyxiJ97UKb4Qq+OggYa7ya3HDHz820xoZ24yUdaKrBEnGI7U1wXQi0GVfWM4M38
CzhdWODoxyysL4W2MpW71K0BtFHdnQM8zqPWzcVyWFqSYgSvBYXBm4S11yH8nMOPPRzgmBAEGbW0
iD9gm9nJsmjXDvs2OtWJxIAJpDjn8MRdeRjzqfP5lKKRGBSJBPrx/Ejb6rT/dnNk29rqG2VqAoBF
U/isTQDNulH4vy68PwwbHR/gDZ8TXjF+NtLg4X8Ass1dbn5izoSZL9yLJ8LjW8fFXIsc5LYN+eCO
kF/IC6AmsKqM6+KB7QIhMYXlivPsKrZ8gLA0TpkPcOE8IsVhql0JqKQgzEVJM39j/ob6BvuP+h/y
mwVfQvDGi55Ba5KFkMYQAQURz1s6vCLVdIflgv12qDbqqylNkoV9wa1ht5e0AU5xozCCZwZ2k+Dx
aX+SPzJuOdINc80QmVZ4QD3R1kk6Ui79KPOP5ATWWFQaH+3k2UiIZ/oilqq12qylfgx+VswNm9ii
juAjQFTq+lBj/QmJZmh+IXSolFxTSdGhFsmCV5TtHvpMB+9Y+vueIprVwh1j9Cjb6G7KQYYEFSHc
RMkVI6SaJ+LnbvA383jaTo6PlNtU9TMkurpMyzKZnMY2ZVEVY0nm3B5u4SMt2ycqjCf4UfN2GcvH
Gqa1By1V5rDf726COJcRTO4H9QLAfVZwMLXqKjN8MXIUQSBtv0Dr21PCuXxrAMhAV/nNLsoiMu6Q
MYu+9HH6kJqJyW7a7s8YMj+f6h8T7uwSMUZ8ddT9J1u/JGY1xhLnMzuBOSBhYpq6uZsWdmTGMHHL
d4hUsnaQ21i8Rrlq3qtYFI8QjPL9mUMt3rIkumAssigEtY5k6/GKpqZ3xq/xT6QU6VKgv0uflF0m
Qwk8xcLKAD8mnZYUkhmEdxUJDm/iEjZTX9vDmhjvqiYV7Fhpj6A+zEETWuZHQXhXRDDg1AU2X79W
0T0VREHuHRDqvdUAN+osxHwdgAyu6qkDZ62x/eAR90kwz2eFqRAynqfD7u26gA4/Py8aZslVH3cY
l5wK47b6tMYb1PP+ZTCCDY0SquTZIu7dObzXJEQs4dJViEu5vuuz7Z8S4iTxFNDCZlyIBFhHdr9+
C6YqwllDbsvMeqad9S7NO8SeDT6zECHRAeTwQcmHKwAq/c/dHelRLaS+b11YBuB1CYo9KplDLefV
3JhpeTTqujpSlEw+5igywy4qvGTc7eBcEkhKqnnV3T5YRTKVQuRepSvVnqMNEOp0xhe/+XbZG4FC
8XykBaPUoWjf1gH+cYEYZeiGzKMBx8PqAkFXD/yzTWe2gXnpz7rfxy5q1EVF+Zu0SDfn3s0EXLXx
r2QDpH19WrTqH0jrEH3qq/YdkddxhY/y3ni1qZM16cR44wnO3aWlpbm4n2J6Q2BPZVAs8tXtEAWb
QRMEas8E9jp86rAVfrvhc+nhLXsrfErFbtDw+Ymm34Zm14iiw4+lmfvLcFiYLK9gMN+6wrOr0qNM
h+wu8uPnN+50BdN8C8t+kRk4EzgLuLMIih923+OA5vyYN5KcNeqV6L8eVHwds0zCQg2GjhyNcSk6
ngVLnlXTsL+RN6H02R3DWgHCNUrZUZl1L28WO84SKI5FSKXAxPvRcQAzNQ+y9P/6vrxpBzILqx/U
Row17TMohY9Sidg1/70bR53wgstViGvGfRXuK8kHmwsqT+xhOd/UTR1/SZ0f2DS2uCVOMlAe2pmw
aW/6NNj15lE/zJi+lrvubLLpzDA9bT8SneQVjd3BXteJwAo5nAWs2x/V+FDigGa9X1smxNAg932E
kP/oZj9zmb7dPZLNNc610/agJktQ3Kj53gBhEjGOZsTbXNbFQW3IhYIUqwh54iH3t4VtD7tRF+Ey
1QqvHAviiJBnjlzMWtPZOcAilXUXY8lppPAnMwbxYFglndWDiUl7yuwBytdH8wfRD7ka4ZyykOUS
FoQtMOKS2RkA4Zqs5kk+0APSGliYoSkTUBK+ii9SSju71h8C/ubdFHt98VR6JyFLYs2T9/7RooX+
tcc8LZa62KqVGfM61NeNguDAytAX84lggRXRsCE4gPn/tia6RodYM5WWx2+eIXyg5yfbrE7yww8g
vDGFvAmJQYTQ/fz9xhBtR+HYKkd6yyISuly482h+Ij4FOz6y3P+j73PW+9VgPJsG8v0Xvy/VlJAj
IXiZ2n+41ytfqTPuoAjOPEmbApMBsoHN53DSOg0UljtmDKSx3r1oshCx6ebpw9ePLve8F9yyDNOn
HqfMvOMd1Q6ZSRYx1kiDqxSobgMsqm5OIJbzDW2dUoHEoo8WuNmRlwvhPXG2W9QWLKmBTHGQxHkK
X3hwMEWSeCXcuvW7LFrxf2o/kmKoPzrOpuZzF/d0TbUP+TWBlmVXgou7v3wlPzdzSzSqqhK9ampq
UA+tXYu+ewdh2ZcpcfjOsyw6yxRji389Mo8BdLGGghhyVDjUc54pSafaO7garE5EPFV+Cs5gd1qM
+KIS21n6Zrryq2exKZywr1nz/wuurSqRD8MX/jlJY4fr7vbnq+0RpBHeqPcW5/ImWMYCdyI3YPUp
7vZzdHyB4Sx3WxBr2m89YQ9A72SbDcKht7SFzYF0qRwwGiHYGPsbcHfsh9905v4fbrKNB1mmcGxP
DCyukMEwxAOXzDE/ldLowuEa+rodPX80FiajJqge9b8k/nzm3HzYYNRuEnyf1b6+nAMDbkQn0omw
qkKMqZOzzdbXah/r0XJ9pGlR7exdMkt8IDMAfyvZUrwiEagNYYc9/6W5+bN4071jg7akfr7hKfzA
cddIKxRk3e8K0gyllacsQ9b880NHSTJcoeyy4lfGPyDqe2HZWuRdGLtJ2wLXSdMNzrnmoRxJM0sS
D8Jf88CGzxa6xrMaVNjY8DKzDE9xofp2T9EWWV9WZQRxPB33ReSPe4QT9mRhTnOsX9pWuiMLzC5h
b6fytpZwJ13Mq2M0fANOGEhYIy3rkY8L7t8u1Kb9RwRR0hWjnAHIGOtjFeYKCZOlOYMiPsf6uAPZ
Vd1muNTh6vikiNSwkjvB//iYIMh8JN9pursRZbLBw0u0WjTD0t8KIb7rnCBCjEXsiQotfI0syP7k
8jfKC8wCll3HBiZyafJxuCciOGsM0B8Wd+VDxXFVESgOLfaqMGZK3n86iUYOxd2CJBc7LOiLST4u
izejnY+5cHFufwr6LhT6lRqCs5k9opBE/1G2r0fjCrixsAJ/GqWSttgkgZCg3fV/B8zEBV3zyTJN
BFDvy7gixFhv9UOXSMLgJk3PuQqBWpnEbhZrPPnVS3qKRELLXS3UjkFqrvD+TvB21RQ8FKD06Bd7
7p3BCUCse6UZ1Q92i8rIifSje1uwfkpMT9LyMqyjOof9HsoCFITxLGDJAkKQvwEPRsvIKHP9rq5+
XUiyTlsSQc0ba3MWLgO9Anxo8CtmFyJGcj9+E2D/CNhU+6D/eZ8a8ukpZLBi3BSKeJcBW+Yr9LaV
uTm+Luo6QJJPkkUL3fSxhg7DJo5pbQ+IUCIL1l/3xqGPxgCjgIXEj/e2hzbG3fRoT6nfzW9a+1VW
u/XfzKjkFbSs2Mk0T7sUh1kPQ/g1lrP7n5QACgiTukZwksd9JaGdt9dQwMw1xWU593ppWqp11UZO
hpPzdJs5o/qOrjKB+VN79y9H/GK8LvBJidwJuz6Imll8w/WTZgoG0SsDNTQ8trZ0WL80/j4YJIqc
vlpIw4PtCJHa24LboktZYFTq6IsMh/bQ4pTDbAxlwgSrPaHju9xUMcS2Wvvba7gDEadmX81nr0Jp
sDN3DVYk0IZW7/V1N8F6Hmr0mxmNYtpPhbqG+DVTAdmiZvOuOewLPbhrOUoNVfHI/Kw83Qwj0q8w
qvjOOSElBZkMVPY+CjfjFizqsspKje2TlNXXemnlpxNtbOXzjHqFpW8ahx44OYrscKvCVZR+QqoA
Q5g1q1dw775TXFOTYcwMMYIC52R8rvVnWYP78CmXplmRBPbm9XL8f1EHbm3NvDR/qYBUDMnPcvF7
Al/2SbWsEC8we8wchnSxvoK0mE6mMpOoh1RFChjl4+Q7lcDWnZxxceydvW28QdTMFXl9aJhBrq/M
tfeaSfC0gWQQH7LjD8wWImBJQaQye0nz6/6j1ttR8kIUklyl3Hyu7BarYjw9lctEe4h4ANjJ4dVQ
PgIZij1ots2j7Al3D7irEb4FbSqiZQ55+m/+9CULSdeOYTY7CBq/ADCCi3aakT+HgfwCfuDd6yG6
qhdXCtFbw/37wsBHlocskEPaU5x3bbmGRM40buRDW+mEe7+u7hQQCyJm9isoVzf3GAfto0GNJXK6
JQL3buqh1AibFMN9ghPkS16dQ0KwsE76acRpo58Gj0VJgV4+1uwhjud2iSLDm1/69xIpXOD1+EJD
QZpsBhXOnZKWNP0dxABarFnP/pyM78cotuSYTb3t9B1E2K42uP8qrlSasGlpC+ckLpfQ0pGEMmfF
kZCmHaFMOKpDMD/00dUMNmyaUDbFtdu3ZuMmv4reQGU0TzFo7Xsd+F4TuI1EaVnzQ7hAbplvYqzR
MYdKhbPIFNK9gJLACgelDRJVBtyktTUW8MVqj3RKf7kElFgIbPKo9IrgbSb4Wwvf8qXOfZY9A2IF
dpH/48wS8sP5CP8YtqqeCkhVvMnJ07nymhrbIup41dNCpKdrjAny7WtKD1VjhskhVaTfyR9a2VCt
MaPdxRmHQbcdyNlCNzcghXsjyqDvkrF3EZF5yvIv929C7AbSqk1bphCyrGpHYKrQRt2buTlKuH1Y
zOHblGSDPzi8mLztVKJZULwxLMhrt6TUgfou/fZQiat8HH5kLqVW4g2ez28lfpehRsNC+fXpNQtp
AEA9lvNG8FmQPDLpyTbZopOJc6qMIm2xHSkLO3/E7cAeItnP0KOFDJpXs09sSfZpo67PoITBAT06
Jliqoi5jvM816S63MvS7VC/2C72lgzkz9bpylz46SDR5yb+kuDKIzdKvmBLPZgHQyKxjHeUwC0qr
CAlr8Pgct5oUKeSTT91W940iterD6OVlVVtqed/FPESog7RkSJ207JSqJ0lXdwcd67q/sVmfFapB
F6B1pF5PrG1c943sclxNBUL7W+HwyExDY/kX2iG52BMdQr35wzKrVTKiZ/vcahdKMUG3TMx3l47d
+Pdk2ezfOG+5bx7ZimGLXWLNXPGhW4qF0VZa6D3w9Cc3OggBRlxaD1r0fmS82X+BtQOu3oPGYQw/
OFYKR36w0IrCTUXeVk/+tk8lifW+D78ZI0d0+sz2zTDZg1005haM6T0zpsbTsVAN/nlf0SlA6nHQ
XL5EsNVxtJ4LFPsweWUnrXxy31uQd3p1dFrHc0G1BrLjN5Ttxud7BKU0QWeYKm779YtnnSXJLszl
3UYKR3MPPgTC3dX/+z8LYnvmxJIn6814qJeiIQ6UMVKbGLu3MLGc23rEByey0HwAGpGS4QEQ4pem
5QJOVxN3gg5Asa3vBheG38X8HF3ZUHU4cCtLf8KslSxu+s3VBpr82KG+BogdQfHmV8UF8N0D3asH
w6qNIhWFIw70Y4f43XOb2lJZJkP9MJVgrFAJhezz/QyFwcmDwYokbdLIqL0wu1YyZAW+nx7s6Ca3
DeJrxcaZVwKHIp4zb1vZMi1Zk+6NQerOSXNcBnORaSFPl1uXBaDLQZvesyDKb7g0dyRTvqUgOxIj
QawHmz/iTAqVhdM4uk8QRlOs+l8SWIp+3iNys+SXrgOhVQdeBl+NGGeG70TN3ekhOsDTGRIbJ8Hg
pgY4wrPjRv4CeqvVKIPBdYIdXW2zrrmpykOcZ+JK4g/3Kv5KuVudvtbLoMEtz//sWRlu0rr0VU4d
HgIdoGQM3bs1gVySIfTxgtmj2O6uKi+aXfODk6pnw/GV9GWUImW1jWEno9crdZCdtkf42NoJcj7V
Gf7CpRq3z73M3iMTSpswP04xc+aZ5WG3C70WISPVMhsB1Le3TLl753YuTL/ntZ3BWnbtYYg37fZX
iAsM4cmXtFLt6yNwhIlOBeYFRqkMEAxFhIOl360X1dGb2DK7//SJc5QkCXb7fGWAflv73JsIMenO
t3tkQpPC8g1ja7vnr0iFBS+zXh28BBj0bCALwYAt2pJ0MX7tKfk8h+q/p1wxSPEdnHQp2dKfFLS1
5ecYTeuXMx7mNqy9T6hQRGWkBwUfFMYGC60actASgqk3l91bPivzCOCdCbPOBMh6VLVOngTr9Lv8
WXmM79gwa4pw3po28m+3ea4MXJwvDTglSiwBodHML58ojAh61ubocEWyObU54Utt7UVxWLkEGyCV
c6in7ziqgdZWhBmAHt/1RyQPumcZIEMdIrbUpUGIfVCbmLFqm0JAC3e47hyf7t0fLGMjVFflAPkK
ANYytwDMG0c5CCQMMzRmwDEnSf7ZAHGDmsHYpUdtgCn7/IYpnMY3yU47AFTHlGsQdWRTBsIVGR6c
N9RKyGiwg8WO+GbvEiOp+3/Z/nPv5GTSOEeenWQ4WnXkyn5ifw8YcH7u9pL5jKSdHFPITJizfEUN
Skc1VbTLgRYSeaZA8J9hbfC+qS3i0XvqEa9DN2wl5WIHgC1SAL3i+kdR82YrLVn2XoaTllcguqYN
hMa63QjRffWb5yf0Xmwc+ttjI0bJjI9jlKxfeviwlvZ20YLxwdNDmVpVJXmyjnKsNFXteySfdZWY
qR3JbLo1xyZqoKS1b7l3V2u/KX1KwFxxKexqiqaG3M43TiLqsQe0620I+tLtL2RFsWNFP2OkIP/p
c+lcw5WUkDxvHhPeTQ3o8nKWZb6junAvi0bhBrpsASPlMcXIE41qwFgSDs81He46quMA+qZ1046y
6lw2/wQThBomdGPCrytsCxwf4c9zNnXr+TFGSGNMZbx7mZ96WtvaGSS6SvNBRoiWKxkRacqgB3AK
4MUr16VWJWhmwL+V3RhHJ8fn8kmjphvzYx2QZ0qR6EI9cdZjuKVqHbxWap46oAlZjXbr8m+F8mmg
UJuHcIFLvMqbdLg1/6/3D5TGjxTQnjyS8HbF4FTI0uA7x7qnOKq1V9nNkew7u7FZ4Sf0ZNaKxEI3
CRTQjuhYxtKmw+7Af2HxhsNgcg+SuuQU4zt4g+Sh1Tginy6j8mJTT7JrvuecQ0sr6KoCJrY6DNRA
oqrRj9qQGnSFHyjHFuWXzestJpdL9OHcaLT8GCt6zIVqJRcSbOW0gZ0lfvwaG2m1Q5NR7gJEllEv
vgfuFHj2E8oj0x/2DAZBSdudu0+X58dveWS7FUz4JYGo48L+0KSbdN+4DCQVHz8RWRtr3Gj5eVMn
uoagqQ2goND8YkrFcwFm6onk1qtZRPa50rN2d5Gck7/ij6erOafpJkOMA/6lyX/6qLCh5XSQJdCj
mTFH+EEWdnGZo4XuCztGiPxt8aJeWAiFwjB7kI4adLOpNVBBLFu5PlyJizpTlajuFjdDme6yugfU
0sL8FovUxIkVO8AM3NIevO41+P3NeOnZHdghjECtY/xzllHPz/72aJJ4eHCB426z82PdaCISfxwr
JxBrf0CwGWPcwADHjwRKkV67eMVTX5k+Lpp/JLRmO2BJQzGC+8tS9HoRu9jArn4/4FjKvGSV4OOd
6mkzRxQ0nxgV0EofG42x8Z1UfrYG10PqMUfu81eos8BSXOYM334P5Ear+Bci6dO6hZ5Om4tYESoL
Uxg/FbZ/JUiCSMt5NU6pSDjdGSgDdvKOlsRIIj2ZaMpQDPwNlCfP5X9nw94ygvKRBd1JgNoHwj52
Ajr7h8z2bDK676SzgFG5SJnkQY5I4Jg6WsfDV2xa5Dvnc5JhEhmmKf3IdhUSKNunNfRSwqySdw7I
6eLc3sU/BS8TUG68rferPWRlGHzxvtqgEBPIeAUnd1lB6nGsQIuhSTNYW2Y0ZX5vi+wxFVIc7US6
9+gk8ywslPCQHe8JryUPC6VnK+dXJ2v6CY5G4aXKOVxuwchOFUebtRGGS3YEAxOfGhsqbKbDWVY8
c1dgY+PHnBuC7ijfkpUll+TrLUvZ4gFfzVKExk00t20LumRDsxsTcL+rx0yR/wpQq3uTqAF8CRe1
DheS1GyU0t/688mCwnhhcuRiWavAw1mjkKDXfCpJdgR1xoYbglnxti359U5fwFz7dn/se0dY8GWQ
bxlQcYE/kGcwKPiyF9+O3hlpSypT/6BYgRgkwNRjxaH6dJPFPIE2SDmoUtvBkK4DhSlhZdMuRqo/
9ik/9Qh2mkFSszmNjiaPC/TcDMb9y9sEh72OYRn+t8z8PoycyoJ1GxNaEti4bht3yQe1Siz2LDya
Bzckr1IksRpQc3YGx2+EwDcq3mprJJhVsOxm3pYnOsjKFWa40HkfCZhEtJbHFgEPmhTX5Ju+0yfJ
vtBDw96oeZTzdIROeT4PEyRFnkrDMeJ0hO2DypGOGeATfrBQJxdbNRn0ZXQIK4v1MRms6MPcyaX1
wZ0MHh55QY0XE/9JQ4FHlwlsEImiS7P6NxNS6LX3U33L/doRxvInEOqCvfxqRIPvp6wTO/S5kfsF
m1wtrknSPeITMhtY9qhjDr32k+OpyoOgBDOBVZEqSsNRlMjIPCiz0NYtW3fzW1ykNvEsjOWi05A4
lWjiMAvyxOug6dFoXhhot1/vHXxhkTdIj/wfysI8jiyW4WvcNa1d09LgZD/L4FtUZv8VjUa29duB
y5blmHrIRj9U26c/TQ1tu2xH/DZiF/WDzaJejV3Ff10DuqX5mawpWhEE0sMWG3r0bcpfoRRHIF6C
GOlH0VStUh5VJkckmJMLWkIf8+JxJJi0XFW79z8MseaNKEpkcWcNKnRsY7fqHzMRarUVYtWWp7mh
j/shwYUEDONzT4f1uguW9irhKvTawGqm4eRnOXTb3GBeNFZmj1LBkfA7Gk83TaGc6FQrNxXEO9nM
yPQDtw4mDvARPuHDARpFtzkNJ63p8BTCyv+vz9E4MdWXgmg3353DksjOrs8xe7Tr3TR2Xt5A8VfQ
xf2ayF0PQOK29kcQCJc6P2RVt3WPcQz9UmHSnfY+9gIzU7Yrlp6sSbh5w6v8iU09cipCdSMn5qqR
ZsuEsyCnAeu9wjuyqx2AelfCHLk+MDEyIe78ha+NP3Oy+9VkhLfLJYoLmJH9p8MENpW9mvl8UM5a
QK7VW/1KXZajGw5efUgJpXt7muoYZFIFGykUGe9PWWHH6Dsu45W8Gt8kqTaHNFU305NrUhCieDJb
hYXioXle5PaRt+JuHCtgYxHdxJ5apJW8/RGBumNWRPFRoRY33E/PYy8S7FhogjHOxdm+BKr+feTg
TSfTGsINl1BefECvYbIOTNkFIz8Tso6zofRShpQ9kLQWmDgtf5+0vf1j36ZnYAeGfo9VYVkPruhK
1254EgjSd+OPZ5mJr71UVyHpQgjHUm0Ey7cmfMXZXIIBbSXA3mScBm/UEhQundVjrJT94gt0Lfoz
VVs1X6Wsfh2X5I8BXsmN/aHfKI3xTXyIDCFrBh6SQeBkx1WQizBuhPDwZs4IPQzT6TTOLbYU7qWc
2kYCbDGB59lYBiY9oR86sSb6awYp/LK5Y7q+OYn+wAr9uxAL9Lac2WtPQBv4HUjfQIsTVOymTNqg
hT1y6MVIt9raFN0/PAo3Lxq7sYhBbKymzBAKOcLPhtvnlNfE77C/lzdEhcP4hJUK4/738ikerVJL
QK7x72sIan3+iWD/F36JzOLol+qOqE5BqJqX18M+fFktCIa5jEpxtf0qyM+OgdbsXPHZtFc+3W+D
+iBjLI1VVkE0dN/S+AIA5umtVEy7F8GeNfOZspI+WubCP65bjEmDtrV6vm2vX7Gx0R5BjpXiF03/
sWEy9i0tn7ijeZ6NUPpDJYm8KMUjIe6XG44Triknvw+c59UCMUMsIOAnGY0MvKUqxDOeS/NOkk9x
ignapQ1jV1S99qAX7+nQbvu5FOkpfRpYOGW8F5lLZ/2KgMm8e9pWa66HZRRGho4NO0eBK4O+UGEH
1EvNs6rUt0XOc12vjh6Ts7ObJnrHiRAGyOomWjRHn4NZu0OYc2oknzIFPtC6Kd0VwiOq4RLXVpiu
DmeQmDcgA5SWpajnrS6IEcyVW3fdmu4hagILIt8HUik/jxCt1fKrNfHtjU9z5uUmVzH39YJ/C3Q8
BQkuW6PjwDw7oRgGdhh7biOWxDWQM0ETLoYZUyURYeXlSxQc4fu2wIlZE0Knaa6u7ilmtdEtvKNB
pAuXUqHHVeH2fSbEPw7pxhLBKf0tT8ADwFubvbJefXsFntsYYxC13yKsGbFtRXU85CMbTTAOgzxV
3Rof307woEof61OW7GMgCLHvJdMg/NU68M1MFSsK0AkFy7VtMEq957icNLDrfVhhEFhIlknbuVNF
Drvu3LVtshZTIctxyR82VHJeQsIawHDnVDvnoTkw2GfHW+XZ51+Ai00UghmIe81RLDXdzHqz12rj
tCynrE+6cuLkZud/uUbUzBCLtGKoJUH5zqbfiLM1HJB4P/gtbinKmEryd7lQp0VusFaM31XeI1PI
OKhBZsMQkdyBhsYgEO3v7oGINGnX2YZrFuYT9FNCkW8yyzkJNsXJJW7zq3zvM51GoqdsC869hUkd
0hKKVKOpV8ym+oBZt5rPQ2Loyp4erZmNTghso5Hsppk8+2vUITQZqZ4goqQVgIvY3C6wzdd5R4Px
HwOP8ZqfJqVkTliM3Io1kwIxXUst+iBdtHdjxtucZxwXi7m/TwZAbMQR7XPNn+Azl2f5wIVXZp1F
VCzn8uKwfSA+mVGQzWo16zQ9vejV9lU1YogS/cUcU89ZywGBTNpm7UwfxoSptUDFc1J5/WzkRD3Q
13Z6fP0Dh05xGRmUhn9BE5wcy/+gmSQBhuAT37yf2Am6zYKxWPjkuB8o4syPkZC0AxeCxhb7gJXk
TL+yPDoBj4S2Mpef4+wfHuaQkNKnrafia2jLGnnhp+LCeg7E/tQ+oYHXq7ohXqRLhS1zzpQ+ndY2
KbIoplUxuZEp4ADCZijvE2Sk0CzOI1CgjoZ2euFqcN/UG9ytP4T0J7NArY7xsUMz0X7c9u1sc32H
JCuMO8nWXyfor28lyB4oXRK3kaQz8ek/LMthCLa1srMXJTr0sjzNshcYuuTqkgZRO9XQB2hKRTM/
QWfW3DM8VrTz6sT6Ka4rNTyyzdJBzGju4ZMV+FX9EIkmNEN/7CckbIUVWJmaGxRMc3Px78Z5Paaf
HXaoR9bQtvLxF8I4hDXMXBdO9vF05nAyCBXkkLlYHwH06N3jy5YAKxTB6FANcFKyVjJaoE1HnleJ
TDWZD5a1YTBsPfAB02iH7Leqz5gj0Y0uoTYDfwKkqp9iBkeSY2YccmzyDJy8/vbTC0DW/j6cbsTa
tn7hUARSTPg6jDknXnwC9McomWxnL32WvoK3hZaCADr7JnFkNjwCbeywg4BdOZYDUtvYvbft5Fte
sZqBd02nEmyDhIlSBfszRvrjKrsLrKKBuVdb05ounFitY+7HXdF/kLNqtUOGwrw0YybK+loY0pWx
NjG8k6jTont1DMqUe28iDYjyiXwbV/TrXd6EWZ1alJUyeoY71uMiM1D95Cd3fhIG81r8R0pkh3LC
8mgJ9acKHR1kXXmmEY/1nEkmqYWZ++LDszFrsQXfTLM/KfD7hyuHu1Pnma1zuCJh1Ida8gGRul/O
ve3v9kglcnX57lCgtsvWNdJy0IZZCv0LMkdJUe0nBriEkAEHz9wBGcqnrUH/juDUZZf/QLCQbvGQ
rLbkX6cttNihe2vNPxujZm5wuP/JRYjQT565rETUjlvl7p7xtoZh2baeieCn6AfXxvjqLfm3A8R2
N4TC7OPm9eYcGH0ahQ4v42YbPBSGuCbZYdj17ymOpQNdT4sWrnh+ZUdJX3k7b3b8jsliPh1Dm9La
Tx3IvPg6A/P07o0z0vqt7I6mjbl7MG4lB6Leo3xc21fh1gP4ipEnUHuZIeNW1FLduPHpUt1D6h6k
UbDCPKooFJtYkZNQUygxCdX4goi1du7rvVPF0lflUuHbx6i3z8hm+5jdESz1X/wA02WKNylLoxh2
0wf3EzvWVm1QXpWWk4286qXpd07ijbvHfcVPwfueJrPbTrAuVSDgk7OCERT4oclkY3mZD2yUMSpL
ejxTtII7cEVoEvWoQNL70P8j22amx1oKoJFmU+xGLukQoHjI5BYWRoYqT4ujK2eTVGOjW/lDQUGv
r37/0V5+Jy08ysLUhXagjQQMEE8U2e4WRigOUqQvM7e1y6R2vvDqb29RhT9pGsxWWQSk2DcxUCoY
4+rA0NMQ/O16VPon5n69l78vxlDMXL3ldlLgdauVDI+lCmNBo82rHunXllNVksyQ/TRA7NhsSkXM
QgRxxr6kE5me+lVPJeyNVyiknSXKSg7u0/Qd83vqDd6kV0cLhoCsk/7tjAbrXXkx7EUKNeREzcQC
sEonMqBnmY4YExD8P4j5I+p/UMGExfZRdP8h+5uWSUDHrITI9QEefOODeu1YiM/+mXJ1kmje4zwO
XU0fxj6SbqaVHWYhRIowUbdeJWT8jwokQ9LFMtrw56msFKtCcxzSa4ccJoCBLImic6e7UFWAkCzs
nby6BM8FJwyliym1bqn7M0+uBozaRXQYLtj+FiBd7nOyKtebQGPOvxdn6wp5lNemnG1DJnZx14nZ
9X/VrWz/0LMnHFuMU1BKJJDaiQLXZOmv9RfCKDLCSdXmlGtrNe6p3CHoVA4vNkwXXjywkZugEbZa
HiVqFfuUNGEIe9IzhGH+EUp9LoGS3pJN/+9vTlXjSPhGKV0IrWwghN0GPnWFUx7nAP7cRvDXIu80
9/Tc+wrgI3VVyUb/jl+1L3GpoM4QY64wKy3/9B8FrhmBQ3jKam3oRaqAy4LdU5iQ/6JdXSeCygOM
SWpqOQXm9+0ovyTvm5lLBOdtUzEBHuVtg7T6iPpI0lDf8MnI9mysntafk4ehyxafcUu3V3ZYaCoS
VUZVClcWmsml56wkcwu2zpPX+RYLzYFwGVEAIZ391eFiBw1WnamEY9sm9cyIhwMM2qF8VRNaS8bL
l3wyUgnH/0r3Ncojm61TiQRdV8VidQzJnd6g9tMqfDtF4z9SHIn/5B3kXxmhclEXn8DkCaUJXB3P
NSJoGJenfzIBaGNPw8Tm6iF4/wwEi6nJzUtYSI4b16/Q/8Rr0PMbH9aD41+sqVmtFYLe5rOj0vsa
2FK5idT4EfdMStvjXE1Y7e5+IkMJUlUDiBHIetC1pDwg+mE60S66KElPR2cGxpa0WHS64v/i3+VW
X8NYnwxDSrSrS5JK/NQQNtTdL8Y2YaYiVZOvxJBHsEr7xpOasbjlSZ0UIgu3hGL6Ju/zG1ko2/Vm
fYQDfdLvAVtyLGw/SOSAShBd7h72Qo1K4L3r2OLlPdR4hSohTgPTjn6ljpG1yJqais7T7tL4KMzC
b0pC9FPPgtZJ2uMvCyEjfJrJ5CUfZCuWjIH1iH26oCeCTSWR3rpOf+tjDOGxGw5E/l3+2LyvewWN
/fqkDXzXdZDBRrl48GGiyszVqV4gVPvO8hkHPFWxjZQdCQXzjC5DMqnAsOWpY7i4Mg6Pa/DSGKHV
gIpbjD5YNNhOemvCe5GTp4TjLAr30p0XvEJxOU2xm11eiwjLR38sdmInPcrvTqrbCrJ9KDyntsm9
AUe4xkJVyHCl6NatlIXYuUo09uNzxX/Pdo9C6/BaqcSMW4n2oVhPX6JDpQ+Hj0WDAc6yviICxzvP
qkgKwwIRaD7vk/a+04KxYkdkmMkqY3t4btEhCxvE6bQbCUnpCa2TKr/WY++AEGjwkdgQxJ+LPUg8
wB2nEszxmuW6GEj6sMiHFlkVQKTUAg3/2b2pEojFOF41NhxL67xsf92484jESuDrpV4l72unoqVK
9w3Yn1JBnBjCNJExEc8XFRbNqBzqEft2LvNqLKxyHGNjX0YxxTQVEtJNyDhvVTr0IOpZuLn4Ir1/
RFxuBG4EFvwzuupJ78pBvyoJgvOlTTbihSQSxq6TR2BZTEOw5bSpsQu8yBzDtysBI/wjjWTvgr0m
O0KadrVJnb8qjafCcg4PoWID0LR3oTHzM4TbztaFLIDPegQ+IsnAuiUZflDi2paGKKsngFTFjBBt
jawCT8V+cq9/6cRDMttoNeLp2QfwyvbAZ22x0h/IuAPk2zI4E3bTIj3b7d3QdSGiQvarqAGU2rGX
NZ9gymHikwVl7hIQncFeMui6nY+oy7dqXG91G7aL/UVrENkptscFiJJzjN1VWuWTAMhPVk2vbQmh
09snVGEH0O9ZltcmxlxyKQMYq7gMjK//dmu4oku/tPLbN8B6XeeKtzrtKLNMfPYdkmh1XtGBlsru
rIEk1PMvwUGK6zO1gn4m2meMklIvTTv/pIDdD8zK7KiMEKpl53HI0oTo9H5YIoO+94wO2y1Tah+Q
lcqhzB7x9kkMBi8R2w+r/Uxx80o22qCyEvf/BOadoDT4oGSn5fcZqaZg3eAjiN7Cg2GfgjmHiVxd
9aN2UkH7ak7EpmyRo92cTRN+lsq5L/v+bIeJUc4EJrVcVuRYILQxzVdZX7W+c1VYWcg2FMa8d2oE
ace3Q11q/2SsjaBX25Uqb4D2W3RaesL6PLVPn95x8o3LW4yqZZcAmc2qFXp0ai4wm+uea4Eql+G+
KjNERipG82iWbaBc90pxaPgpg+01XRi2Okp+9avhEqYiwKT+753SlyawQ8jM1iHVn903YUmR7Lvl
bQC9yTDeUBWCU/jCc56tY0HRg+vlFhvR0FVht/GUOZDmk0QogpFVlVplgiu1mxPE7jrS+sGTXZue
khls2iQunwOPXooHxwEkVeXXL3mu1fZIe4OIKbJ0S53ZCcJQN6LZwNMl8zEHsGvUeuXLqjmBbNDI
Xgk97fpsF72NUqjURUPNsabqaaNkHj1G4ZSFyFtrLAX+cGIeAIsewnmFPwnrgUq//vGXhzoMxzDw
T5MM8n2Lu/eSefpPuni/zFrIfyQTyldowiR4xLJp4GfkDB0qUDeAUJYfV8lv0OAJ1VBkbw7Fjtsf
Y3lZB1w1YBh9OCczF+Ylium1cXpacfO0N8Aid8LoDYGNDM7UaHSXNciVvDsE9u8dbQZFWxke0ySk
Kx9LFLlobuduMuwRn4M+GLWJVzylhcCQ3BRS6J8egijMWUqxUj4e+3hKfex/Xkte+aLn1lrKpdjp
6EJrJA+HyF3L6NN4Qt27knw5XEQUqnsdRzEe69vzzOko9C6V9WtVWjzcKudMdRnRHL3J1/N72+qK
/fYWjB+iDeEp8svu1BRq3zet2E14yizkqwaf//t613FkWKM33+HArjW4qnfK2tFKxEuyB7c78Upu
XFaDmkhgz1s1DBMmW0xZ20auFw/cPA647EmR5b8ocp8cXaw7yVuJL6oy96M8qZ+LwMiBfUaPlQ3C
UxeR1fesBLuEuqSaQLUBRGb6wynd7IPXxwFIJRAZCjJvO8LzQNAPAD/Jpxcbof8uUBCynwKziPW2
gd0/o8NBmM7QdK2p0lxx4xB4NifyXPEj8YYEQTWXyUZK3o/ziasw7kSgNF/cOqphukYTxCnZRecE
TyT8AQgB2kg6krkEej6r6pTdF11hh8fqjheACDsJkfRP2MCu0erlHK932/0rCwls+shHXVefl3Xb
wFWPj/TZB+e1lTv1gTktSf5tS5ledoqyaMe1+/csQvY5TvG4hvt26mviNAhrFqhrHtJ9S+BcaNV6
kFsmMJweDJdvNkdWA9b7mqS6PPilWi+0+P8SsSOk1mXuziuiV/psgDYpkRlDXfYm18Fjbyse262D
Jz+DxRvW4elXa1Ts6KuFQbdHFdZxGNcj750B3KdiEp4o2IxJTavPI/R2Qt+ApZsba6tO4WpNy/qD
ehwufTcCYcBTWvjC7Jl2n9uhjjN1sANN8vTDIRfr/MJtpCKsqtYQZMyEFhpMGPPBlte2Y+qAZKYH
72ET16L9vKiWDBgfhbSH3/uUE4yRJ3wtdnXDP+Bgf6OWdjXoKm/qgFb6S/LTa8i149O9UKcy2GOD
69YC3CmT6lSNrJK/5X0C7+guulbyv19rKDSSs0ghLLNOz3w4gQyq5qdBGojnkNMGPy7PZ4L9Qf38
5OLlIp/kvqq/3B4aE+NPmzeQ9GFpJQk2EpNzBzNfc1Hafqp9+UOS7I9C/7rdsTyuGD2F4hKgtus1
1iq6BJvZM4yUPqU7Qj0nmBJQtYTWuTffQpLUomvIgc2A18479yGqjyxQaT3HbM/z/UizNuaZ5ESm
iqaZZfLXpeQw3MRLIypSUFVXq/kvNUlhlXJEADNh6spwO7CiRPX56HjLjmiHMaCjVJ5ML6EBHhBi
EH9w0aA8bAJRU/kHvPBBJqaUq8EL9xEp3/AR8v/Bdo7joqCaeLIRMxBvwt0OGaWeQO1XmcN34e7t
YyCQP0fa90ULjYnSJlDwEBg/sUp87Zl4PJgKTA44e8hxjtWVzzK04Sjw4/Dw5KC0WwECjjeinXx7
36WzrNbFplm2pgN9vWfZZBEmFyNI2+YeErq3sWZrqB+iuMwIqrDZnbI0ZCr6E+mHS9d3x9JtL60C
58c0ZXOgdnVMFaHzwXxDCLgp3lvCHGfOH52rgM/5K0slw967qXRMP0uzi12Q1Cg8x2JhhyrYLtxo
UdOTWwezuK/ksNLChgvg6GDE7HNWskcVB8TRev2/8HYpQxXLbqPeN3Nwxg3ZLN8LtZuQqIWRaCW3
+deEPUsj+65QJvFl2/2T+U1NitWY2LoqRjgCDh7kMOqZYP8IXv7UaZvybcAIf6wa+MQNkQCmqvVQ
nFJlozFYZ3/yY94iuHzQaNUI99laCjsm3BSZQrfOvu4+BPKkEmcALsPco+d8Je/uvTRzaDYuC8G7
Mt7jzLqlrea44BbsD+y9pEgPZ0omiYRvaQI/D0YS/VeL8r+oSexWBqmJiuhGCtah2M85K3FjdvSd
uPlU+HzafqCxoaQkPE5GQ29hb6BDZfDxTdFU8RxGORKW30j8d7ZkOREayN4qICCh1/SSaQdNg4El
BqJvo9vMSDNFuvQPPoafwVLiVknIuW6dNRQhL94wsyHNNrYLhKexZflgmi22/CcJE+KwfoBnvqZL
RldSX4TiPQkrGijv4smOzYbu+3WZCTCFtlKcasUCnQJb8aDgv94iYYV+T9Ym8f3Dxgi8i1wf3gsW
oH3wUCNNYmiGISADpS1DzYQDR9E/I8jA1WLinUp65Mr0MdLtjkOSlPCLEozKc21GIexBoEdbNKlI
qrEzOL+CWI7sFChclny5oqXe89nvRfJrsxOh3O4/xHSAeD17v+1rkuuuxVvPvSLitSVlxq4Jo3SR
ad5gpVjqJAjzvd3V+pHeEWuX241416Hk+syFEC5shJzvrv1E7rc3m0LeAWZbupkT+hqlJmos8VXg
VKBS3ZLb5fizsK3CU7cmZlNb5bwpFRhma6zIdfWAre3IPuqpbgQzHVRQfjOhSvXIri4lsbNf/D6Z
ovPuq9j2bdMHQ7wUxVR/lRrIXyP4/RRpUBt6KameeRZeZKYDAibH/UeJjXHbYyiSFbMTM4kxu1rN
b/Ek4zNTTbygAmcOh1nJB6yi2neNEi8jkGDU/aQw/Ti4KXyZcgbQ3mQCVnSBzuyfPZ5gfYtPfA5Z
nRTNE6B4Tr+mZdAlF70KGs8sMC+fvxopm7I+vAaycYD3m3nBh75+rIm7Rs4QAySyvRGxK8PCGtgk
2OOhXp40DjJQ67JYRdufff16g6gFJ2xjQ5K7CPwBXiFdgP7GITBZlavNvsVg/KBOYsTQd7ejKXzs
5uxVzCdINEydY3SBXUKA8NFiMZ6ffvy84ouAdAMj4dwPjYRL8o5wrih8wQ8qXQVUgh/9h+PsNNjV
MBAbtbEhVAzPtHKZBZazuTRU9rN9SHskdUHJG27MWohU4KY5Jqq0FKcQEOlelDavLmhK/GwTPBHi
7VlrunGwZfco8u0+WeRLWxTh7VMJO4WI7kTBa3U23SruOCqB8lQvTbnWHIMgmB3AwqfLDaifWGUn
CJGvUtQGctTW4J9YzgeYPNdw4mvNd8N5QqcC9mhI2KssCmA3OuiTnAhs7/fcTx/tsyNwqZKov2iV
t4gdVON85fsXh473s8VXp2V0fa/OqljkdwOdqkMzaK81l+8yJjUsT63aQsZEw51HWe6VcEsmhuSG
ptaXEnJhrqdAqOjN0FKwNh0rzPPdGNEV0ZWlHiYzAQe4+XLpjUGJi2qWlygCjM7GK7ohbEgjTZBw
0717l4YoEa4hYfSKxOGovAiT5zS5m/0VYXgIe8tbmtDIBo/xE1j4NuH9pHEFiAQ0LdrjK6umYGrj
CTD3QQg9z2/cRiQ/Jay84PQ7xo6WecJEGOGWeDkGIr+E2bF0J6eqJNg9V1WE6zaPFFWD/WsSILsj
xLF0gnwoVMBrkK1nMwLGvxYlDKAnDVC7L+lDWUN3Jn/igP0B6lbu0cpTl4W2KMssheyo1RtvgvV5
kBoSUXyd7go7jmoqlAhJ/ABtMosYwBiGb6C9v18IN5d+zwH/bQcL2RV4ou1q3pAjpXE2jPO9CiSx
AM3NZC9ZrmSxBjVkmjnwZfs+uwfX0dHDvMqbH85VOH1AG/dTTvXMWZyHwH+hk6JyWw8yW/5ahi9S
YeBe2nqjrBlKkaFrpO9tlYWB9JEkSNtPSjzHiMwfctwwTjzTMfKK8Chv40B+NWZyLNzVYggAlm6X
v3iI6Auwg3LcYbPJ6RToyoPbZyp7oKrGoAAkjrWBSoFpSqbwAxJByXzByQKbSudUTVIfIzpZFD31
xjieY27Pq2ZAYxF/80GNj2l3xNt8swehoKfhtg+HmLYMVUlL4SlOJRTLZaIiKBbW2sn7lFSx8/iA
6L129w4KDrOJ8p+oVgLN+kj8BN8kaLPMi7f2ndqPAaMZsEP7HF16bY41pSO+KoPdxmqmr/D8fxvq
w3KfaRAF6J4SGsAR5+vlW0WdS/Idj7lyuMCVNfVknLHO13VHAH91Ssbgwljpq1OuUrhdn3EHhI5Q
BJ5W7573HMjE6SrX4XeUFQhb9Qe/U6crjoOzWzKnZJgtpt6n+Vk78xWiuWPmA5nj9r/oUuMpRczv
+8Q1V2eE/gbc+WZ5ujZXJK/pUnHC9vG/gMj3vUT8WqTrwu2DF3Wd2OXS/qThYCoC22VBJ/AW3C2V
5qcGOJc2OCzlX/bI0Ix2Cg5e0DqcdJoX2Qzp8GEr8D3motIfTaReEuMUcvT+oFx9Ku00CT0Zjq3/
1qei7kVVOal+40P8uDGL0UjdqOSm0oghDZOAtPIQ+7MBc3gIkK3TjS6yPkoCtk1Csznac9GVRnTH
74FI8JglnTA5ASfk4sSUFdenTrzzcwhEYhxZrd1mTZOUu8s3e4nVQntlZnQFTETlFFD9RxJtqqyX
rJOgfApo7VynGRvHC5c4uF+FuJzrHI+oxnqnKCE1M+ozl4SBfGTBRd+V1HfW3pxQ7dR+gdw2YYzU
/pYjq1PhtMFAR3+sVpfSK17i+qkOC2xzPBbuXvf3zQifVyU5tTvhYlGZNng4w8iNXwJ7A9doHwlo
nB5sEyxPPHY00pXXo3OTswDRqDdxCuFOZlNO7gOoKPGkL11lM+HLEv/dyETTymTKTIWQ5F0awabw
ATNGX4vXYmvFFsGoUGoiHICrJFVseWlHOxKlPmoCjNwuQtqLJ7MnnngsGC1cgx53eeDND8DlX7tA
8JXcDFNh0UOuepXP2ijlC6OTDPc1DwpQiShsorIk/9xvAbg50P+boR7kihbuON4YoxHaQdOsGiB3
9JUzRWhPcSlZgNaAJA1RC/xvR+39jK7GNMb63ILIpa5a9pJuYYDqXSHdenh0coodQFQsQ+J45Db6
pm0phfSX0KM73TVk9KOEeSIWVBg1Jt7O4gxr3bAWp1+3u17eb0LnpRec4kNXgYxzI1nOdg/exvY5
+whV4be1zxXuqGk4+8qiu1pzeWnHrdE0veWByHIvyR6pMApL/xBK7LijdmwOGt3qv/VdvW8aSmtQ
/TJDTee5VZ7Xef1lZSXjetg0IYwjwY+KqBYAbwT8B0ReC5G+BB0dEbPJIRTMmw1LAtRgk8k+a5zv
s/XxxU9ZZY9zdz66SYxzLL5fAEMf3xwJT0Wvtj70ToxTkIa6M2FNX2zJ4QLLSXtDGmgZ2wjPSCL6
wbT9sjlcN119jSoGmoMZlN2r+P+vCDDOX/ORJeoj9g9DklH79qRQHiPGLcx4G7N10UQ0jCTJ8+zd
48/UcjfeHeJW4rIVDfvvaQvCJJPCUCWFyTDJGY1lCXa3tKS6HEukC1Te4BzbamE3TfvDy2hwyOLr
9sqxcTSTXmdi0cXWUOOnVcwLktETAMvvlBycfltv7sD5qHW56aAR38iQ+zUX2jQ3L0rkKDVBvDl1
5qwWjf4nYekH6fSA2mPA+GfEdoz3q+lvNH1zzffsOy2DKLKz5WtkH3ffgcadHdzA0Jf3VAD27aDx
8rMio2ESJPBW2sFSZNDvfwUP1gPECgFdalqxm+kzBOFOVUJUgUd+mBVa/cbnhybsj4LKZdu5arQ0
7doq81oRmelvwayT/C7o4QYg61kyZ4j0VQrkD44049ajKWOw2tY98WshAJZnUvSYzbXqOPf90m1W
bo6V5Ir+ovMOnO1lU0R5hhSsgg1Jm4UsqTrYs9reesoUO+33Z7XNbLC3zrLyUlrFeZf6Z8WO2Jmg
g7ULJcSRWa1S4mquup9FDwyB2UuBx1VG8zZ3quoLkWbHM/ZrUa7bXGLJGmrC2GhH79+ubNJ1BGXM
+PMsrUpm/SNd5VRoJvcMEXJXynz+oOl3L6Go1JBXQ9XK6UTlfZIJhrQkGRDFftohlbWfCoN2W/or
dHyLtJLinrPqoKEB0cCZMVdjPXYFqjLwXw+LZeTPQ7rwflGMq1FXKEkXzmfJC9BM8BUgJnDacDGJ
BiwURIkgsDNMjTMu5hxGSTMPqa4ZUY/CAUQ0M4qAjMzBTwN24eSH6UxFavbmIb5Ux/c/5Ktopt3s
iwLcHr5yR64Y2Q8DRU9Ai+R8mV69wIC9QdEzwUcK4Cu29aD7VfvzNuIefvZ48ioIHKcsNyKcRbir
c+ecr5am5hKrZo1SYNPi8Oyuw3OC7UrRVON05sUuwh4MWwM2wVrWvPlnc3McnB3kufg5eSoHFTEt
uqfqyv+ccWueSv10GZvk/qy0vCsP1krxeb6/qUvO8nQAgK2bBHd/lGpw5xNYPEc7WAup+LS9Vk40
eIKsMNjPowmVeSNR6L2mcmbew2LtRNxd06q7GV1kC2bOb8EG9A21k81C3Zhn18R9wfs5UcTmL1dF
2y9F9Bxyy1v3kNg+O6M4sMo4lR49j7wKhAMxqeIWI72sKW4ayuYPURrttgp25kd3NGdzxKur19mL
gv2ET2f49ZCiabGqtdxcJjv0u2bgyX/Ydexx8bFxItf8Imo9kKhhJA/Jac+1DN3/t7H4UDDNmph3
RK/AaGqbuh4u2ezKmbpnNUEF1n1nzBa2ZlSWu3gRMeG5ZRqlegR5QnbhzT45aqd6VNreaxeP3NAc
GfR0r1BoGofFrVXXtWQ8up9MUZUrtK1ublKf8f6VOgyO+5ikijkX+gsWUUedps5o4hTS9OQHGT17
4gj7EkYey6Ul7v24w9NBnxsYML4hpKCQsj1EXUdzvHH2mTRLWKJhBrFvsN/4jBwxY+6RL2XuJBqm
Zlym1EAovQUwGzrxXvZoyqBaT5yP6TYv4x1ld1XIKpcV1z7I5iMiZk3mpcTeL1cCEccVWiZfXc5A
8LtK4t8pNEBrm+vPJ6u0sQlUGW0ffo+SzAV8V4EJWFgYqrDV/rSwRcbHsQyLt69UdQDpOIY4EMys
GywYqXut6Uz/oIcvYkrYl2sNMeN0sCUhJXJKVYzPlfneme54U7yXhYgPsI5UK+nrGNGUtptEwCQH
icy95Nx4aDCOb1nrVyj8xP0dn1XEOVapl2Wh9pn6zrbjaYh+D3/ndWD4Q62KxENsj8hObEKAAhWO
XViyl/PS2Hicgn+tjriRgmNsdAAeRyK39ChEQz1CBgffTcjzNospRyRFP8MjAEJVj2kiHnMxNn6+
q6Ohwi/im0LXOHODFiNacBMWaLXh6VHK3hIElrioUEq+3Bk0bFO6fQkFUm2JINhtlJOWnJpqVGUa
rg6CCqUw6pQ6yhqkvbRaik7q2OC7esxQEXpR7VzDrf9pvRdCjc1urix5ELBOoZf5FmvxK60bNgkz
AovbVTEJIvw929oQEPMB5pM6FvJHdQ1W9mqPFq5u96unwLwVrlxyGsaHDSSqEfFZtuXVCPdPohkR
tGOdhn36EJJjyEYJYdBsiqmK95dF+2sVjH4/nfuNzLIdM4Go9wVFtG+F0yi9vQKT3LJ298UsjjcF
ulkgYMABIQanJLKFkQ7+9W2/Io3kYvwVxnJ81YJKlPzUnfgfsnrFY7wLNbe+D5MqjDr1VXiWmogZ
t8m4kK3/WPNaSw362BrGMi6gNOO6Fq/jQ3zy23RW443X+opATeLJ6nEqTLxY/C+cJtUMFeMwLluN
+LHxoR7y3TaHlrFwEjr1xp8XwjaCzAKY4vUL7blO9w1z2b36PbDlhZV3grxztopBcMRMw59cKYhW
Gr/80HQbAEsBvKuZB/p244XeNJS8GZ+0oYdH3fESfww7nvXp0bViPlYixBwq2IMopSof9UATtqsN
Qnw4xSOV2w7KkdX28MiYU8dS7mGHzaYHGVs9HOSTKKtlyeOG0I6KjP5bHSzhtMw5UpxtGLPI6c4o
n4SY2jhbKuzI2GUpTJXSb27rmr921PXUAtcqiIzWqqzDFhftURJ7BjbjfY59vE7qWxntroEem6ni
68SBvgp4P2eVvpw0pVzQccwXynxCMqtMDlw16VHwPO0zk9UgnQ0GBeVo6EB1E46/IemQBkl2fS0X
YKrOIn9dKaT6SjF0iWdd6YXGl4uhkL+5ktvEw/qJo9oqs+FGoRmUghhSR0nL5qS/cCqY3QQZC9OR
+uGmRG6GZdJKL3DLn+MIqupzjUXM7b35YNUrrq6JhBItxw9IvqQYw9GJRvlb2mrroCXxP+sm042b
LC9+3iPbdzh6K9gUvKQkLdxGCkaO0YWLlCc3TZGi3c8EGa1/zi85TvwFNcdnChpopy8yimZ54gTt
YlHi2W20euZTjVtf+XbQpMSq6O0rZrtrTKkfm0xlxsIxINokiu3V+F+xOLjNID2bjbVCY1KTudHI
2EXlVT8m8DCXUczecHfRduuXeLIYg9DDBhy5Ehi0M1h+U28aWDScAxLGxaopayRoGPVfZqH4WraY
ef+BhavFynAwMhVItLPRVJ3NebXiVRh2SJeVaxI4DmJpc8YeZqGWq6Oqx3ObU8qFuYoDLp0LSSnW
Dkthd20bQKSA27z7virXRLj2tHWxUJrkQOAIvhFJCyTQtNHOsbW6WC0TPMVw8exFUFMUsI3KH+Nb
An0t5YDkwnfnpekHa23Fa1fO0tkXP5ImdCNoDzHRuc6yxUbtTLfGU/xhKnLadApcTP7VXWYVxA9B
1mmFH4BDg4l2BzrwXsgy4uYSZSiwFrL0CeW0+PNEmxc3o/Eeq7XPchQnNYYzsDcV2mOaD0xTCy/W
2kJ9D/EJIIQpklofSbFoU8B8KX1lKl0d2sW4h/QqC3PapQSoQ2K52TB5O3AP80B3wIIyaI3FH9lQ
awmWK7h8ZOlelwCZR+tszBQZQu26tHzBWRiKAYtMBr7ARMmnOoh5TQeeTGm1sbooHVAchLnTkaC4
4fu4N2MQ3JKXndfW2mmb/QNjpHIH9DmUGMOXtpGhDuWEqiyqiYyJkJRK53Gq2iduVVpP/0EXU5wb
yy9x8H4rohdb5yaaFj7zp13jm1ysl9nKqTphVrw1UC/mI2AFu7wcU93yCszGCkHYSqAQ0Eq+RkNu
zTr2m1nB385ULDYwQQYcIeQNpVpbzBmIbKJ61M0cpfLj9lHzbSYmsWeoR6l8lInWWseBKUqNT5rn
AYlOOQhWqnDG7UktbuRq3xULDfEKDXt1IUkevO4N5/KwmfdTU80EyGr+/8Pzm+z2Ny04H8WeuqHA
c7XqqhSobZmt7ve7u9zoeE6KTLaP42vTMsECGYNN4hAnAJEPn70hWbRsQDqId9yoPiLph6YdEUyF
ZoGWjxPHUbQnN6XaONVma/P1OTMeBSdkCRV9xUpCa1rO9gMOTdqT8RM2qlyyX60jg8zcMlbn6cMB
60HOqxXitnBDR/b9OtUnIHUcB3EB+xyLoPzwb0dVWimkbT+gi0dObIQ9buoq8knIBlTwr3hCPf/5
Xrcyu9N6KXuQM+eZgF22Ql6rRBmpLrKGSpSFHcJ5ZEB8kqmvsh5rrVt6NhaBaooMSWmSrGQHpL9M
fiGfJ6dJcWkexAvisq3Et07e9P+KOJTw9Z0UQCOuswiKxSe3Bdw97NbnSRxIt++VLU/v/Ifsd7jO
yix9Mp5gWp0tFMGHDgAYUJXw4yyZFTCB8tJb4mH3+GGU50O8Apu4HtoBFh2zolyH3riSeXg1NPGr
id2oKWno4Cy6xXR272HrOVBxnaKG5FNxT9+bdG4xrgL0IDCvs6IsByVWy4jdrARMnGJLvfLnMxkJ
rFiZT/Ce+O35fOVGb2yxPUP2VPti9+HYIA7hBjpvnT30MBz91/1DaQAePgeR+3txwsmesIipXXFp
PtNJKnDig+Y7HU/Lm47udws2p7x4DkHpNi9fZ3Nf/fVd8RL75ui5nbbA9PfxzOYCCYRNT5ZI72mW
tpPVMiMsVhmJ2j4tMxb/xX81W8RwFMn4jNuX8wBMjPPIYVI8xrVO6WYq8bPmJ7Gg+P+7xH/w520P
A+69kglyf/BfVsnRE4ssgeLNuMUgxZLroiEvOgRNWL4Ga5Ze5FA8mfcXX2Xj14XA8wXY3dbtGZ1q
TXUM8GBQvR22WFNCyoCClLwBB+I4d2Pn6J7v5LqdlkenpnIkvvLxOLXjsagIHBxbf+zLNUAoFGi5
F3F80RhhZyG/zR3zOQSHGQRaCwpFvEUW+kcOdnvTPK+vtIg4PS6P0q7GGOksMM9exsJRXEzHLsIm
MFPCIXn1Gn13lMvZb6ZNB0y1CAWhI0AKY4oYBcV5aaVDo8cEGTm1J30ikdUeJmv4xS3LdHpLfolT
dT3i5hMMBsPrtdTKZk+YV93gqt4ImmBACUaXkP58IzndGKzae8V72B5yLivSnB/99DtiYvF88NGc
whVWHSSr0dXF/8HOa+Mmk7GzVM5wjGQZrrjaroR2H4Zof1LCcGn0+OFhBTyKEvGtAfUmeewmUy4s
+iUu6ZFF1iJMcGZNWs4XTdq3Xk/RCWSIXVQI4LsoCkYexybjkLAQTw2qTChV5cg3X4QNVloewrwx
SOXXFnC7VH2Sa4SM06jPIUBIuL3kYovShC4IvLCjTzsqiBkj6b2DtK3vsbKE2HhLLQTrVNjtdjBN
V5SjteWTqrXM1KjCKYxChUJR2yQYfyKQ9dLDeOycLEJhj7MIyNmuavWCTNk713ENHOzCmpXFJiy4
p1Q86timuZJbs6+fE8LXRw+C6Vj5Va2tUQlqpqpMDD98dHwzHZW37m/y0tkDDh7O59yu8BCbfMaY
veHpvT/N1eII4MM9BnSHMNa2o8U+GBT9zyh3+X9D0tNcOOZnJdSg+6S6biUg6wdXteqdIUs9lAk3
BP6Qo6wH+mLCzmHveKIyJYPh4O5VQI9buLsOeBK3SFw53SW5aHJjCX1whI0sAFAGUdtkWDUYsGQ6
++CQRSwp1qZ9Issbv/+ucc/Djeze6L7H0JXab1ltr7ACXl2qqONZ/URHZTIHqzVXZx3fWawzn53X
Cw8KjO2XZSiIh2pt0nAxjbTtAGsx8hRgnrGJvmefXcyhPpuWHNNoEl1oWzWaFXhbNuhWrwm/0NXn
8rooQbOsvNGK5ZynCZZ4gHOjCr5i12t6OKG8s08eFLBQ8er936NLYYe91Si2qVdsKBjcuLmd4nEc
Vctrl977FhDiiABG7N84E4QDk/UG0zzinrv9O/rB5LKY6Ss7OSQY/LW5gjNulZ3aC87Q7wsR50P2
pnNrGVgiC3rKhn6s0BYL9ML6mKs5IaL+CQJsE52FbqAKPlR44xP9/lBxrrTqIKqZ31rFD67uPU0z
tD9PihedWlcPOn9wmxWcfpcnuiJJZCqa2JNCkDUsRDLSRWhUul68RlslAGkNkVZNi149yCv/nNAp
lRq+XrNQGD0/CKvzjtYI7mS6J3eylbqF0xlVgVzliXqxAQ5bRRLHDPBmephzNSLJLOS/Puk6wAPd
/g40+1xxrXul+hyZLNnrnoUaqTtYG7LHWPPgtgT5jrSfNtPWOaQ1c7rYz9G+/DaCCzr2CaXIpYqg
CZuUIgjZTx/YBVzpB0SyotsOaszTuxykpTS5B7EnR/tqYaxheWkmveszhpOYCzaJCRn/gxXAKHhz
TOdEhS5kmYCBp39hoyMAyA9yBTgNnv41R8s9UQy6xjyXxA9FcE8imFTF35zHKOPseqbAwm1ky2ta
qX/+7sVeF+xkU/LneB8LMk51z5eIpb3TC0KBvOnV1fxYE7RAtMTptiJO+QBkORTqa0Klp2MZJbKk
7R8zwNIn1i/B0EZ7CHRKfFV1p/aERAUmq2DQaUw86fLirvUDwW/sFlvQFN75UNdsdxMke5HEzwJw
Qzx+gyHpuhTg0A/gj4207ASW5nNU/Me3FIc7fCOTrJDZiaNRh8VMj235t5aiEsJAVtShi6DqUUMZ
VfdbDbGxMLri1X4u8p6wIBH71RHoRdeP1aw5y99gOuugd98hzV40ciNVVeKkYMAzSWp/AhAj9KRh
vk/c6U3nQh2D/dQxCLFm7LK5T8D2ue7ugw8zmbQKSl9vlNLziiQ6MjiliJHD1XjlfZHB12wab2dX
AYvrUTsl8LXOdGt+4ISmouHIJBfTwQl2jksNnco1mPJqc7XwvZHRbKjYg2MA+o0kjaTO5GJmWCRd
YePp4FdjofXPjX6013YjuGvEccHr1vXP1Mnho8fV92/OGwRbwsda3QBRxwRBWNhX2PrHqGdKCPWd
wcnSh1QWolVbO6bavxoJedRdn0IRA2juV2fiYgvYb7fxUeRuwXoqGNLe2NMLWBQXiWV4kiTqrp0w
9z5Thvrx6ijHQqLsdoiy5lAO4qbiYjNiD5z3K+plPBeKjoKDB3aO/Dx9kIE3Uhce7nBt3e5KmhkZ
vD4V++kABkWtjlL1vJ4M9n2bKERqymkibJLZ9PjfSFvSzib6oLZ6iRxvaWwos4GSwYCkYTPrbYYg
hqo3PEJPPg7JvnUK2zTGpe13WbQylmOry8nWS70yNkiHvaXEOlsKOpcI429ChbOPRIUQSHIWKh3s
bb5B6hmUM7mtXpBAYRHJNakI+K7nU/3N6vB/fWuwwBCBPoWK8NezwALnr+eoP2EKDV/C9yXmfHwr
lmWDh+7OkDKRYlepHZAIsg1NMRzY9/upU2c6nhriqSHaBZZFGWH9X2/beYzt7C0OE20cZlf9rn0y
uQcjzO+xj93Fe3di8odlu76v7jsI57e/16HsrjnW/M6FwqRkN7w96s23ZP+gmYJtO7fEpEv2zc+L
puBXkkhT1bOoXkWBQ01kh/akAw7DWQVogVnNghHow9AoszwJq8phgT3Tpn0YbbWL3lTVBZYyHdvd
sk+UNpz4qATWSV3/QZCSIy5nvnhfHa5mSLK0EyDO9eWo8nbDgkknBmm0AuCfir7Xf7+UzPIV/SIn
R+b7tkiMKX/8ai6j54rWQeb41tkI6Pau3sIMy6LAGjEpdch+glM09mpw8WRF2W3qiEMP0TFwNU46
A3MeLUukHPWokHizWywkNWVrSGGQw4cHBtzZY7Ytahaj91j00qAI7WMMyMlvFSJ2ZlCFGoH555IN
zbkrxbk+LApqPO4+qVC3l1BRHJaQTcrom6b9q5pKc/awlpeK3EvawFtl7mBQtPrK1tF4ZV/3A9Ai
mHW2CgU49X/JcD1wiBvBiOO1v1eXO4DnqSCpqrHXUSyjynaZNYVoJOrkGmnq/lVP+Q61KYRelCAR
oXEijMxT+0vZl4wqQAEKyZySb3ilTC0NAtzBsxWjKOBTeKb+8kDutbOz5nn1qDDhG8a+0Io9dap7
6JZP0Hv+qPIveo46qJ5vV7lM17zePamllyPCmLyo0H01RnQPKCYpqjtikibr1mCcMXJVMZOQLRRJ
ElS2qA7f40YLG4Q0vf8pXhnsQ4Q8lH3lrHvp77if2TilHBNzO0UagM+EtjAG0wRxE7pdEQGp+OoV
ujnzLkU0X85dyK56rMSIZgmobe0SvRvyUvJu4tX3g6oGIGMNKWEr0lnCpN8B9w4UT6YnIsAuCmin
J13mrzfvfwayZhVzC2TzhWPJddKeqWiI3wWSyti71muFDsASxxGFuEm9RfnR0DZH9i7qy0cHrzGK
fW/2OUzvLzgA5Q2npSxJV1TaLuhkuqxXOiS8cBK49Xzv/PBVOOSXpSrglcOTUSZoh00irNlhodzN
qa+ZUfQEB/HkxvVR8pVIyaUjsCSwV6K+GPCie+M3jK2erYj3zWnzpbaBSqmEDRSLvXByizkh9mCG
8NWQUQsR0DFBnhrP8PMP7QhsCX3q70zWz2/rNOO+szalX9ReWQAWeyOsNN8WDmLTGYkGaDztm1cf
4F4ZTEyt4xNehHdWkw6XAOFQZHSRUkHCB1dqWHEv1lftT1ksdceP1yNzGlSVbaESKJdsdSHIc0M6
O/M+4dMNC++uGURUP5VxarS9ZDXbo9acPJzWPtUUrnLMNXjYRA1Sef8C3hL8zt5EW6rh/9vZK1Yk
K8f0Y4Cb86IH8JfdGBmCm1OlTNKIauOK80E8SgmAumxJe9BnziQGMe+aVWK7VRQ+3rq928cUhxJJ
Gj2+/5e4RMMHE8FsegQesaE5Su9Z6K0a3JtBkXGfWJXRBVCfr1QgM/cTT8fBWXoA+8SW8/mN0DPp
a6ZjAHeMa0lTXtPgiM1PQe9IqXesfZ70zkKz9lbPIs0O1cuoDtTVKH7h3/7pjMZJUtvaJ9i5rpeQ
0BpCfs7vZ4BdNW6tfW/BwGeUdqBxbQcPMfcfDWRTQnHWtcGEB3XIUi+1uUSA/erQ6Tzfd/EXNh1F
2ukOUOc9S0jIMrQf0KBi3PlCWSFujP8HYzrBKe7JZQimTX/ITTfXhoc1XiQuKXBw60MmK6OQc5JN
wggui/18Qdd0Y1N3qn0vNrwdPHgiHAufxXlvKM9qRpxUnegRrIJa3ti/8ueW9Kw2WaXBV5s3Bf6T
KZ1urQYpvIvjBSdfIbDHdc0UeQd6/mCbT7idgo6WYTqHb0NeLZWCcWoVjcjm+XP1ITp/231rgzNm
MmdHaZAdnyoB2k4Qbn6wxTmy1r72zeCVIF4lbjCZT0ZZmldR4MTYYOn5YLiBIWfjZzVpzmhEA2Fc
ZyzUZi6NmAyjaLy23uRuPFAbKctMviuZeISwOybZ6NHT9gcxFKtBJIjsQg43DCdzuRkeN3b3YI5X
lD/xr4d6dPr+RUOD5hnJ/jlUVGwhwQyyGnsMcM3XBHAy+X3NxWnt7lJMF9bcmdrnEO1m/sKrS7IZ
lmVUsZMh8KqaGjDmMlTgrHtz1HqU9s9gvIfll9WgKeibQrRb/dZ7NcJOoa/dhNpXCVrVrRRtRtKL
8n4ss/XI102PM9R2munQ55z+A57tUMzRCDCywLjZdtFSvZ36d3kdpvQOWZWgFPMSquKFwHdvW/uJ
wNBQ6i85iyAuTwR8y2KRkq5CgmLB6Fp1NrDoitaMq4uq1XgLzVg+g9mPjRsbL7ITWPkdE7t3vpY1
I5j5uQIqhj7ll911Xpsiu4/qFs3BYm7Jz/wo3xCpNttcIHSEZvpC8zalJz+YMX8IU7W0Qc+o8Wpe
vjU6pSAFIa7s7G8we5tb4PwUwNsy+Zta8F5rIZ7rYJb8/YvFcCZDHhCLJnef+7fqQtut88McPmJA
7SOU9g65hD1wEuw7/kWFDwM9v2kpbsQCw/24bo8mLnK/R1qGDgNOkc1/F1oisYj2jPRwVsFvWuyB
z0mJ5yL+ssIp5mr5SnQfhJpO0w0cTzPZHm2C0vUgrywYb1oSb9jYrAwX+CvR/wBLCzp1yEwt9IqF
Md8nr/dGGoLdztv5X7S2XRpKV5gi8PM9Gg7V/+kg0RRhY1+H7uFPR5oc0N7AO4fB++r3m0qpOEmv
D/W0Rlj1q1md5d93ZFrqQxJ7n2KtLV/gYpjmqsJrtJlAcZ2516eK0KfxJBOcxKYGmGE9SVXblqS0
CJi6rovsAByDqRAHqh3mEKyHbx2xr0IbxaJG6cJZhVv37ev37uRGgtWJCX8DxfEQnHXBGJao7E6c
LbuImwVu4QbiyWfJLyBydTpl0ZH67kd+8G5ELZd/C12wlai0yeE5+jZTd3GHJ69l9W5HLID73oxo
4cnB+4tjrDLJ0rLxtkel2PG0QFN0cAsWYPlHjoYPBGVQswi+/eU4pVmo81gSn1qMA1FdkXHVGSW8
bQPsf2iCY2pcK4sqYrkBQGbTbKK6Cv19BMF89esqcixOuTgPUxu01yq/dleH9G62wX3AZd0nbuWW
hdv02UDlaI0xkt2uYXdilsOoAsFGPd3aDlL0l25oVcWfWd0LjeADeZBgzSsVQSTnxWoTOkdKWQVo
J5L3WPrVlQv94zRW8mbu1YIAgJuVJbb7sKBuz+Ohxflg5bozi423/ufwuK9Iy9pEsax7snb+9wVC
LyjWlK7wikr+eurOkzlK8XXKwKhxx7jBFU43dp1XOmK2mcKbsUZ0mrvBqxiI15LBHIW73bbjTqst
7wdtWjEj5K5jIKV/8ihN7f/z6+LDGtyHqy1y8xHpLzPzGB8Jz5NeJpAeOtpCwkV14rxD9xbMwNu1
EpoymUt8tpJ+xnEjVHcxdmNzzgYq5suW2AHS14cxXhFksBojmDTxiJne6L4xn7Q1zXfZziZv0aPv
IhMwMaw8uGkU4B4etk0Ity6/jSoQM9rO8RQiSXgWoNctMhjY8Eq9EgcJHQIoaixiYIGmAs9EUQ9+
jC8eiYBHC2bsHbUSrbANcp0pVWslgzUYofIrtYqYGtzwL6xXbRkaJAMGhDpZj6YB9NwTfJ9pjC6+
WYobRdseB0tsGkGZrNjI33XehBsK/lwKOzooJZ/vSLe/LifqWo8ctcS+vx65akCqIa0Fc+J9wCKF
LlaDlqJMg3AMn1UTcPsXn80pyQ85KRdwRc+mYcHurtDlC+gVIgRzSaIUdPfMk1A8P1Ym0EAAmp5Z
TIk7i5xf+WKfb2840J3sounKb2FRsLrYhrGHdcBKUDOkMwsXowaW5h/DtqhgAtKrz+9xBCNfeBhJ
MWg3DitzocsJkswKhX7Bep1Y2cahl/0VRi2WIyEOUxYy9881HLPyGHukAAVj8elGkxHgH7lnblEK
jq/xnYJ31sABd6U0vuJMzapSwPDci7p8Igm1J1sGVat4e9iGJKROhh4KvC/O8Oi303TQXgs1y81m
cfVdcuka1melrYSRGgNQiTIByKsNkq9c8UVwwyxPjMwXgJHE9t1M47Pfp0j+2+NIKlGsFMaFQ9BL
p9j/chGmGNM/1TgOFv2bojuSbOhSDY7iyCN4hS4eIh+m5obbiSMrI3Ib1WrZo6npiMjvtLywZDYR
OqICF3VzJun0zXUZ5EFk3ydOsoCUHuTZYgK+9btfi7xdWkLcEnoFlE9QmHguraSyAq+kcdhwcS8w
dLYVrE054y3VRYQIWk8OnZ0AlcLXB/iedVJZa9nwI/yG4P1LwRQiilwJTPanXys+eVB18ZEBx6ft
BxSeR89zn5xVPZCQJRC2vnqKuMrKWrIQp1Te8LZEFYO8BtOrizkG3156tMVo3IS7kAGhwOGT/VuV
Ob00t8KDmjzgtyT23onSkg9xRG1Lctk2zLCZOwxvehyYdC9x6Dz47ShvFXj06Oa7jGJo2o8x+HbF
6LjFOuGdb3K/HueQxVxSiU+QNvJlOy9j5G/Gg8yZn9mLxcV2oftnvhU/hePHGVZI8iubWglYstHo
2F/BKSm/QyfOATW/PPqpEW7Getm34mSb3GKtrPyw03kVk5EBMmOdSenGpCIY1LnES+mYNFaZAozF
+WA522Co7VOUrYbF1CDUCDrH0yZeqOz/IJMzBjKzrphhUCccPnAMYDLe4o7844R1cC+vVNtZGAdG
T83+5yncXfRtc8EL200c2DPGEko4l0NEUAP8A8W6YbD4TRjTpv2CxE0xwcdE+M62gjgxMUp066Yf
K5NCjdLsBjIfnsbjp6wOHfSwMuIfj0sNrkZpHKVlmdxXyhmKqX+MJmL2AR3q0nspPRF9YXfxysv7
BapV90HNCz1+hRWdn84rbanufU3TQf8K28Ynty8iU1X1gcSuucIiguNwyW0mRieUYdt2yM1FIz2w
WhHljoH8XA1rakkrDZY3D9mA3D0hcBwdHVQnyqdpZCUIztoIQdVtfzWvqZiymCGrt6FIb9KJcT27
u/Ksq19By8guEAVcHHfmOpNF07afPVj8gnEsBjxA4oYuA6xdSzvDPnoL6VtTfNHVW3S4HQVr82hn
Mu9FUktQModMfdRDlMX0BS6vXg2qXGuUpAHg43/wjCjm7Z3VphFhFC5vH/c70gUw2v2ByCryk1Es
po6mpsh8iIaJvhjyCiJgRQNJD/+wArKZC4LBiewGZInIwVBKStUUfFolNG9AZveFUhI0BXuyo5bm
4FoDaHY/eYbNfEtAp8IP0lKuEishEHvCo7R7396d+7iKrlW2uaNpSj6JmCohPo5sruE3ViCOZm1z
z1fqOh+zYpNKfJ41YRMOV0OHkCSAL8R/qg7ZpY/awkS1czmfp14ffgwU4cY64+EfQYioDqd3o9q9
W2RD/YfQJQRxp9WnD+yt++JxH4qkf3dNRs7ZKXTJLADlpt5fGXOZ1nxWFgtCNzwvfMcCVwyKbG/e
ySTq+EaqWtbc9DVsv1YwLPapTvIJ/l8pu/0uEs1fO7WNf0xLrfNvzsLcv+aE0FGdzlxe0hEL7GTV
lc515D/CjnGWcONU9ZUegvtndDYixuxsyviqHH6sJaoX4jd7YWlBirD1rsF5DY2kMuqxRtdskTFA
YFwn57sMgxFa8sXN7ediS5jDxq2Zv/rmjsrQnY1x3YiV6tyIzAD/vctMe4ZPHg53UtKX8YB3dzgu
v15Fcz08kYs4JpyYHAMx4oLJ+BUEAifHcMdQfkF5RlYXXC7xaYRxM9SJm8tAp0w/idsVfF0T6v6D
0VRG4yhzNMYtmOtgTrBEBcQsecl7aQf8ciMCgLORy69P7fEPXkpa3IMG2kjnIjA134lfV/Snyou+
Hjai/1A5WDsyt/KnTit3DOZ/jC+M6R+OH4UhXi6DrAR/YmJGc58UXWUolY94tJFSeTR56jEgYS+3
8szE6mTQL6PGyQHY9ngpTykBD0t4MF+d7hBnxMG+MTAzYIvJZfsTlcHvtnMR+A2MeC3PsddTHCvd
cb9Ho5Y6FK2m/JHYQgmLViH1ntoTDE0E9xPT6i8CzpbC5EKhGgcFye38l8gOsUtaYFI3H71mTjLU
NN9PBMhLMlxocsk8rFRi5ipetWi9K9shQZhyQAU2Sy75aKq0pqAjR2N/BW3ZItxzPDlbL+g94KXR
x/LYWIqfLiR20niG4DlXYDsQsULqz/+mDc4Zl/Qx8RN+HGOujpA58x2YaNceBC7dV6SW/aerEmJW
ElcOWZdF1yDgfM2OQFpLUBF7OBiWOSD1ilBCo8dsDisU5OLMD3cJJZDVsbrMNNm1N3zYJ3MN2u+p
za5q/lSgoLygrvWemv/Pvsdpt3wWJcY6KoC00AGPU9SpXI8Stg1X+9L886s1yA48MMcdS3LMhMwN
OWvky7AKp/KYlaVOvMTO3niaS6IJmv0gWK9rFXekTJta4vSuJlJN8VheLV6+H8SLBFnDAGbI0pEv
ThUM0fjVdj4qbLO8ECY0hobic4eNwK6/W/L2cu7G0gz4HyS2mizPWda+vq+Uum0cEdyOM3OfYs7K
27Oa4zZsoqvOwCv0soRNDfVeyiBUshkRpYhPiFuqMEKTWeWbLPn0DXpJ55DwgdPNaXYce6pew+K0
3Gtcx7RlDQfl03d+WdFRbpFZu4+rF7B5/NwrAH034bBta5/P+z7twML5Eo4Q60mvbbaafyvqYA/2
0cBWkTbItGpCYbCjPmqcvxmlVQkIcR6OYsr4/ljq7KrHRF6GFeqLMsVPAXPQ3TZ+KlHdFdC/l04i
6hY9mSTIpROkrDgETyV/A9nzX/lYDqvIhG4JM0Jaw50jWafp+rEhqMocWVJbPnh6pI/GD749pZpT
vzygdL4Ly2NouAh3Ar8iDv+MSvWvMVc9efShTfEBYzCGVy2uk4YU6DYzd3VIZLDUOJKmmfErAobw
UlngoObLRkuJYBqT1/MExPlpIxoj28j1Y1rXfJRYmtDPejU5SRrjCeeiHC/qxwHDewWcicLU8XZd
JZccH0r3cviQ1AcLG05OdQujjfLInJY2LdjVP2vx6BBP30V5a1ScprCzIlRVrSzjJVO7dP+LW7vf
BWC6zzxrsMgP8rp059k/+hBNnJKxNX+xPJH5lPlFfF4GXSrHeq+O60c5YJKtlBH/LokWF8gj0Mr+
Rfv2vXKREgRSqFugPkxBMKO/Oeoxp1IHYej7KB8i3iwM3k3of0MzAE5EiiSISezUHfwX2ahB3KqT
6ZCfPg2DthB/IP2XGZf4QVLKQ5YrIguV+mmPT52C4a5em4OToVOM9jmREU82R7vN+8WBqAoLABAn
hlxmkPrbpl/jxyTu55gOzcFiS6mw0UshD6bHFTNrPUpKryn15zC0EeYANi9hcU/cfoR7Mwhz3kfk
020NX9MMEQMkMsUc/JiMyDKYT+F+SAroPu9vRHE+v0TLdR4gqBOcwVuXllWxlplOWwqN4/qXb8zs
EeMwYQ9ow5ZHNrTGOonkXxfxmzWlsBNl7dsmIuypqYXw61w8qpO90d2om0jxX9DyPf32qrZ8zeCc
Az5Er4T6karJc5QUH5pRFkn84e0CkdtvkcnpF02nYdf010PRuRCtFQj6+gB1tOPLdogW3QoQUn76
fUJ79dTnEiXRa52BJzbcXGt0vrEPwV/lvqrWxclD+H4AyKxU1PJcBY8C+rfSeCF9+ILjQYR9FHW+
HMz4C6GaXFyQyHiQEjZwFNZARj6rTvIfmMWdzhmhopWl+AsSGBADJ7m29+GmuY7cXyj1OT0mjWKi
o+jionBGhmaeMHQmFgmBev591iiBEgQ4TIc+ntMJSvL26S2mVAl6vCLmpT9nAVe5p7drfkbQ6CqL
UoAXkW9gO0HiA41g078qzpPNc5vCNrsr6HR9GVC6fXT4bpo5AbTlpO3404zfsjPB+CbWsLc5oQYc
kGAFl6A5aZtwXLhfq+Y1Xzd0p4emoowspcI6o3r7kJXCRHcWfF2II5hMy2pqOhPzbufVWCNdi7i1
PL7x2plljvbkhlXXI1pC10HQj6SD4dUpaEJeNiKcFrpRmFVrIvDNoHTRYJLzDCFmg5+2xPdQTsIf
ZoRlPmPJqU0ftgmksxlnAXDboNTXjkPlYQZ2GgDs7Ju2nG9MfflVVhDfki+V1bC8gylnJy5NXb0+
BZ576dDdbI9LQz7mdr2Kr3WeJ5GnlWQGVJuyyOmUieczDxVyzZngW1LU/U21+SgdNhugTU6HEsVZ
DSmms8ienq5MqZYjj5hZnI9bgzwDR2SNMEFUZ6TkI1RJ+PnTOXr7vqx49Og4POFbNLn5c1bVJdAV
NWRIxInvA4qLNzs+u8lPiX+oHt6/1Ewoie+P10XdG29Jiq9okGjyBV8uvh58X3G/FM4RmBjyKzV6
1veabpkMQJuYnld9xG2gB+lETrgVDidlAmdWn2P8ydeT45MFUcBJ3uNynMqfX1YAratBZNjHrF0e
deUXEErHWWkkUjdVutOGJWx9a5WH4f2bhnhhwRSEeE9mOYUm1ETJ35srfE75yMItJVu3p5EGYxA2
rz+70X/qk9Qo/pyKWLyMx+qmLUf4JGWxjCL5IQ73ZiLG2mOeoiR4X7demHXw2xlb2vZa+zjreDbe
MTvDvQ+7Qzf6Al+p1CiZYiTR49vRiop0+USdQlY2rDMxc4r5lyKHAWHv4FQ2CTO1PHRzNRfEMfTW
fwEu6H+tPKCiFesGgl/hzlrXcJFBjbTkY3uhLKjIhVHQxdJyULLcJYJcrAe0e3fGD5GxVxasPgBk
DGVCllmAvtEumu6pFASZlzp+hhdvxjYkSmidyV3JTrzDwqschEDmKeAlasFPG2cFCmV8LTyzqPcE
eWMNAa3t//+PDl6t00LPBfajFUGXBYKuct8O4dmrC7l+PJxHH7tn5WS28Zsq66R4cRFwnir25X6t
2VD/Rk8ngVz0H2VLAxtm/6tK6BiuwQdf4sJMk+QuMIziPJdVijgs24wAdhzpEZHbPF799E8Uckn2
9/IjfPgLsK5vFhnjrQW0PKmUTbwRNX9m7o2vK3yrubGeWjUb9Rnfg9TmvzGDpf5J1fRSvg5NmsTZ
IBVUnNrxP2IbUqlRRvV/wDSnnyqlq+9zuUR6V2dvl5wWGFpQjNFpffkCAwM1/oE4VeA59sFEcCU3
O7iQW/CWadP9dZniK6EY9SE/rD+YW5fyCzl7+UZNS55iRE0acTGrwb2dEvi16Lv6Cs5xjandit4t
VsflhTJkQlQi6IxdPEY9xDZNiDqcdhzrxWyu94mFKq1MYleJtHVh97RbcItyWUedj6yKkSlFpU/4
ERSdSo/pqveIks/T6jLBZZiNjzHRTF1P2G49gN6AEtirVXMK6BWwHLeQDXMatkm0vzu36UNvBSOt
aEvP/LltUtu/grTMNm66J/FpK7j1xnEAVBEIW0bsXECrutleGMC2RVa4/1UVDIAY2sZu7H1jC57J
DVZKQuEoQ11utqREmyYnqG7M1ES8FW1Pcaee1EO+9Xgq2KAk9RohMbcexIzwt5CeCeJxkMgH+gLz
WJxbF0Zy1tDSO15cAJkkwHpziGAsv2+vK6D+W6rk93QDRH72gQjBhb884E7BugHGBfGeNC6+VOBE
2M27yrr/j95cYwu9ZYhHx6tyqUEGOf30DURNpMqHk/ocGzOH5hngpjMQCOmwem4yQttSp7KhpcJI
zc5La6KCIYq41UI36csOsnMW9AO9yvM660mwDzUwVOfqeZDf3B89isNlsctSiDZBzdNB79x82zFR
jC3Cvqt7IkmiKF/jjg/PPRD1FNUEC1GQCBnrzCmmc3Irdk7mzjX6xZG2YP8wmyIsMXQCymwd9S1A
Z9HFm7U7rk8EkzQ8u5Gjf7I6trAWubd6ERBnjcZYJkB1k/Kt+T6WGa4iAHFlvzZ/boKIAW01CmtC
lG4lX4ULxYDj45MhZCd5FPYhsLZXm8jgxGh6sW+4nO1gdMJcOVkJa0zw0vmr7ESlx8Lr8VXWke9u
JIRK+iLTLdKX/CWJF3AErRypuQxqH3wNyvLSnl62HTny8JlCKKw8u9BX25m2PDtN541bqq5S/Zwy
k3gKXSIFfreQBwnxmanskBeWoKL+o2oGX+tCyPQEy5p2hxTrj5PJVRzmqu9l4l+P1j2NLkCU+dJp
7bfO531F80a/6cj21IPX3rY9TXKIhtUNYg5/L8Rfkj4VH4+fa0s7Bip7d9mb9jBQFnpcAhg+S1z2
ZD9xP/0svNGsRoaZQndpehwWKBOnKucfVDFYpEqDqcg2XETczbP4YhSJ7jdq5YzFLHbjyo5tMmqw
bdfKIaOCM7Y+LHsIx80Qy6k37xEPnYhLLKUWI5SlzqdJ6CbsI/4aC55QxQh4Jmdb9MkKW5oZMRUS
qDKuW8f8lnVumXsGFIj99bm9kGA7sxaYtHJBJLBrWtQzIzs0oPyFEEBqwdA9r+Ib12dBlZJbogW1
W1pF1O1RQOVQnjKw+rvC3xzUbEcCXQkg1K72oPNq5OVk/DPuexx2awflDWMo5TC7cBQGxEYTQAgF
2sY6SVa0bcMPvk0zRJE5aoNigLDEyLe3DvNtXzBSOlnHK+8TEaRXy/MJVFdNbB/bcLDUsFb+5mFI
tqfkK84Jtfu776nGu7yQu0LUuKVC8Hs0xc/2NRieqvU2i5MSlht6RhykmrXRi0BJia/ugRzbQCE4
Seei5k3az/iHpBN8Cu4cvFMDI4KwZ8QDKrP14f4ADU7nogNNGYDC/+E915T0Tt64XefpWmP/UX3n
mfJHXTQnBOFmT//mJQf73Cj9BydT+CaE5tTlkrGLDY0Q0oRLQOAY4ZaPtMwAG78xd8R6ZHNIiZcO
h5uegEeUbRq/ZRL2+NV/mYGfzTRHaJBPomMpZgCGBMQFQ8ywz8WTloJF5Z76REO+IvQp3uL8x3E4
RyNLwaz6Hsz9gUhInWe3uT5sOFwh4qkfMPzDUlzXDwZ5CrIJ5OVZrRC/+LA6aDFrUsIBCG5Le0ZP
ydFGJigW9g33X74ByJWns0PRVWRgAfB+n3EQWtBcdm6K2HcxykCIBTHLmh5lJmig+v5IumachDyG
P3hyB7On4vSz8AkhREYCPJ8u34v2+NF/Y/+le+Ijck/NOJMeoCqFNjne5jNnSk1wa/Ce/MruOt2u
WmRE4vWk1d9GZ4JrYQcNrlABTmtKiKQFnNTlXtLJtbiQY8BGVmJmnAA1c5maZAy6ND2yj/+InzvT
br2LJgCK7NTGZA0sUK66+nCovmM4R6CTRXjHyK9s75iSTKq2F4Gl9Csx0R+9ElJgDdfG5rAcO+8g
b3qKQ3YyYdJzDWBUsjokzM/97XDTk4R1xUPYo2ge6qpT5/k7n6baOLUSxNr6bP7c/ibROgX8o4dQ
7lnHSVi38sBCeXuws+LOU82x7pHaYAfYEbR1Eh8QHW4FcSCLWtIjE+Zk3Mn8LHk8/aFBOF1H8+yl
HWrOl0Q9xS6UUtTW8PtMI8sEghYEaXktee07YCy5/wPfzadwm/K3qsGvWHnswPJ1BdOPluxodt1J
NVFL5aZmHEnsxujWmM7lefWLYamLWjkojdj5z8jeLwXi6HAgugvSsM6DAVC0RiOjiqRPIcnSVvdn
TQlHwRuSrJ1XAJCPwSxPfKn/EenSaLcl4spdvgtH01/MWXNCPheVKgX+1LF4aRjpE0HxsnGtSCMz
27HeFcwH9sPs5A9XRkGbxjz0/eTsjNHZzf6y5WQtGgH3X2gEqlmZTA4eGE0NuZWsQgvrb/n6wX+f
z/IuuKhPdye6med/ETM0107Vr4zI06cDjca3TtTv9ejs0XNoCQwSfKaZnfvlgDC0wehRV3nEKi9X
kls8A9RO8Th9ZIysi2suUAEJtyTd5oqajEVIBHotamSTtAMwaCYoOIxZ/+FKwm85UR5IoezfVnxl
A7sNbQfSh0N43PJY4H/+rlw9bVTvQC4ehueWPU6J5+4bXR0llbfLDYkrcj23Hb6MvI7Jw81uA/BO
3ff3nOYHNrudSTg31ATGqyw5rN9DkW4Jjk673k0uw+uvls38Ox2GbyZuGSSEtj00XYc80cyKWYTT
55DvoU218chMBPiTXAxb8XVso2fImpDe/ZZB8ZZ1PMLzgjL8N8hYzSaXYp8KqtwG+KFjcZR4IWbo
BOXzPDqLnp8fNNINAAcvQvYfcZsMklmVsNfs12LuseAOtMbABUfWrfHOOnbeRBzWDCtwek4Gfvrb
MwKUTUS53Lh+pfUJYrcuIrRA0qVPS877WksQ6Hd7z1L5n9+CMKb9ic7a/4cy4fKapmwnV8Z6gk6D
TO3T5SgPMBYAHyAO7QpJPZTdl9j64Hs2v8LfWpAMhjWf36AFado1TfCiiNcgyWK4vKHRe48HE7tC
OJ39a4IY4mjGV/i6ppfXS2ZKkk+uGxLdF8CrJeBG6z2nvgK0Vm9URAvjLu1lwBl/v6MhQlxmEVTg
hP+lHSwaX4zhzrd+AZ+01iHj1GC3JocdEaUZ3EddJrFOFF/muLHxP7eTXiLeELrJQzno5BtHZRWH
GHciLqEG4WaGwqeglbxGDOWmZEMhUaqQV5/X+KYzb0v8R7Uk4e5r9oDMhKs6U9caEo6vTFMLGTk0
eQijBbsZNfY0MKlPzCTI4DjKsM+D6kUCR1VlJjZ896osO9yFprcHCSHgCQskz+SlWGaEyViK8Xqw
FGr8U0THhpDR6MH/Og1WPGR24vMkjERKrNwazRHfxLbx4Qn7izxlH+SXv1KxehuDW0DmLonLMwY5
2ipk48FjPT1DX4yNItzoXUEZotY8M5HlSK09FQaEZGsUr3Z+ZbhUiwa/8zSJVCbBSPCaHCpSiAsa
yDY/FZOob6yggRfTSPh7rMSsGB08cuQuCYyAB2qKqNeK1qUWAyQF6FmmhoRDF3QQ893wgH1yZoiE
PhUOg6E5Tg8Kt9ZqXWRInKR7n7PQNw3RomR1/Bg9X5PTfyL2BQ6PEt8/o09+AH+WtL9+s07kHswT
0DH4Swd1UyTu4ZlXW18GHU3lnCb20s4XijH5QJ/QAUiCO+gFoZLyTKwTKzliLPLtQBHQ8ZfnyQix
OjXWiQzp82fMgAMNXonuGYGw7oMAXb8VKD49nVyu7gdhsLP54m7Qo4wof7bBLT4AnEaKxJrpuDPU
5IZSGugKmmZ0s2VWJMSdNXzCYWHcmEb4BFpnrsN6S8CgTPeZuDyCk3DycV5xWiOW11Yu/xm8A+FM
NuSSaj3tPi7+HC1ce9Z8cWzRxfTE199dGYAWMs3jRAsQt+YgQeOqQ7NQRONnexoWgMlI6VD8lj+Y
DpG24JUSw6yNvqvRQm2xxoYfNxH2D5lJQAYdlEbl3OE4D2w+m7QUlomNsHj0F2MftrzKBk2GtShP
tm0ZvASRH6AlqsmeP8Lw41/1+8WfGUoJ0XfXioFvwaphKYwSqgVQjavrjpqg7Cu23IPlfDwRt2AN
IH+9dVfNFnIhpeqNIRDRqL4ErEjPvmpgb2hMS+ALxa3INtCci63JfoDI33rzr9QJF60f2N4z+yLC
3H1eLPBOXWg9PQSGHF/LFd5WrlN4kC6VVU/THhvbzCaJjmbAGlM+xH0hp1R0qp6LF4V3NtzBYX2s
WdoXeQj6hKU2ArurGq6bVktTJ5hGfpQqUN8H4t8aJghdsEahVqGXcvq6bzKHf0GG+fiWHk7hoSae
OZhSxbQLz4G1lf78g4y2+GJRbPKXrzi6hQT20gitYWD855zSVHqItJQf8njqSB+xwzgP1L1DjBP8
+HOIxPkyp9m+ih84yamvf8z2spdesOfY5rXcWo4lvpQE2GI40SIRnitxokvaHiHg9vn6yqll42WJ
e1KycUe1Gp5TbMCKPyOkwAdecSY0P01bKYT6CXNPdRX09xiYKlAzNINZVSXnIEingcL67JMCfmEU
X2O/Jqh2OR5CqY4wGMH/ba7snNsb5dd7MfvPaweqpt7rGg6g4dx8miTeF5Lo6aK06mpYu9k/idNe
pLJ0RHkgM6UUSA8kLacvXzRZQytmYcxuYtqL9k5YKFqvUCfIe7QS0Z74ASPYi0se8kNnJKt2aOZu
EvILawK9EJktPMrkO2tfYI8QaoAjX58Bz81FQvDf1unI+xixUIPEmoMEbqltIWoc2fb5KCLSY1j5
gOs2fYZZwnb+OALKtWKfwEFw3i8LyU0rRm0nAoRa3gv8Afc1lO8IG9iZ9159frA9ZDwajqfiZgeq
YLg8orZLgyFpS0XMAducG72at178i+SEGfI0k7OflhZi0lHpjiTPsN1dXJP5RXTjUg3tjSB0pUa1
UoHIoF9qeM7q93akPMGcjQECzpkpbhZMFRCMxB8Rb23++r7OllCrNHlrqhP1xlKMHrZA+SeKHZKa
KhIsLt9XKRE+SuC+YpGaU3q95izpj/MsepSSzE97a3ccN1mp1KtvrjutFTrOITWhOg5jrwadD+n2
nkQFymDkncQzaPSmNTBZZwVoYEkUVwiG4Fu+Eo5bOn5HDfdEjoA6YlrGFznwtV7R0u/O3Fo9Iuoo
0C4uG4u1nBL3aBtVbwO4a8OwxsI1VqpZwk3mE90SdDjA0dwGlWsAuA/NHiJTQcOf0m+h1O+gK4/a
dSAtjqvP8SSRhuaJyknXCt8kyStg8YtmXxj5ylK5MfLuVHwqADKhgiMd7F8+GeW6ytl4tjN95Co5
eZOy345VpPJhZH86nGgQqwZIhJZ/cVOxBH50UXqZEnz6lJea/44rUL5tiUDDROoBEzw42adb6OEo
x14C/kftagqfdwUdk4DtdL+IytJ1dJ5/VxLRqT1LgxTo0I0kn8/Umqv6pPAgCBH/1yEF+jCAdQ4h
ZsZrBemAWY++M5osCrHkV4CJtwD+Vjipp5gEobJXzqiPri+Hp41rLHIEaqRzjULt6WA2XJbtIxEx
LSQ89dT4u80BCdJkGYr+rKxk6qA/0RV0lpUtNQJE8SEZqYzkyY78XfVFLwiNc4zKt+zd97kw5rVD
TDFvYVLr3oDcmu5qgd7FMXgh9B07wnBe5j6Z5vv1P2mGbzp7Fthi2sbNeTsrzqtSdLyUzTT5hQcH
fJnKnHSMtznUl8mDqkjGQY2MumDZrtqaOhFuEICGv0GgbdqIIExnHU8WUy7o+o05DQI1rVMknuc3
LHLHxmw4ooQbgECY2/+z0V3Q1mqq0IORqC4w4xILmeqeQa6O1I+dkks8sJI39u6IW6m+hM4LPjIf
OxIPNYtWYifQwRGzlE0RHtNs84pNyEjeVm+97SqNmxEUN7ht8pJAOAU8yDbwJFYF0tH/KHB1kG/X
aRfZzOtgnyF6zTDj9hBv1IEt7GOFSvGLmmVKcarxm7ZNTqffOQKh634My37g3gA4SGSjNkquz1hv
IjFwrUyAkeIW1tJ9nMuicWcYTOsF0/ELOmJ0VOGL3ybjLaCyZLkM71TcAwKaZObG7h+QOoFbTMCv
XXconKf9OSvrP6osn9penKRM3Nli4XSd7xye28MCFxR0roGy8RUCcqr/9woP6IiMzrmbzRapt7yy
lMxJcBg7ZAdKvurYsPJ2DcKoCF2QDjbWxTFwd3UISZVC4uvpPvBlPD5cZxRhzyl08ZcqDIQIAom/
WpL+tcuMQk2xFbDGF3oOEnINo2ClGQeOJgw/lAMBNEFI1uoAPjIfMOHfX7WG6nunoNGjUhGKVIG9
6CV16TzclCPMBYy3xFqIHITUpO8SiTcpImS6//WWZFDUyWOUnsxkIW3SySmWYc/GivCJbgLs4c5L
WkU6K4Xp3uL5UZhfLmyNt9xN7GzL+04jpHqjVrVXie0QvCs6UiEdt2TNU0zauDXypent7uZzRl8I
6NXtX7B3dX/YZqIGNfJmcTCMdTVkMcsNa+OZSKSv7z/JfEMjrGjOWVwlfwV1jZ0qoVrKogvD3eUo
8FsE6/FwIR3exxhv4fIxTnvoomOy5l0I/R0MwxqR/HWdIQP25Y5ZaJvGACtheI7hzjyo7Wucw5Em
jK19bp24EPwMS9/Oadid+NOrCWGEX9wPXLt9hFuwmNLhoqx7VqyouAzZTrCsoLPHiquNqAAsSvGh
Dln6H2IITJAZcQ/cFnGzSRKYmcEYTn20P7hfs8gM4yrM+Ve6kCutd9gTbxSO50jB+zdt9dozKhaa
Bax7EBiRyWm7LTeh7jP//9qSIPAU2PlCVVheuSgNV2u3wMJI89Wr6ciYZXf5oRzXCptMsHs82qfr
5oXfq19tfhJi1QlaI//5r5hYeiuS/5LJfbY2c7TTCKTzQqhIRLb0LtFeRs4ScOOl3SFkVySo8PYH
+Zxg1Dr/R0nBCcAUwuYLeCcc5GRoTVW5qNTuoKOugghgcmi53SRMbgkcLF1gsSk1FUJUbAgtlWuo
IdOmwBQOBrdUyznhKAK9Y44NvBpLvH5gnYkEkDeT6xmKlJEYdofc3+w096f6XiUg2SqS3WNVVMlB
cJ0lZCmYUrIRiCHsLAJ2+dA5+Bi3VLpK1fWUXvFR6rVtlps6LSfqZbjuSmuft5y+4GUVNzsti9lR
UXYze4fS9QkMG719j4PrKxQQ08r3lOkR70EobnpG+5BNBWBUMtEi6fqCDMd5GyVuNOl9LAOw0W85
wvJ2fTR2BlZOmPzgCDzdcV8JJp/H10ZckdY5GxTGjEwecwj3L//E+cOXCBs25evdf4bgqEnj7U60
n1gWwJ8vD41p0UAKxZoX+X0lBY5R1+CW94Rk5h0/z9A0HYRMeBDpNEyssBolbVRasilM50Hl2YCb
CpuqptLMOBK2vVAqXoxT+DlttkjuZFccw5Pl3ttl0Jx+hD+hr3DOXItB0sw93d5+Xq94U6Ljky/Y
tEYFbYyn6werHzBiJCriTy6cFNh14jF14ebm7UQw2FpcYOdtVwLCdP+cCGH22JmhKFp+qiuqxm01
QDGEGVywHTqtYDvXN1mVZW6F5GPj1QOCs7M+f2VWACnCyygeiwUNgaV0OVTdmcKWlvjiTA7G2qHY
5+UEdeaUD8s1CyOxuoiEgPtPZZfZQz9kWPx9+R9ZMYcD6H4q+jQ6l42kelMNHYbHpyqdFPpwR1R1
W1trsfZxhnE7lpumk7tZ8/Zl6RpbHsd80BinjbHIBoeWPT/DD6DhigvIjzzgMKU17nWrO5UYr+yi
21/udDIiCZLI5F2X1iXKkwnByCEd9h0el/xTDlSsDISiUV0uLaWQZ2H0QcDBzS/Xx+P4JzCk3ZcE
blDBbpWrJpStVkpxy7dyl7SJf8WxEtEDBlOxpwV16cpa0RK08jBbB/wotZa3omJYZWmYC0j2mJlI
orxNRGKhe/V81N17uQ3A4ncL8RXRNIdecktafhkOojJziBJv08BUVnrgZDz07DlfDRWeDKclQeMr
zAXcXv/xRo2mYV3rYIQ/B83r1kr8qdq+s8RGc7EfyUlCOD+cpmyZzmwjPtCgH/SPhLbExXU+i460
kAhP4ifaG713pRVR8H/6J68JMLyml19g7WNYNvthiuU97roWcXP4avAtE6c/CQEAMSH+wypeot54
UaiKjCc8CSW96nuZvNJpk31GiSwNj0F+muxAq/HWPtEejiLUhx4WaQTmHf3tc98eqcV0cn6/WE9q
7huTdOQ2Xoz+V/wwiQ25PI9AdNvzN7RwxrvrN37hkiuqEOKA2rf9wuGjC1uNoCMP68IuSIYnZQp2
GubpXWZK1b4g3rCp8JRZCaPPiRERBIv0CySj2kvagyakI88yWe6WTbpmO513dJwtWZ5AvRaeoJ6k
g0NRUx2msKVMnkx5eJmJzuM7gNphrQFsLRzU+g6buZhZYsOo7Fiw19hmIA9labnhbVDGYefRguZz
lSo7ROt0gZGs+JZF6VQGRTq1PvfVjyaUHp7bm8sFKCopBNynZNA/evGKrXkVKhmi163wXt6JTESL
nOiJsJh7hBckrbVGzdMXE2TN3jaVjVR9Yce/YDyMWt47aLsLe543tRkTI+QtMIxKnatuWhMatM2k
0496orNVnRRus8SqjNil3RXhhW1tidluBsXsuMmTi4ZMdONfUezBSXZsKOwz8xO0Zevgac/gYAHt
PaV3Yx2Y8D6qf43ZoNozAiJ1V2g340WlH7L09t+vf/MgkF3f6VYUndxO5UUHAJQd56WXqpFIcIUw
mLSpM3BxBdrQu0RU5UMEKqBW50m5Ec0JjCKlnqV8OtkiK4DqaRy+rUTDrvwH29i+ifCr0BaaNYkr
MY6UNbTHg/hP6LAapZoxZrwd1QSDdxklg/IBLjR0xpHFSa91hILmyLaLG1SQdnFRElfOB7yljRRN
0gEGFDdt8dGuQmQhLULCQ7pDD+UQMxyWVOnweOvg0gTagX4wiChXzGtTfhQC6Cl2HrNiwYvrB0d5
4cyotI/63TIi+BmnH8pPzECkkjDlQyLEwksfUco6Fwe5EeZzTTmvb4pD2bld+02iZV+9CxjfIyn3
CyiQmwT2T1kmO58W3y+72maAQzP2DJ17OexWp6gYYTk910hduSTft330CdqcdRJ9BHH/BBLc5s4n
f21TyS4ZXjTw2TmJrp+Laq7ZSWLEErhxcZXGHsTPiRvmq7RKKA5vqkUf1/rJkSXbHaBq9GKEdiBo
MniGG2D8cSky9vuHaWRejAfR0GAIzjKAz4RFnQFx9C//9j+bRu4rGH/8hznfzY/peRPfSTNjJwvz
tnYsd4KqkJnueiBlc9lbsBYnCSuqJwLQDnFh5f3VTZn6IuB3U6AZP+0BC/pZzzQ1rbrEvDBD4tpZ
6o+pcInR2/zkej6K2idKnODsJ1h4JM9ssAV79dFYdHrjNF6wK+Rt2/FgMcJn6sfSFEcrSTdFt/0d
94zYG6Qk2JqbbR+gWsUawkCi+CwWprb6lhFfzJ29JKRvLU2ZyWlrpCgua8yw2w71/WT8CTB+pu52
+DfnJGYQLs/ghtxnbveWM2PJpU2Wpjr5NUD9Fl95UWbJvJF9OUJboi6SsS9pl3h1QeR2rmR8qIEj
TgK7Y6qEYOyhXOx2Hwh1HXLnvaRiKRJXTeubhISXF68xi/vbhDLyqg1cV0Xc35jiKQPw9F24OSHM
YuVWNubLmvyyx/rb+l8aJr5t3i8FhnRwCyhdPFxXU9/I6K8pSMmzxz/48x1Ats2ffR25eWpUaQ+v
xDz38ym0jZmFlCcygZJOk6wkHtHDQRMDkBDBjGz2QIR6Bkhp0OOkr2hL2RHCgt/YUPZeOG+04EVh
ygHEKkDDPdEZCQQAkUdphxdKxNE3sKWsDU4GiCKJI0qUj7/eIZX0oLEjnMyrCLoIbTIirynbrYor
OWPkEoQyoQtvvZ7aK+nvfQYqr+7rDezYYUyI4/EYC0gEjA5aqk9WcAS+1n/p3EwaPZCteaRsQzm9
8LxD3nAwyAm94ffSon7F0js7Q4v8JkGq9BBBVYzyrcMV/LUABlm61aryV7W9dmfcHd1bP95SfnXV
WfcdpPeRvok7vMDNi9Sm/eI3riRODTf8FtamuAbG/dktNqik+B7qUcsx6p8DdKbtTVhndAxYW8Pl
FepsHjBMv1FUEx0tVW0kRiFAI+JGC/ovwytuNJLrWy3juXFcZcfrqDwVq+B1kEXmYtIoaZEk4H1o
f6g2O5x0naC2yjwA0VP39MKN2kwiSW3C6j7HORfP/JYQAzIwqgsA3+biUOYr3LquovnBYV5txFWX
ODEPn7Di7c3kImi+kaIe+Wivla+m5ss6ONT+mlsggniG9c1By06O/tPrrdLeJoszrCpEQT1wzD4n
wkTdjT7I50fIaow54vNSJF1SO5S2rQL8wVUbolLLjt6yyLrdVqyGagC85F2z4k2ur99xg2kWYpS4
D8Gzww3KLsjmb9/sRaog+szyln3h/3HLuRMJ1Pop5zN/emQvoaFOtteItUYsqUXqlw0RHXEOg6aY
GcH+z95+MY1AJZ6qRUj2n3X9hKoFh7u5plfuOktljoKyJnX1XUzn7DWHyVaJ7+j5yB9N7wf2nOmi
4oiNq2H6Q/fDZdkeWYVJ3LNPcVUeJtSAV3zmlUhuzT5dOcroav/j5TKeohM7CVGwwdksmT61IbUF
sbeiTrOd8OahBjP7kqfg6YzLyT9OvQhCBf8J81YbsPQjRY8o9QvgHeCeSmpBqIpbFY0ol29zIWAP
FjjB1cBObe9P21aSt678MStGYaYW+xS8/qKAlRk9xVGxj7E+VBs1IHgo4r+sHXmDkLPtNgcGe+YD
2d/0rbQCEgLi234zjsvm7Uf1uZ7cibXvFaBZhRd8i9JONQna95gIP8BPcJi1+KAdDrvKJQQ1G4sY
QwcVPxK9AS8f2qtWvehblxGyqJ60Ps/Q5gwc5Edz/w8Py4lUcwIpGoloZvMxHmi7odYmsVi46So9
iTQfXXo25BpIKQF1mJchdxVCfpPtEDHtrC9J9ixfLi0RO48p96dZ4U+U0Md2uJG2mS1r0CSXpr8H
XwdpDBFxhSgusiuMPeV0NgtzeGKXon9yBJkUhU154Vhq20O8vG4dPreIfycpEjdR1k0/kgjTu+9Y
cMOEWlG4y9cmKExaDb6V4YQkz4KJohOanJ2hzpgNkZKBICu8Ertm748kV2IIYUf6zgdopgjzE1fP
WRCPNNdwL1K/VoJd2rXpIk1KxPWTrJ8W6W5ycBUdVwF0iB7wHfdpx3D/rotJiK4zSZXYD6xz5mja
mvBcOaQ63Nix6V3i7wNZFKati6cEeIVsP5/RhxXSIBNruMTWZ5vbqjhtAbIdaCzb2UnRJlxGCDEn
E7KJfIz3v7zjRirWiK/EkodwyS6IOGdOBhJ5aO5gGQT0EjGOFJ51QNArySI9wcZhZ+080FP3lULf
iCkVQmcEjDvdded++d161UkCicvKTIn5MeV77Am1dvFL01i6WTOj1xCsJAOSGFcNVhxHxVik0+Lc
Tw65h4pC/Sa/1TkSKbs6yZd5LEJrqgdljo+DpEKEic2gn3mQ+pIml6OuUu9Laxofejq5Urz2wvuG
cmNFPkix6+nHyiprtiWaqeu9oIxxz0TL2aG01Fxr32vAIcicvgT9sN1KjJMlCWT9vxrG9n1oeNMD
lDfA53kythPfoguJPy/ngQb65wENb+jn1Kz7Yc4CV4mR4vP6mg8a7ZAMbVJRPnFPTNT7MD2HJ460
DqAfvbnL8yj/0xgC6ZoFWaWjA5uveFYHyzgpOBXrd4hkrp8qYCioCqIJtd9Mz+r0zIrQf3DvZSmN
TcxOk/WdDq+fWHtunmFgrBuIuZYWcUZ5L3w9wicw1ndXLhyD52IMcRJ1fNMRMvSAYdPv65kISRa3
VVYhx4CXQhhfYZE1f7UX/5jbNMzBEJxZV2DEDG5zeECnzZ8aUnWazM1v2JIpKSYXgpUQhI8z22e2
QLudGLhqPm0vcaKM0Xk5p2leJ+k0v0T7PRWThYKic+6SEa+9dmdZu+Eu88cO6hWPjeRgfSjzdv7d
1c7UsgWZiyJlwcQiCj8RFggqdSoLZQGUtZegFhWU2V7Ac2mz5JzXGO9oGcyon8upOHtkjkiT5c8N
aK6lHxoVb3t5fkDBlu1EayQqK4ktE5574H2o2d7reQBdY9NS4zIyFJtxRWU2P2lRd+hl5ynzsynW
8LEFyhi6jyJ3Xs2VGYJchRpvOBjx+BvNstn2mQl9S/57hkgmR9IQ64RXrKI0YyfDi5AQVL8k9hTI
uYFni0KANcpIHmNdUKJJE9bOP6BHPbFrv4brorMX5Kt/h+8cihyZ23d0KchEsl2TfOocv8pNhdv+
AKkVcikZxDCUX0ikcDSumvjyngJT4M0XNhxPj57NGsJjyyLJ+p9pqNFuRQwVVjv5/pT4Hmt9PtDy
jaYlTBh/Vz88dbfbAuO67A6XWycVxpAI8uQkJCrQiaKtzenXQlC6pmWSURfAc0VSyladSj/SPmnb
H2RGBJltbvkrFxp9W5/ZuJEuOOz4PioBflcJ8oNezYY+54JSlj1iL1ShbTXnT+6Xuftoys/YaK2h
Dl+ZX9q9kyDc+D7gW/7YerwxlhpDg7zSd0qU4fVPRyj4ZWTXut/XG5MoWng96tkwbKAlCqCFREO0
Ea+eqy3DE1WNuTqDexR/ZaX19wsexI4dC7LFNew4PCW8oHPUxqKroPWrSaXuI0LZQzMRRLW7UzsH
/kP2V4YBGYqy9QBGaJeqjGCwWIeUQUiWAMZ1ek54+id6QEINR0jjWHAnmi/beJ9+kPhJ4JQoV8Ya
pIfogKaG+EUCaOtedvFuYtid4pDBbA1vdwwzpKkk/B54Ow7kfnlGMCUxG/oKsZUtArr/mSKL8CzH
W4dnzuVwnAytY5fL1sUDFxaWYddnEh4n4rmW3aMooOdIsUWfOylK500Pk/8hC3mArFPOGW1AH1Fk
1IPmlJDrz7yVU3byUV/8y8lTu89rPmuK2rmsGfYX+crPamyE+Hs3apT7sh2y2dFxBcO5SdU0hS07
CvaiyEdWxC01cMHf8JZnth2lPcsjuVAlGNo4IQlmaSrQ8ptzKC71AbJNw+tyeUoRazNZt0O9xmsD
Rl2VNUU3Nf1UwdG+itRtETiEveSjgtQX2VN2jUFaeNrRsfrpa7+XRv1YAw/UrSoNtdsBOPeSfTa4
rSaD/5wApA3MckESwVD/KerohBjRuQUQ7DUoobPAO7+3e+EZBOeYDztB/UyU6TwDesiVjdy6+Ytj
gBpz+vbz1j3j7tE27aU88KOnruaCUHzXqzuI2xgtDMSOWDLzRDd3CS8LixJ27Y8nC0v89ma57eBo
B2nHMBXHmOyuRXvZSycvcTCk6HdSWrGv7FVxr9tXxmw3Et7tsuFOII5M52yhoSWuSFrgKYd5sQ+A
KMhc/6mp86YglwhU/bEQfT/2nEl8NF+i4K7nsbKDNd6piGYIILsg2kMjY3CuFLiJWGU3rbtEcDKJ
KQerCRBHmdCHB/7oCkujxxGWvLrRUQS3/gMsBiiJ0VPn9bkBWQX4urXjLQI2RnAIynIu2E0+JVTp
9kQ1sIEYR5DffJux/vOMisBgDiYntwzqKGPuuuef/QvyC9AnHMvDRPq5vB6e2TNDmcZNsVrUIFLi
ko72cHh6eReao+Nz5XEOBMywP1gLEQusUw0pBF3C5IX4GgjFMe7uAbdNJHUcY/CG2tgRT0+Mk5A6
17uuOQGnKAOf2F5bcFIYhwQuEeC1+jCtygyl/G9O3EKdj63zixgPsXAo3Mz+7nn0uBMJIq0+WfAl
dEXllffE4UzYFrUkfpyqlsocqK/S5lB9P1ySKPwi+3Fni+8SLwSrY3PYHZK0RClF9w7JWPsHVlS3
dD78U7bOvkC0g3ldwm9CUm1fMOBk0MZf2wMRVwl7upSP6mjkWJcx30CXBb6Gawt/Y2dtf0ZExY4O
EoZ8risimXjWkXFJrESeVtNTL7KX30vduQtR0XT/+WB0PYRpkx7K3thMJALHq/1VP2cNQTlmTYuy
b0Jv/b3Yxj3iBvcMVCATwzkQF2zJTP2az+1rh+kkZjYtJt5WTNzUn5ErybPKJOS9u5J1yYaQ4ei3
32k0ONdYmvT/F1os6tBGEosvvugK4bvLQQXLLNpsyicMnWgf4KQM/bTi2EUHZYg374IUWjgUyACr
IHbCasqwpY1DPZCrks9X1qCEZhYLkNsc0VDzlMKa+qcslKGAbILtb6RE+D4VdFdB42Sv7IKIKrLe
FDhLfNzt2FXfr7TTSDVmhjb5qq6x9SjNZ4vRopEAugWaz/9qjdG/yw3vFq9kHiOmfNQ+UufR4oo7
fw9JeTtEIcKM7IKz+R7fNYAUCm+QO/Qj3DhYgC8Sp7koR8jxTZqZVPYG/je+RxB/xIIw3xbUt7LY
2knDopwJqtppFLNuEZcRXhucik9dJbKHK5nXxlL9BL/PzqhrGnVC7Te5e+0YCJkyE0G9RY5YQwZS
M9xhLTDA/BaR79zL03Fg3J226M20sApTHBSghlnkhwS2ZApQeBYu5aLf/Vn2PWraFYvtXlmAevE7
1nxanyqB6S0DljNyKoPnAsy5o996TlayqUQGqhkOPwFdz7zypQVyTMr5FsvhWSdd+OWYlxt2jyXi
8cOyUtbMwlU+fzr2GGyxDzm1rld5qK9D9VFESIVXVxPnWfUjeqqxcZExOLv5i4sHiEh7BB4PiSWJ
0W/exxoML+R6FLxIm9Rl6DSPiERj0AI+UCQH4YO+rm5iFFSt8yYpgc91rPIXtSKJtcnh2IdpJWAK
FbRByMC5GtH8BlK7QzHlgTk/R/KoiqDjgHjoNH1tbDs2fhC9Yc3ZtsrBvc1ra3hgpkMLHrzWuELo
PXRRgKQ8jjh/OKyGz/vM/lPTQPQ6XiSwfQkJONDRQBvtesLlknrD4n2xD7dERday
`pragma protect end_protected
