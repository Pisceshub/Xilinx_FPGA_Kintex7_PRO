`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
BCC9rc/UvLO+60OKG37h+5K6XVw9+xBlmGSPNNtCyHiGBNAs7uE+P7kAaWn27GhAeEpR/kFMWCax
az/GVqBT8w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KqqDQUWeBjbeC5Do4n6RoTO+nx+zDp05oc3Bq7j9aHdTCyJc3x0fyRiN85/GGjrUv39QuhEX8Yfc
PQieFCLLhIDiLcaO3g03QeMtoC4gucQf/+wx8FMN+etUNIAKvGSpHcDF3sE+QU2wR0z9UkcquWwd
T7s+2xbq6nw9IgjIn20=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ArQFRYMFjfIqnM01+3BErkf89TR7vHqh8+aVuOpf4ehtdLgHJ/5eVLEiyKB8J8p19WP3coK1LCXX
zKhiKuxxeGtbGwfm+yWYlBx9ENRZgRCMJMCvUsDVN2so7XdAPwkjqSnh0W76/Lhaf+d+pvRWlgkW
9DQk2DdXzM4eoYWj8692SXfxs2GVr/LFsjE70VNgWii3g4b6hbt8arRzcBGb7WdSP01/Vrfupwes
wvc5UsRUnFw41z3BPXfnJG4S7TLMUaKkpXt4XkwlgjRwtf/TFvPay2nUHGQKbMhpn3k11OWjCVq/
je5H9c1eGYvQsLZXkrE0A7BXPj2zxOkaxG0eew==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D+ZRBE6u1yF80QejORI2YlK5RectTc5Hc3ZGgcNzOnHuwsKdRLXxgO2EwzuQORFrUAcI2O1GShfJ
cDaxaqcC2RUD7RA3O2LsbI/gqaNLWKfE2cPM5kyY4LL3UpWPM0Uo5ak/GypCYQ+UOf0Kv83mOrCw
gTGIytvAqr7oSLY9s9w5ayy04DJKSe0dAiinfq3BJ0yg/LnSWrLQBOBrA4Wdb3lM1weRawy6ucLs
RISAq5pL8KX5nYwI6yisEb3R/a68Gt9JyNzCGetfTfKa/ZmZFgr4Mj4aSY4hNGRM3OGia7fX8MI2
J9WLaNV+MP1mjqAewxP7QuQOtPQpJ7jXaieBRg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ntat/Y12i+xTz2OshnCjcnc8y9zrqQygo70X+7SJQZtc4rY0Zflni9gN8Z4mJ875xuUjX+lsIH9Q
3xBNfK+u4PKka3FGIKhp3P9okYAJ4aQHDoQHPys7ay3p9o+QjpDu+LoKsYOvKcQvSTT5h4JB/ADm
8cRL+CJAT0lnMoC1oD+FzJaGD6rbUe/m+ozDAZO3EXBxQhmIERbrgUps+YqPcCfIPBOirPKyo36x
gPacfOHCAyEnDGqsYlZ8/OKD+fUUWGYGW1h+tcsLksdUksFOzpwjaG/aylVqeGnpGGdju9YCZsxR
FTDPxHHSYbWz1IdEVen5mJ4AEFHyNM1FWcDu+w==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iooVi2sFmNJOwue8KHSUPRW3tf4tB3uu74gs8Z6LDvu2knYgcu9jq++JPYpGEqao7R4n5XlVPf2c
k4alUHvp6Q50up5xf2+TM6YAlKOh56q9Kx06TJnkavZHpzcVUxjTO8lhG7ZWXd4Gx6jTrcXay9Lh
hZnVvqIrYIf7F2M9BVU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TKJ0HbePLQGnDE6xQ2nS66ju3E7NpHUMIS0eN5TmIrTiavo1ur6LEw91l2unykROGHhJ6ADO8P3+
+vp5WK18tY3bqWh/q6bhiVRnEA2oMtztFhG2JpSy3iPMMzKWi7QDcZAMQdJjnf/G2+bGK0FCj+pn
IcyQWYXOLQCp2MP5UnYVxp/1/Rseo1YZ2mplACxSxS0C9v44JZ0uWfMD6EGmpBALrJusrcpykUXD
E/ZZoTwRUL3BWG4AsvhqsJUYITtSPAjRUg6DenJjWOgD37PK6P1nngWyf9Jjbs53XYO39akVpu/l
Uewa4cLxL6R5/kYVDFXX0OuYcl7BxOYxaBLIeQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13648)
`pragma protect data_block
eAOL/opCDzBH1z0QvPCIvLtbT9rXP0S3MoOX8sbx7cgUmGzbbfnSHnsDbxvpXxYH8/vVyAQtbxq4
rKpK451vCkMK/GHqUODpeoHaE91ICrqdIZchDtP6KxdABLX+zlVsmy0BLH1aj0L+3iON4jr1iN0o
Ub+oT+LN0U0ccaqjfdM+LxJB0vkvu8WtFKU9MXNhf1fktz2hn/SUIqEfZ9M5GVeU86Ckp+KHBE7h
PwH9s9LU/MVT1Bhu+BbPPlT0Ovzl/o/ocyUXWwLkaW4vFjM4TBfAWF/NF/HCPfqBo1IIVlxVQyGO
fc1BdKpbIPpxWEZfoeJ3fi6KX1z/fCtr2qoizWQRZlAuSzDFj8fT3AyL9znTK/qWiHzdXAfPiXRG
bpNPtJOnyHPXwdov0M87sZ7hntGl9zV8byvJU0YiNUsxg+Ei67Y3hfzCfdXoXoMMz96qtDZn6MaJ
sce8Lev5vL5yIcNIVgPPC9H8CkKhQH+QQT+UhqClzuQQtPekT7oROQhN47F4g+qLGxieSKm1IZzM
PqRpL2mcjTqTGnJTnC9GE67N3RpFlbwubQ9HjRJmfeGvYdgw2N/6lJLYulWQXYa9Qg7HOlhbXLfY
azBJxFyA32tgcboq0GPaDXDBhLrfr7YXLEn212wp8pV10OadwnZ4ZkQTGZIM6dbeGfgjym/FbHjA
5E4iPtsZ6WkK6WAV4t6txP/q7EzO6zVFg2izkPS1eAog0KDSbXR/3MUpcoA29Vq1vNTK8Dq+Jbib
dIfjTj6tzFeJDhkwY+peTw2C+xu27JmK9uBik098bNOBec4KbNmvQi0eimNkHy1E82znvbjQY31D
e+Jy7q6zdJI4tQDQOj0Nw0rpIu/g+BzuyiU2v9TVLA75LZEF41bBhP0ec2lWYLEYnARpYuF5aAvH
8A6t8VnkXJsFAfc2nDSvFx4Ofd6gaA1rB3P6wP8/nspAO8XWpgw49XKzIwXs635kTAZHw0dvquQv
KhsK2VtD/2HB2uedMkwV9Dqn26JUgWJdXbhP23l82bu2J0z55ndNDhKY/jalNBH8PuEMEOC9xpdv
SmQEV5d49mYTN0PRBV/5dkH0fy80MusSGHUTFbWyCQX9ciLrX9J8K4x9HwN5XqLbVZw1yjRudcex
PupEEx2w+iDEu8SWYDO1ENJ6eHpJuvDsSu/RhHSPdhfnHI/Ex/jyzfzLpXXNPKUprc4fVOdd/HYA
8BDwp441Yxif2MYgU1pTqnHdHOeTS23c8/DaEAaAV6n0EtSAolpOeSzuYmThjx75M81YI7ZFhlZH
xStLdSPRqWoabAWVFUhNRZAqowm6LkyPZ//WVcpvttBkGcpEjpvhk//IWhxxNMiCOOhMsgCFQSPB
5LAIV2RODP4oPxTaVcgKnj3v48G8uwjL1D1nd0odR7J/ZgWTgJ3CrglsGFoU0884HmGjHb8XsXUX
G+ylQTpf1dEHkaOyOjTdOUceS5VGGCh9FlkYIYFij0fxc8/9JF+G/8H3EkUPdeiJkVudReJH4eyi
EKQ9LZJSZ0S5NlqjmH44Lmh+CYtane9sfTOn3YOi2kXTz/VkG70dpMsQkOYPyu5e+UDnFs1lNXfn
TYAWqD0n5u3fwmbm4DEDiHMBDzdL8RYrfAz9fxXzV47Tf5iYkekowTTv8XbBRjwk+BGm5NTZbWmP
e1FO/61e9JWYMZFy3AjrJ43FM0Q6DIktO2xKSjEJEsNBw00uxjiIi8S5yUPgyEvR/hSUKhLC4Iuq
eZxdtL3CCdCs6ZW4+z5Xd1ruVVE0qX63SSfhhFhWTYS5M2ja+G65OA5NtXGinkwQHBTxQzcfNPQL
8b83bF6KctS8MkDz/dJbWpIMRy5aM4mcFnfkGxtgPR1Q9FYj8e0badDyi+XxC1j+8W60Z4GMvF+b
69hv+kXLw9FI4LzrIBJD7lZPiDtdVQcaQDdo2ZuodYAgPs9CATrD+YCi1XzCTpYMJx7bLeCDq+rq
xOpT39T+IhW+ByDi/khOgFI+MD4xxDZIHQF58vDHkN/vdiAlxpWOe6m1LPd8LeQrqjP2qTQzbOAu
iHcLMe2mJjiavrGrThKHJfjL41Qn3oXMS3mJDuOP5flUg3dYG7aZTVuJ1y4Hrp4h0BdFiguQUOHw
MpXcQ5B2xRiyiJwQoXSfhdY8gcYkG6l5qUApu1Rr+aeYk2WkEsqYIkvo2Ded3DneEVsLFDyuzatG
EE/8bgK1s/Zn5tX9TuFr5Mtqx/ZEDufqjvFCCuV9sAzf4RAuQUKhjc5jHWJRgjpjJXqBuR/xdPFz
trA9M+I5BNOnmwmSVbw5rmjg6gufsO1EYBQEwzCrpPPJOb2a0IhS3zAMWsdantZO7sKXUqn7usaa
a43IZTQVaNu3Lu9bMPtlLFI1iUFPyCTA6O8Sh5L0DNNF2zsxMdCQzYI6I+xwAgnqEEWdBG73Erdo
zdYrr3H0ZjVmEGvGXNoADAvqiKq0gBXIEQaHkoTQRXEvt3SwFJR3B9aXz5lrjFulrMjggyJtFSb1
tRTcEMTzSL9I0CO8vXewbdTpLTQ/R/0rWSTyEc/qzoL913Ujya06ieuyfez+Idel/Pgj82rfuEeY
6bwTShBEof6t2sVqqeN8fglhAf4k7gxDoskXeEilZGfyc/AiIuZzqn5NgKn6twwGIzkI7NMfUCXT
gG463ZGTIChE1WREMj1bcRMVWmfAtFtfYCkCsqgIV+2IWGmVT8UJjOZ9QZ/PEvbJyWMRBQRwpx9h
Brfe07l8aPpXaHfaJekcXPdIhzsm7Mep+0X67ErLUOS66LFNDJM4w5IJ2FpaZOs47MP7mNqsKiey
FS3qSbPI6eyBp+45gwkJlhTMwtXiPIuJPzpCJyR0vxaGX3OK453HFrzb52GmggC6UiM+uc4NkSdE
ODu/SkBUvhRlsKKV4S8g0iU4AqeD1GTpT2+y/P2QnrVGFdatQvtT8JFjJP6ZAWUGhGmRdQUia7s3
aueAO0HEQsAaW78k8zwxdE0pyzhhqz20DE7igVbivNM5yR5ZkPgUIhRLGHVH6hoe2YFBpK5zsGEm
EfcspUYuODNWbo1JlK+RopfTggUbjZu7Lc62JR3+mYjoubYXscp6UvJeHpUZYAlQQIGkiKMWD5/r
+BjU/PQKOrD1hMdXVLqlIbPydM4tbVFbxVB8V0oDUPU1NypAIBl+PRfUgKeB2ntv7CyLAXGbb9xC
GbcN60nBf6Yac57RfL4F01A+2AFTGcOkZIpGGaW/V5PF/L+xr12tVkjnKKAknTy2+vQbP9L9dxMo
eCQtsZUx/79UyzBYLIUfhwGugxsfsyi46PBERvE3ynJe4C6McwQTUcnA+UitIobdERhUU4TUkVtR
iLIr/8qlYOfUR2gmhtGsvf9bWJ1B0Qt5wyu0Oi8nYJMPh509kUVt+IX6OqCOU/Y6ETEKqzGfGsT5
sL9thk/vxACYuwHIqVZMesdaCZl+4m082i9ybWDLMjaOFCnOFmEEvb/jnTnvEyVv5XKFj+2UI8V+
Fl2TiykUPCXqzLU8FuFVSkOI/zXiWY8/b66tI+J1ik7WeoKxqceIiSGZglKgy2U0kJQhSoFGyNtq
KGfZAsEm/oO9sVDlMWqvVdeSDoAVMCgP8QfzcKG4adVyqYrcy5lnkgp9VzARfJ7pGhnC3DMMr52G
QTgE+m2zM6Tn/I4hd9WjSo6e24Hlz3iMBSlfYbsYvIxChkOubWKvT0rXopjuHX2uGjxCsuMI9apt
J9cQ/vHsNvCWaTqEEhp37azKt8n7EWbckGDD/dHGPLiTD6FcGYb+ZisuOruFbsWY5bwZ6+Sao6uo
77MlCCU/6ereeQNBte1JE++GVMI3tIdCwICUkDHxqUdksr3H9NhseEPbJmir+G5dXiQAdvajBPcJ
WrhbTFwy+i8RN5DGu94a9skQ8KJU3O0UaJuVVzLV5A0/hw8kxRAOZDBF7pwBo4jpfF7taazdGrbK
wun7hQsNer6muUZZJDWTNMHPp7AFhEg6j2zWo9cWutSIsimgflwO1ovViJupK9nFwhUoEhyCz7fx
yfCZ0ASlF/UW5sBE/Y06i/HIwP0kLYR4IpdCSbfHT6BzjFpENhbk3atawVq1hq4XD+X153WfZL0l
sey1ZTdXYCZOUQT+f3KMcyEBUjEcN8Myc+Zb5dhgPVD4KherX3B0UYnBpmyW1hKMc5r8hYrMEpyL
DO0JZDGphd151Rp09B0sviBb5+RoZu7tnBmv4lqO5BHaJ/p80U3zHwlegnO6nmc+oLa+Sbt4q0+G
OgyDI+i2XPnLO+Cig9VGKrKsNmYZL4F5mh0Va5MwuTzEGLcvQ5LwTUZ8G5R6JHXPUj3YGXa6/3jo
1iVMrHerWR7w7VhK9kMWWbcMxEm6+D6ByJSllWkv+3LWDwHawZiGuQFqgb2ZKsQRAqcnwXjtgSWZ
0Ul7C/Z4/+27a1ZQMNPMHvBJGtckloMoPW7zSxPPROY+qGFH4AKWeOKraNdnwfemc9igVovoylaQ
jKZo/inVaJ86P7gl45tRdzpb9IAyJaKUESnFuRZIra5/VgQ/43ZL2cecqlIsrueax/+ePdt27p4/
l5oGxtKCtmj9CYAbdyXL3BvrsxxQPTpUpejgVwTRB/hv4SeFM0/92hKnoLpLZ77wKzDMHrtOatX9
OyPPt7jsukA8QT8xiQnd6p6eEd9zQwnDmft6bYY8WSCdC1rAJdlli5qvHnDjO4MihrxUvRXXCSie
Fv6/Uvx3oXHh680O5lC6Lk2898EO/X/0jTqfhKnLCEyZajsxXWAQofxr0MYyUufEWCYwe3XQnlG0
tfZPf7WjxyzmYW09wdFSPX79uP62DcpFHI1wvT7z6g8O61rWDMtbR34WiiqK4A3h6P27UCDcfwTo
Y2drMUdWt1n3cUxIn6PxcFLFvOui58b3k+6AS8MyqIZNASAoQSdb6WwlRYRpzmC5ElQ07ZA6tIOB
Gt2F7tIHT6Vq/2nXNNRHXPD0WewmIq9/kmT+kZDgJBESqpngLntmHNmm9b/820qAAJU5SA0SWG/a
NzSzJgxM9ERuxIcmv/NpJopj4r2Z0FKp+K1TDN+EpUM95VpE0Tm2NWtfRtKxKC3iuCQq3fHc2Uh8
zA+jYUcKzFIoWl6Fm1jVKAzm3Vd+D7SaFRMp2WXZ8LvfAlnheNfY1yyiBcS1BPb9zZM4DIVV9N8x
ZtMNIDQ6X+vrqyoRXVdfKWQrEn0CfxTxOKAQO53TTmOkMHi4kvyMWLOpRYASjR/pp0TAv92IfmXK
qUAm7isPFvw8o4MgkP53b8uZahf/F/S/BlAzsmo9d0NPYp0ec150AowEEXhipId+NoQ0yFuaeVok
DdasIhrbWZOjNraFaYNANOAA9p1/fJGOxl5+5WeEesUpIIcUaTaQ9XVughBJ7wsxogpLtvNrLDVS
Uf2q36M/kI1FErPoTj78FTEsXQY+X4qxJEOXXR+5AN8MW8QRtX3Ri0vgtMjEo6cU75rDOx6L6GMu
bUbJq3Bu6TnC/90N53q2VtRCWIq9HUF44gKgY1t27MhVQiIi67eBlxAepoNjOgch0aBmuk7P3/+I
ZV7Ih6lqo9UXsjbm49jDMvTV6Afffx1EemvTB7v6lfRovKVJAEjcb+OKEHqKC3Yh3uZGPmwJ3J9u
ZucofWzadgzT491U4zrIlhKqjcKPrzboTN3TOFy6A5jlVueRQgvfZnQvKcll12tR+2I0G6beRanE
l+8YLBjUtwPhk+IbxprCnAzEdYlnWpXqkYvOg1oNApb0wl8H8Cn3D/b4arx2iHcTTgwkeR/OOYyn
E25yAML8YRW2EWdLVzR6Zf/vopFOhP+TfsiHJqwc77mXVPlSMydFpzpXJfEaPr3xfZ0j0BvPnN+Z
1vyTXaHwcjIXn6mTRaToSCc5NEoI3ydRDNaFhfhhMTfsgnVyIVrHR8yaI4mw2uG7yjjfgHN1OlYL
GX4GgQX/epyBaMknkqWWX/hQjgvVfb0Jgy2y6R8t8t0TELnvh5DZP+e71VqbECILebw02ZxW6B78
JYyxYAw58LzYVWCr2gpOGP0XSNx9BriHDQSrE7+KOVD597CcJRagqqUKhz6g8cwmAGTmonIGo0SR
OhkQAAuRboX5Z978gxb55K6fA6AuLfI8++7vqMN43D2Zy61Qdgu6rxJfx+Mcle2sDJMLfQgkoLSy
u3AI5bhLVcXwZFJyXKibwAbVqduzFAFvpOn8QYKJhlAF5avQl7CBda6cPmleaWWOFbO9iGi+2tjP
cQvVwWEl5ma6NqE3BpFbc+uFpxh96sOYQzbiGwd5XIknaEt4a3YtPvm+vE6OCAwZHr7U8iBt4G/i
WLmG2xpgGL4s8MNaK/ZBpdHLE7DrjcdiOKRKBEyKt/Ax7nmU5Z4M21jT1gC/v+YYQvkiVzUFtMvT
GYGo+KSs29BnymbYrX1sR7zBCTncomFGjjCy0tZKQ25Dz03OLMQrKYIJo2Kdeo4h2MIF04MzR5na
e81df10Alw/5bXnKoPKr80p8Oml1f5foRGwX+10pyzFutVnheVw7nHsKPs/vezvBA+inE8o4GhXL
h/HdflhWNZsmnj8h3+GIbURJwLTZ2RiscFRpQspySCEXln2j1/4trH6b6FkWMp5CpqgkpzF1J11g
j6mLfA45z4RAB9anAQqlppKKPtNlxAH+dqGXLhFjXMcEmchQ4km/ky31g1wLqHFvebpOvz9R+Evw
lxF5ya0jwF4DRQiKhjw+N9npwMfTyG1Fp3sYGCABSpUzqgAUC/eZAYpJyVhbgm9xnguwyl0gMpKp
Vfv4GHJukJVizn2u1oH0QGZyf0LKQerfcnjS0Us56nhvVllCgauRMp17xomYdIecFrYB+P8G2R0M
PhP9jMbhlBUS4JXohjwflbxVvx883BkZWWa/8AnH4CHWcFNGlR9TsW3L9fZhqqQNDyAK7pVtrdgv
KNObCR3ACapJ6DD3Fu5ZEjsrSpZmGqm5w6S5SrdmLb54p6JFzfvNlyA34wVyy3/ky0TipSxA3eU/
LkRtocYquuCvk2H42JvoozB5GJVTXA9J1BaLkBf23aky27/sklqpKLzRdtfTxID2gUEwgh5l59sv
Un6Dzw1oCqHJ/meyq1Mp0mFFIgzbGKgQcVeS5lbVTowje6DlAHlxGOCPBaOxZRGBxeEWs3mRDKae
nJWHyGla9kPircPuBAhxjSsuT1ct8DC3i3ViDXgtwQaH7eB85lVHeiKCuyncZltPiYnjZEF7UUtw
s0Me1xERI8585KxZ7K6Xpnq3dXYIi5B2FEcsRNZwK9dFu5MEmZtt46IhZ2xu2iKQTn/34TLFZ3jx
CjD838AzzX3Bvsiyzvy0Hr5gVLpc8VX342qUOZ6ugp53mp4GaGzn21mVEbU3CP+0ukJvnvY2jKky
I7ii4sK7vhiwSNrPbPgz+sLuiN/mZ/fCgGccde9hhDLyRGOhxlvgKTaz+amUB0FUrbRR54LJ3siB
eomu6oU7F4HTh8X6NcMFwNgAL+eSjYbqKWFe+xd06g+Kp9zHriJ2v1NTohXKn19KqytaI5NQz1Y9
ABbMx6pyjwH5U1WTbxS8qTjNcLHga70YZOQkA+C4+KycbFFB/UzSNY3neCd14tS9Mp7tcD14FfSY
eB/eIgmLlgtQ31+Fc/aOvPWh1Tl0dJvL4J0cAaqfrOnZV7r4Uojoz/I2MPEvqbIMm2JzePFSOFe0
WewmAOmnvJ/qrkEPn0tnvKZkNN4x0wd5b6BvHOBd2hMd4xdtkGXGWQmWHy9WpesPKqv8PK9erdS+
+0aM8reWRWQmI2/oYwRF86SMuIAqb8Go25Rfxv7yG4TtOt8lInctQuaNXjHCCD3LcQG9NovoJHOm
y1pOoBcpvsKh8WZcqAd84S/kLoEZYQ0CTyCQzLKiLOsf9Y1Pky4V3GLMyV8XejDcGO4zC1FFazGN
kIvmZSSDlVN68b30BhYyosK5Qzmbffqf/zWpSBZ06/bFWEdeR8TQBierX40WAXoAOWw6dt/nilji
HpYRB/wONA0UAC97wUFUKf9fZ38qoqvnY9KnOZvl89FOAT9d1hZJ64tnUr7+xYjTz7hymaK9nvcZ
4eZAmICce774b7WNvMvTPpncS9t2NN8zt5SRYlkZM6CbPO7SkeuGERsnC4kKCX2mEGTAkNMJ2cop
L3I9qrBf41xhCLgcoaU07q7zTX8R7y2uMdJYrNwV22/MilHpfGUb5P8hb56HV/nIjdz1qF9YTzNR
kSU7vd7fxEaVGVdiMzkXXzy+WU+xTB7AJlD9lyml+4+Ta6AIGWPXc6RxPX8YhJJdL7TFWekl38DD
VIr0qi5cI3At2HLYgqrP1AWkzDQ7arte4vrBBw6NLnCwfdnrLffXcv2Wlt7EGa7TXpszN6/B3qnV
gamLCV11UdKv08hBslXDk7paJfoJfVDE+g6uL2mJW6zribxVMxRXhYc67KHxqqdCo89ArL51XZPZ
2V2EgJcPezJp499HOqRI8oSWEpA1JwUf5Vk2E571HDtXL/dHOSXKfADeDR03Ldd2Kf9+kR+JmFLx
J6u3ZozJWNeKBuUNKNN5/02yYqG+/ZIDNJZtWoZuJTSqD5xodMfL0jCBke4bDim+D8lCNhE977mZ
edzqdhBM4Utq7K9AoFxAZv+bU4ocCPft3xo/nJlgdP4JdhlT41AjzWF9lisqH8WCr6knhkemrvYr
Znvd3IKYa8ptEsK+cp4YE4ZWXS8iXJvy/EyT/J6RfBShitI2d3FGa0mENOv+55n77Ao2n/vwGdcn
cEHYb0uTPMSjtQTl+7vlEY1/XLe2+TL45OnmORWHKq5e/8+mfu0ypnkqLxsT+Xcy5M3nI28wsgOL
mZeB4hMBLCTf51DKST73oNCcMrKlfQ/iNtZMDpqen/7rnCKNTcZH6PBzk95DKRzPkNZ7REfXI6uZ
DSyGkS76PiJNvOwdxsMUYIzVeNI8/G+v6CCO2EZfhp88REVj2uu1ID/K7nmpZzc3/4bJkjil7o1T
reI1Dzy1wnyat2JllGMpIiVoG/L14PFisnGYANdoQ3j5hXj0NsCGQNL0ngtuph+/ifTTRXTFjaUT
YFjlh+q9apcXJFf9EPp+J45b6Ov+9Uq63gpfr/Jdw22fYX7lck8SR/om9snOvdIBjR8nJ3sZ2NYB
KI7+hpcHnRQHRnnPwvmQBm4SNtQhkUup6OECLKaSpHhLm/afM2Cb/uQdyjNqxJTA/PXCulTkCkwg
YmtzocMp742DoVyRQuBKyRrhAejnrRR2ErftSGNkXVqYptduj5ffQq0cLUOMtAaOean4ts0IU1E0
QqXFisKdG0DHTvG7oXyNQ0iZF3uGe9k0J1BHnLX50PVoSHh9/jfDHhr/9UIWUZjVFXKTWAaxXWig
AihQK1nllMgoow3Q0JgS1VjGJPIYbUf1RdGlcTP62/nM6Hp8Y6h2ROs9TN74YhYDuPt7FXZHVXl4
OSarVUfIf5P6OsF8G4T2kF6wpoVvNjJroFEhTvSqX5YPgxgHDpILIJyjmUt/h0zLyQ7BtCtkX4ch
kMVW1x5hzDu7LmtPFO9OxzYXF6XTJK7SZ5OCyWhpsLYDYEsCa8tBXx38QRXE7t8BtQKo0PXHM+4U
4iQqNl6E25dGIHwBjzdkpKEZNiUgZLADJLBQvJGUIxOVfAeoRgo5bp5PBrfEq64QyvMiY7E/18wI
Pf1zRC66TiXAYyLd0jujnK4Hkx4YrB/fc1ouzsoqZoNqNZn/Bgj20pJ6TiycELvEtTjh1RwEk/cS
6wMXr2N/cLLRm+oTyOMa6YmTPkB1yHgbrwnhtB5/9dCVqYMysuAbuOCrAzvCx8ZKMcKVyXpR89Rl
wlA3N7mh3ZYTuNeWwze0z+hGqKNYfW927mudz/y4o+JMcOvVj+xeRhcp8hPWC6tDk74MKHvNGRkB
BCiRditG7G2npzPK6wc11i2taWrzv1oWNQ51MpxpQo/mJSy4HvAEshPIc7pR11Ogou5zRQ995S5F
QLqjvxWhH49tKNA7DTR0pnlyiyneo/XmEoNeSXuWrYOqpT74Mp0kiP9k3fcYG0A5BFCBGEUAPETY
yb+pFJC7OuOBL8vzqrV9MU8fC2F31j2HrIk9dxtxLHKPljxUyxSqUjzmGTS8A35g2VA2cEn2srpl
Dvz4qk6SsBTF7IBtCbwAmmhloO8D2mojDjoa8OYIogcPVCyjwtvDhL9xo/0QdBISwFHZI8BKkdMh
05iM5CuQKyClDFyEzi+7EHCoFFYvb9YJjHWV4QGWc95ixMrg1IuSgqKopvdkIRAEcmoYxq1nvgti
DJgHB5/DRteJL31C9rBcUUqQ9OjgiAuGfpOAi0NKjimO9Q/N2z10XHzKR6B/8zl+NLu2JzglPETH
BBaA9PW5R+ez05s6UIwtosMyMNRhzry/R0iHALgbg9SD4xBPS73zD6FmlEpD5+jcH1gwjvGtAR0J
XRJST/WGsNOG/yeBTyrxr6s/EoXycoxdHF91S1HjExo0hHTd7FgUz4ibfzlnptIB5B3qM0G9FqQH
m6m7XHAC4j8vOZpVIbVhXs52YP+ObSg0RbpNveeSYZliHwwfpfOu1lhl5YPS9rn/4PJl4y7aLMSK
De4bip044XFBpAWZKf9fvkKQlR+LYWXVdjMX57GFhWDCea/YbKxhUnhwpHmuXofge4oRoYkWknvG
3EzluSoCDkzZZRITQSTLWPO8hA6F7+mQoOwm89btJMuDuHCufo9Fac/CjvVFJG+HZUdWXCbBdBO6
vHDsrRlWNBxB5ZuzPlcLgqmhhY7HEwfSERI0BU/U613Jye9SZrNUqAbc8C9VXqN2YGYGXnrQmLB/
jHWdP1pUcS0eoKQBd8yyoN46sYWqGioddrKA5lV0UVevWAUroVWvF4id4sy0xPN15Ryeoa86sujy
uiHcHuGsztBAfyTDzhc+cdCrTvQ0A7XPBFP57BIDyaoZwCtsFBcQouCBeWiu9ET78Jv7mP0s0FTr
Z9gz3U/C7AdofYtVZ7ViTvy2xjjWB9gEspaQTrE1mXyHrwae+0OUJtBRhY9miwL8ZU5is52WP7Ju
3wQ4Z3LZypFNQoybE9eIOoSRKgbAETs0zo74S49MTMIQFeVn8kB9l4hhtUdJgjAmUPsL/8mqZkSP
lvbboVcqTohbzkFemjbU4M4FA6plYOPP3JxOango5fxEuZVK/M7e7j+2Ap1sltfAblx388apCTi5
2mZ3RsDez3BbUH/qn/Wop9ubgLjhPPNe7lBhVvvocfuKjusESk2RXYr1EYaaN44Ff33WHbSdho8s
kNLFgxn+I+UTR0NcwCAlRK3j6UknUSMeCsAhgzOLKHfavAwxkAyE4U24pct64dJxXoBgLwa+pKyb
XuS/2Hz5qMxqHt3kh24gTx4SSG7nw6cKw2jOKGYJsMO1HUQL6ZgLbBQTBc6tf/4v3NtedhgChjmf
BFmJYiNenwzYyett81c3b6NCZu4qXIthYNWz4SD2HNpn991lgzWUR7rB+mPIwisbFi+ZbSIWwcrH
Ti5I7GeFyaNTjzDWo1hJ38FKRiXEMbbQUqBqyFsmzVmVupi/W4NlsagJ7tl3V+QJDTsBknQgBPLX
1U95gmvzbJDZNE7Ziu3AX6GwBC+2656pHhxunEFPi28AFkXKNKnvbmU2+iMHueS4Ttq/Qt5ZiuF4
2AfUkyxaQnr1jP3RmbPH6IIPwWWror7XKbgEM9FJ7tn0GaBbypGzeq87t4J2HZlE1ppvSIc9Cd8J
MfC7MFv51+X32WHzJJoJ52hpP07db8okrJVLaGf7QBjLZZxgjOEv9UBWq6Y+4cydnqrJcx8w5wTW
BEvqxiy+geaGuzXRVKilLzKwJvYpbaXZBbHE08T7SsICgiQsoJKnE7OSEqUfQGNGEaCwEZNYLS1T
dHFd7CaVH2UNM7HMXOZVsHrLAcqNSydN2oZbNId1nxKu1vA3Zujmy7yDI/dSH/eKFQRjP0rzMhZM
UecloRVvNJ9PYrg5icgGdExqIRSYHUsMY8RsFHV3eJyH0c51OHmQdh2sX85dVZH8Fz1XdDffEenA
VItivF9D8AYZRb0FE2CloQdA07hpRhhCmVVAjgQi0Nls+e53iIXU59DS7yolSKM73D2oPDEgD4CS
gt/qfvQcFoKx1+8s05Qagoi6iYXuc5dX5XV2nSm6LrH1dz4HZXhxD5NMtAP3U1TWVBnP5CvB4JhQ
v1nKepG1JBvgv7LO2ggpwH1mdMw02/7qXmW0uifNPNZ/sL43wvsBNNRsWSQNN6RIeRz1Fh/Xi5wz
Z2u3wgs/+x1uFf+x6kkjTQKTR0uZ1xevMbm3jKjKk9v8r+e8xcmZnZwU5Nf0o7o4qamVuPe7FwVW
UahEWtQAk5OI5KbbxJMAOI2BX+4d4gmyBAl5yQ9FOqO8nhh3FDowYpA7c29/uL/ZLio/bBGvBseG
SJ24PtKTavB5dyYdHY6Ly175z15UnI59VyWljleI7Ms87keQz3oxqZWPEUztnB99HL6ag6zSgpNF
KWF+oZ3//IoyBYtm325NHiB0hTTch1ZYbRWGxQxBfIzSUFU3hQN9zSq9rLgdOvSIOgagTnDtsHEF
GQ3Vl0DGx7QOFd6qk6vt+z2MdbXbpcQpgOUGdvSgNFG4zW+50WmRC2JMGpvPTC25c+hwtMRO5c7i
gTcJWgPsc17bAoe+t3ENL2FyJ6zUQmrCiOBafYDiXaDdv36/HNRnRF0WJV1QsnxAq+yMrevdCFmi
lDIH9ocSbquiLHib8TWT7tQ5lLomr3FsxLGmPwIOAPAq0CD0mQBarfiII65DpgtizfKzvqgi2mvZ
6cMC0sNBBGPtBs82Cs/2ZOhCU4FmUmsGXneudmQADswDXK5ZAgzF8vB46e0YBdh/tR5q6LNMvia3
GS8wrncv2pFNYyHq067cV2+YGhLSLGMEJP0a3p1KyDWcCFzqJ1VLJy1VPxpFKW9sJWuN/j+luukc
9+Q5ZHToI0daPgq3b3Uzn/3N0tB14cymu2k2++Sb9s7xw/zyc1C4pL9wkzXSL8pfR0APvNeD9n+p
rGH+hvkWq/Y0Pv7pUbUXdD+kDEJ1l/rHZGOSrJYGQMqQMCJ/GdlIxqgUb/Sweew4VsYRfoO3beXv
jJtT9Wa2ElgLfD0xHK3pSC4+8JOb9qyB4yj+jiRCOa6+CzN37JbCtaOKNRCXY8+r5TmiznWN+Uoy
P4KM5D9TVckKMVKxKMflBVTz7uYgSmgdUVwPLnBB0P8BghE+gMBsC+LSx2ptRD6JDuQQI4uZ0E+L
A3+jSzXievqH4W6gKQlwLmkvI8+a468F+e/mhn4lEXJwxHjii5ITgL6JGNAUWLXRBaShod5aibPF
s0DbsRSW1WWdJu1eiazf011iO32JKERjKX5984JKwDPspD0ZW/T3zQEhBFnpGR8ruaFLCVuOFchx
FnYNMgdplf09MDx7l+kDXW9hOr7keihvDB6DmKzcHedSsPUnJuwx/1jFd9xPrJ7cZ/DkwteaS43a
9nOMgLnfzQsWUEvz4nmLAVwqRdcukudqeqqco4KwzpKaIl9uYxljCdym1giR8+lXd6u+2Pz6x4xs
zbih+6tdixn7qW8e8+L9XDf56N0RkUGarVtd8L6KrT3qvdUhitfvPSEC67Au5SF/nrTT5TvaxL5D
SG7STPhTERQTwdm0KuzU2TZWAvS8gz4XfttogfSUC7Fs9Tx2kxqQ6YlieTbX4MSqOBGDb9ulUQR5
wvaom9eumLKYiiQLsLZ3KXdzZEn1ELeByQtiPUWoaGC3/jCa57Ug1FKtLaU3/HvBBhgqqQM/6tN/
5feHP8hLdnEiJ/04RDidXmyyTqZl3AJRCsAolx5K9KkAbnTee2IZ+EY7B4FrCizPwxK1lO2BcO1c
C0byabpAvFm6v7O6CZg1w3NTEZ/Bdhf9p3Dsnq8nWaso8ug3y5UjyN8QACgZrh6SDd+HQknz+As7
8lTKq5/5nicG4qSZgp9YDla00/kPcjxR8KxNHZRKcAXI3ugoaXleCQVu4O1a0hEo9K0F7F8LD5XR
eipE4WRXyXhUUaOaXVi1hMeXPSfTJW8kTt82hpakJJ6DNh8wn+lfB1+GiAxI0vse2KQ4+Z32hWWh
1Yvx37VU3zEu7wprZJcL0myzb0gPIlXhGihchCtR0YoGhHJcYFef9TLO0PcXYqWR3Oeb5/L/G3lM
m6yoiAHhhKZL4KBcY7+AZSZzzFC3NOuf85hDJlKCldNA+lt2W07o928TB4fkuSAZCTrOzvV+dT58
e0ZNJU63eeWmj+7DXCzhdXHgEwTcV3qosC2K9ugZHLfYCyl+Ve6VorMC2kdVHqpudZknnuvv3XEi
tH7DRS8yojxdnu44qJYfLN5vonCxFDljtDaxF1n1vLz4ITidneNmcIXAJnwi/Jc9DRSO0XtxKPUa
EgvJs+PizdXx/wz6Vjmh0qAGRbyEu7AwFB7oAh5wDrz/BHPNG4nMS3Cs6jUNz7kqQ9TcRK8VRfSC
bfA5U61E1vfRM7PVU2bPXPi1kINY1LNyWP9mF3BgMan4FsL9vC3Lnc9A7syClJqvqfpXoqxEr4zF
X9dxlDjP/N1NYQRF+5Nuwe8Vk2xfDTs8EtoQCTEaO/64LxMurrpQDGsQrlMG31M3di8LSa1new/Y
9/guAVUP/dIfWrdnoQ/cnrnyqBhrq66y8v+QgOMJEFW0loAxbwP877LTs7RhUXdySyfMUYgKwPPC
+k9Jl18FVVxy1f1nvAB9K+jTd55+m26sUOJeDUw9TCY6rsdZl9RsG7IQiflmJ2dumtGWD+65IkWL
5F5BBiCy+jSH+Qiwskp5wSCg5ekOlrlfu0X7nbfMWXl08IFFWt0e1YCq95ys4kj7rwHFv/N2mKk3
6KQ8hDgxBse+n2dcpSmdUaC5/eRS3NBRhGLex6uLbLnhGFBSVVjICxYhSuYroFBSSFp7c4xRy902
+WBJdyTZS2MQkLq7IXetfcPVh5WgbrWTGzehw/v3WuL/z1a0GIYyTEdhuFHx8ffXOfYdWeKoWgKI
9cgAv2IENw+ZBJIK38Do5uExooFUnVx/38dXY+vtw30Jd5FFwg9DdJu2Z/gqjf/1ZBHvaO3IWBXC
+3vq1rpk/5PrlMdXEY2EfedvTjcpNfM3Lf00OMkV/2Ft3buV/6BxI19YfVq/g0F+HFXim6zeaPzc
QLDBRnFmOW37zB6mdONT0+L2/9yJ8Zptpz2tzmoO97QGNYa+oi9PT0KS1VU03+Ppfh+8PXdS60QF
YB20NcM7RiJDKY9NkJo9aY1zmtPVFZmUTUumIXFMmSzM/u2BC4Cnxo/yXh+h5JaJQ/B5LQvGe33H
RrGDxNgIK2hA7LRC31RBzBtbLkxUafdyhcjKL0QNKsCoPPPE6IXJ+AXSkCRHsm/kPfnfH12t9FsK
uV2g0ItAxbPNoUGOQ+z3EVnMAJAUmFw41gKrFq3V26LDAjKV0m02Jm5Y6Z8z3W+unGzv+AQQw3Yr
Petk+G7UKy59em20L+iYPsh64F01m3frztRDDUTpdoXBSz3O9hGJtNHmrutvXezpvL+i4xiUNXk7
2EC9zX1bkCKDK7mwLMGhrFDoYBz6pnutzVbKEycwNJHVwFPZIw6fWd1AwcwxN4K3Sy+ZvxO3LaSZ
tOgC9oJCL00ys/ImtSKwCnIhmmi20R3TbDSdE5BeEqsstL3qRmOoD5ZnRLMYXUnTZSSgx0P1++7w
qhSxgX80D4ysTNQ2r22Ig38MHHaXz0uSn1cP/9Ce/5vJLZglV4PzqebkhbP7azwO9ezc2MD3R0Os
qyZ7eVTwBvQqYxaLkKTJ7wWQuMQsTDzOHre51+pC8Md8AMffX95+oqJUD/hJNgjC8zBYB6rS6TmA
Diu92wyuR7T6WZ6RCFWBf+K89aJ/tZaz6gE12e/mD/CpnxjIpJQySOpbWbWdZyiglYA9tfkaMNuz
EWMJ3ko9dkZUvAO7KwYwPOHwHj5EgtGt1mKz1Md4S/7jeN8CE2/f5+vmp9ox3JW31QziTQAzdzpX
6p4Ab+GdKwPCqOYxUph47AgAGqLwMfuXDpBer+ibX074gxLsVinIB+G7GILrQQop5xpoCjC6x9PS
tV3UsKjx2JF8ykrf9ghF01xi+N+slCRJmPRkSeog0cwev2JcpL6cHmWtrjBwKUyoqh0LsDjhBEzb
vH7SHb9SYfsbvUwPtibcSa9weHH2rii+O3VOZ4HmPN5IZ7Gzkek64hYXxe5NCaRtk8ot1tMAPElj
iE5GA5hPVv5tpElTBw23YrYuUOuq6vDmcd141xYxjLSKmlpA2iup7ZCDRT59261kEuIqnCts4d1y
ffwta21bk2WYIqL8Ses6eUf4DNGWoQFkA4TaMJQh8ukbsvojE7iYIB6NE/wxQXu5XCocaDs0STre
ZyBQ5aR/4zkhiFgIEHv440Gq+3P0rMIrDBQcZA34wd4mxg7mzaiVMHRnXqFH6SGEzEyN6I34VdiM
/4e1o4JK2EtvmSjkipkOhWfqqv+QiDljpKtdmPnxwtwpy/IOaGwnaS8zXnXyaMIAqQG4Ip0h8KiO
3TPOv7le/GcKGaDt8yQsX0S2mx6QqmJpQgrBWn68ui7P4ueV2zw5iM7OWpJphu32mujC8bBHVq/C
2v3LoBPUMWARVJFmXt/ZcDIaq81KdxC/v1avu2pa3hsGrKveSgOQKMplVrMNulBBuvfIVdvupvLt
rtEzV7v2lQYCPx7gVWVvWOPY+0TsY5jO6TKIG8+ychyuH5vrmuJqU3xus2MG7lK4vZIgb5dD4/Qy
lKXFNHbKl+6G0cu4m7scYB1FdHOArefJwvbs3kVXvxmwVkDIQ/Muao4Oby2Lpyr8LtD8Kr00Jr5a
hG9c9wtLHRbGvnvOcXJn8NoPDqHdZPZ4k9osgZaxaN+c2JB4jdO0iX5fmSBqSZQ+oJysonETqgaZ
uX8AG/nqzg1soYW7FYM/nym5wCv8smz4Y6wuwNyynl3PYNGWj+XdwBcPVZdyAirsnpwL4dARyyMq
0Mp10khTtWw6jZ8gKIL+hZFVgNgtWUwqyaYUL/bzkG8JF8UkveCKx7Ww+kWdgD+0qSv6EWYlOHhZ
bbB52EwZF/qrffNf4BGrvvzsXjaT1HL53K0qp2cktgZjD4OlE6XvgW7KhWq5TNyhRa1DfspDnj6y
hAlx4/G1sjxY+rvtMLI7qpi9ScIFIDUJuW3Yvom+TH911KmLAOjhVOrXg42qmNyZ4KDaE6erjNV2
t66l4zBWRsKn0prd0O8Jm5y8ZvLJt3OULrt7isF0e+uszzUwCzdyYUPSFbhVNEeDnJ91ZOQUS5S8
vG2qDEcy9Fua2g14lX1HqZS0Qz+0c66GBSj0Zge9WYCdgSSLd7mv1soJ07HO+oaB4v/6c18q/pl3
vjaBZs0M2s8BPuM0fQVPx+JXms7JXFZZs8WkxidT+8EPNzW3MycEO15oPbB6Chrs11zrSRIcts2a
bEsNkjn8cKJNOrWa5gByLNDsszgU8jAkYwdcnG0t98kpbIjP0fZ7W6/8Hgjcrri3EFJvFUAVYZEF
wZm1lH4bgGmAHtUmUpocF/0oEHlRUdos7uuH7ZxaXntRvRUl+E//5DpLk7IZc5hCYKyK+oBKFrf4
vAw1v6JyfVZBixkMGPeQoyQ/VzJn3BDPC32gto8XUYwnv+z87xz3oHWbaDw2TqizjjxFa37qiozs
0m8UxHw04Tk1JTFRM5OeK7wPfFgWBOJYny1kQ8cCDaY9f9y3fWHazn3SRPS6llcEjgM4z0zJRSYT
Q6VvyiOyyDJqJlJg496hjer2Ko+vmsONL9VpniXU+XA323WkpomOuym6+Ymj4K1w5CYPg6qNFxdx
b06ae9cabz9KWFetUrT2WSsWtjlBYSLzlDH9CVH+xAXxcIF/PX9zYs0ut6V+mWYu1UFpeYQBDrie
Zj9aCGRdq+VqJFpj20QtSMXPYJzY2eo7ItzIox6eZmgjns/ne3EDE4atjDF6iwauLTNwdI6t817s
Yn2yNQ8aDjcsZthpjLorCl1y2ItMm7xSqbj5MOdupRsd3cmIcj0ppajrv8mlf6CLtc5o955E4Qvr
kf2IWk1FnHs6o0oG8piY3bu8ev05aGMbigBfaNzJ7OEa8xphxxzxOn4k1nyT0Nm0XRPYomDPOtHt
qlGgJJj/sHzNOalyV4zP73otaEajTi5d6IQzlRwM8Kyeuny+KsnuBiAoYoowahQGD6OSYnAz+GhT
PxP6L0NNASmrt6DjoC3UsU9w1dNDm07iLA==
`pragma protect end_protected
