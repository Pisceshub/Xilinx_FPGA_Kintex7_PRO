`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3760)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEMIY9k4JfhpnaMs2WbrOTeH3MZi5wwG6zm9AZe4Ng+UTOxxzVNu2qggL
mFWIJ2NErZcvu8WDrtv6iaiTNf4jEvA2EDRSA5ni7Bi0k/sm1TAKApZQxZgX9Gcz5UGtm4YkGWMJ
q0Y5S1VoptM6vo22g1j24CVCLz6iiFCOUICwAV0TWAS6nbUdRyR3qarUl/UXjpwaH6vFRl+YjSlK
DEELUE1lJhnolDbqA6kEnwuGTG5HQ07bLuVvh40ykqDVJLy5+a2LEGQOs7sjNAtzKrT5l7niF1xa
7YiYizmNx226VvjzIr6i4eiAGbP2L1IXnH7kIsxuUcvutD1N976oKwse1PnlBA0Sa+Aw0YhogQV+
3Is8T61cHm17Uzlxxm12GO1dZyTrD7DRzIn89i9hdxmUT5RWZ7N850EAHFw33zeEw6Dgo3Nesea7
Rd/MQTYR/vMZsY0kQRyR2H00pUbaWuPIFIRFiemaS2I8NHwrzS7I4rqiI3JWjTQ7/2/Suyy9CnE4
mqaMLR+3em9kgTelu4VGxnfP1ha2h+ZnoCG3RUMuuH2mkb5tErNUIMrwa9/OkKYjp+boesqpF1Gl
5RNb7SBNKX8kaPfnZhE7D/O+iopJA/wDMd9bReYbMf4WNZw+3qZF3kaqE62WH4HacTQUXok7+6S6
M4tWhxuZU8AXiH+ANayMmvNMjxkk3dDGHgYuDG3tS40QeVj+Pjv0g/xLwKYJ+ZieZ7eUHf8qIrGs
5Q26TqN0jD6uxB+uXNZPYT8zgqmWlY8nogSMo8FRy+6rCf8wmE2yt7DR3C31q/FomFfe1SwUBM72
UXj1/q613rAkpeXJUy7ZsXXbHt3Yizg+CwFDS/70t04PRt+u3iIv1PGAWAUe5DRXOS8AZJhHd8dO
bd9K4iDAv/9dFS1B8eYkltpDzY2jIRoipr/07s5Dp70VKUXHoXHe5ASVIqLhGczkNCE6qU+ZMWme
GxFzo7PkMfwHqn346GvatP9Bh2ZuxcsU5LMlUd1YZLp/EAdpdK+Sd0Y1T5XV/ltyzZSeQslS+2mc
0uhDBQCuRnGzv8b29ewt6po8kI7d2VFCQ7DbAJnpLwfXx8H4Pq7/uvVFMui6DP5ByHTu2Tow+msl
p7JUd/huzCLhPTcSSc3uH3vA1lLwcrCJ36EV+2QaYI0CM425VX4EqCaDgADV3ohgMR2MM6H/Vd3C
sIsUWNwjsWLMjVY56soWwKl5LBV2jJ1645wMJVsY162tft9pAPNOmdCnNySOnPfOUXdSrw4vglj3
t1eB1+eGJ8DXz4ydMGwsUYdS0jnFNA6hMr22eb2E/rgfNdQyU+whqgdgI5ig8rXO0TOEPyOhveW1
AA8c3lk64p5tjUjrGTv046keTQWKIFn1FM7f9Cym/KexgYz6L4RAbXUnzjV5K//yWN9ete8Qm/Iy
uUkH+x4lnutu7wX6o9Rlt3gzDY5z/mZiYDpJKNyK8GEXAPKmYQWvNP31dHDd+5+a7zPPLaK0W6Ls
jEMOayzd6SNjRdefYzUvo/dqlYIVQaEbVYOaVjS0IHzqmas+Gwl2qFDzRv0QDKjPDzigv9I0RsEV
rflLHgtxtFiauuw37nLi/P/NlVjn3E5XnTLPGOxtBMAfE5yZNKsIunDOgSyOzGoGptjxOuwlazjT
lBqw4WQl3BlZ6pc5BiaxkroPB4XYRf6K0htu+isLYJaZXIxnWiduIqxLO59XvIe8Um6tG56upkVf
6Yy7vA3W1WAjPW6oQNJAdvLD91LSmWFDI0hD/X75TX06SRuCK+69Q6xTzI3o08sp2/gUjvECbIja
YgmI1Y5CqTLvPzFx8YO7q3+joa6QYKMFxqQqWI+EpVgOxeRctfmDzCmXrcfuicQg2p2keRl70nbB
O6xT2224Lkj+n3ZvSMMM1RzXY/4o2AsCmFrbjQA9gRBkY2nBdB/PJDIc+2AO1X3bYsc4C7TUhnhj
gYAuZb81Mo6vu45HCFcHQe+3nJQ6yxBfceRMacKMFBjVh9c1OGmU5i5IMqJw5KJrmCF1vNWCdz1f
k52+St9wGcdS1AB2HZ5dumcIN+/lckpXQmINylQkJUlBbJ2Hsz1EbNpBtuheGXOnpgtrvPcgHGve
kmR93VAr5l3BXDY+u7Ryf21Vn8/AUAEz6MqI02u7qQyp1OzrQBIaBrbFtZaiBCfsagVupxVnAk17
NL3wJNTlm2q9jrQOznUeExEh5QPrkT7Zs31+ibFfoF/ykk+gdDfVHY8Zti9NjjDM006xtLeYDCm1
noOC14JzcuxIlYXWx8e8UfhEj85vJSP/536mghtWWf8nja8LcaM25IKEXzA59muDUlwUHC7SwmB6
lujaY0J5gBXBjCQyEh8Vmw7ktAMa3IjlTSI5ILbjCpfGyUqTDgqAdbnZ1O01rVedjJItKeP/m8MU
jiM4gPprAfmbPs7iKrXPPy8ttiTY09Wl8wHEa241bYcecqhxQGhaILrRRe1zvs4ys13qNM4KX5jQ
5CvkUT966t4UoskiL0YDwf09aqo5lRfQo0WrZchoFsj7oDzjfS3QvjjQ2GKT9Uyj4d3vnKsbmTGq
Dc7Y9v9lNKPEAjUyPaif493bNTGSsjLb8bKOqb1rtUNDXYU8J2BkLXu3gDaacp/UPUEMFwuyqxom
ph1z1CRlOimJT64i5bkpS+VzmXzZeDrmriUsytCgIE/c1IIW/zeK0rltPKsSCiMf8gcN1Gko5KUD
1ZaiU0reL1HbDSUKUsBGqhnZ8++9mEwRbPEnjPvkomeFrB47Q+sNbdNvNWvzS8SmP52+76ANsAA8
BeJPFOKyljy3M1WafGYinO7uAiZ9gy7/djdL7o7sMDbw6QpZS6Z/BOfY3jB6vieGSFbLFOyQxm5I
/Plh8TeNWvKWGpQ6yRtIvRDuo2p0ygGzVtqzKqNIXNc0hJbCfOmCMzCH67h1Z/ssHAt5+v8eCG16
kgXbHWUYv1NrlHUOtxkke6PFLcSQuvdRzxzXCMFI6V36WxZ1I73qbTH5sj8LkwvxdbhBn34OqMUi
2v12/ejjfoPW6hPZnhA3yeosGThWwYkKYGesKV8frjnYKQcrvL5amWJ2LKnBMO1QjMqszgx9Sjnu
4dckhoqRnvqmOYBV4T56YpzS9C6SITC6NGfAcaLzhFxH+Ao1TPqH8yZoPLe7ty9klWAcrmrV9slZ
V4nHRHrdIW42RN/ouxOf7+9I8AWZgOY2ns+w8If3TngXU7cZ6CL0FrFXhS2zMylzgBwqT3AhTPCP
EM6jPqaGyYJG9vXe2o/zeZa3YuuOhw8etLFcOtHvBrXv6vXEvNVqEyf2Hm6c41W3YhTClRNPreNz
KHkP4M82Zi/U8hhjwKpzSUNw6TXQ0f9+K9Gsut2sX8CAgY6bRkBWswZIAwJtIh7FlsIDWVmV/uzU
fzHqb4tB+UklKcNWDQIB5pfW6WIySJlUx9kbxL8PN+tiGnPURLeQxf/lqE3fvNYqxivIm5q9xkEK
IWrRsBv3B78Bv9p3zaYtnZt1JH5tp0qq10OQsqicZZMaA+dtSJfN4tWV5hY2mhD7wTEBAoExpiUf
94nNSQl91fNNhpBcSNxKzsRWXhfs2Fjanqx/MCYyCLTAjKnkhak1MRBgFSWS/4kWbwKh0Qzodrub
HC6JW0WpE/4IdXpyEtib2h55WelkXL6hQo4qem0vFljzxow5UBeUIq9klufbJLGbfGEtKP9xDzdg
8KMMHp/8ZckrHhKz30kWauTcoRVySEyodruRMcfj5/Gofg++3KdRdGZDbB9veTc3t1PKlj/UwKYV
SNL1ZO5jz6YMhK8OknPuWcRKMI66OJL6fnSPk5Af2r+X7B15HWEPLzQEK2zZEBlxivhpKyk3e2ZK
V3u+Mag4+r1tqqKH+WIuVSwTaRGoRiUnyrptmEf5LgV97ZulYIAxpaEb86nmNaS2zEU+9N/xD+Ke
8sNR1SwbcG7/2IKzRRBHTUanEHj6c/1tk4cn1UDqw9dT4g4dXUviIVpv4Gh9EVpelz5K5K7DsmyP
VUsPhQhdj0sBTHwrQJ08forW932JnUGOTUzuh3vnDp8ZYMEsrKTWPT02PhpBy33GTzjDrw3lI9fH
OZLvkx74wstKZjPg56mUvjkXklsIs7U2XmkBSzvz/YEghqlAuF/DsZbiXdJJ44EA8tPifE0gT3ld
NvW99j/GkZ7ZeG0P+ERilNAIhXbg8IJqWWVZx8RKfrYYPxSpEJcmxH33mna9b5HF2y5UNiXM9XIb
tD2KtVC6h1QLBVITlrIf7zPHOH3HaI5wJw9Nh9oSFbkWEI2rfqUICugyerInC4B0eN8VwCUsp+NP
nQYMfkkigICplERk71K/SFBTJSl1SRbymsMt2Z2ivuYlrgsDsdT+o5JH9O5NEoxX+w7KlGvhVbHx
w3Z1AV1WDaYlYob6OKRjlr9fGtBiWD4tudkLTWlsSbqndTFLxqyHrWSB8l8kpTg5ZBmVyZ98Hi6W
JfXuNf4avZc0cBm9BKyp4S+iU27Qyk0DhdHBREmuzF0DvhsrNyL/3dAX97/Ncz0Aot9hIP6W1JJc
eGksrIauOH9ZkBq58nYF5MtL9BiiNzixm88ladApkomhEem0DHLpBUNzM3Dom/QWbJ+Fjf1MEWlr
0SeRzoZYEGzKcDk7pRvQEs6Z2VFK/QobzzFizi5/pNqkYeSHDou8g8qbhciBgaYXmbNd5UloKWQH
iVM+pL58PanRPaaRXJrs9mazSeKxmZedbtdBsp6UmCYLMup7N2EzGgYEjdBEQX0I/67nuNxFFRPW
HSzjc6FycBEoV9Xe16YzG8KLjetTQABQwsPjGH9P0Zpx5byavs0F4pgEyBdB2dimWNrQi4vCNJ92
HS2YdLmYjy7z/spf4cSkk87vT47ftsLoY0Px4jwEX3X1fqrhJ/vPgx0YZ+GfU4cGTOfHClNrZ0gT
QupKpUbdwEe2A2v4GcLVblKtw3gdsAuWnoNNhdQ9gAiMrFJqY7YCjA2Hp24GDblEGG3pwawAUQ==
`pragma protect end_protected
