`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33728)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9JQaMgpupSUIgDmsbAQQ3DJSs3kPepPm/ZZz3gmd+ukRNBlIpnkcOXIl
gXM9+wLGs6bJem+o4GuXn6si7dvgUs+WRWVole0oR8eGTY89US2CXt3ez+fBAep/rhlMK4nVWIIi
g6lv4qo91VkXmmfqGsuJnESRrv1p6mqItHizPBG/mCWZS7zk4IcH+TJPfWWm/u6cC3AXqQP3tNw9
YtuJqm9AUftbrfT5UvsygijmQcgW5eJgpKYrEtR+XHByWqtZdcERz9yohixnj28o63AVXmtunb25
bGMPdR6vdvmYcByrvBkpbMoL5qUKZtKzI4eUKSBJVs4xFzQ2sjFU0zsAVWjMWCCHGdCd29WuBV5P
KV/lMO/JiERawSSwUPktozMJpjHpSY3Vd8YMUeBR0q5jIe3+Ay5Y1FDFdOuCtmCvUQrVxbPp8TI5
Ky+EyrZCXGaRIVJJmu/pohhpHTbJdO+dNiWojGeHx/E3w2k3jH9NaJSOQbNdSDBs2eyOEg1JokD9
OR/gyNfJZdxuL2bH/w3bZQMPxC7VV5GbHxS+TPFCuGZGAhxr4QUM/gE9Pquo7JEdiOxq0X8GG+Xi
E+l+KGM2uILQTAy5VSzEczUTzUS92I0my5OFBRi9RKHyD8u22Aeqcvh2NqoF5/P6rP7Ubyr1iwUW
taMOpGVFn35xBCmuhYHAt7aWwbKeO3jxDkCXcQB1jfk5Maaq3FKUk6CXc368T7zoFnNgx6pajeIG
DSt2InpGa5eHYunxoZHqXrV8b5/ilDqWO6DvRICXxqKkbC3r0DE7YcmUzQw8C1o66TqcvR+xlzpc
uwAYWOmrjyKnV+2jigEV9cAZEzV6NJu0KmWIBo9vgzzTiBTWfSCTS5CNro0Ac6p4QmSWhzAwF3+9
RtnREEgj5/+hvhS3MGxSCtvpfvUm1mIG90mM7Cb3vP1RvaNaYd9IQpqPN7bLB3YHkGu+J1j7u8gm
LC0ChXbWma5I8TRi0jbd769Ag4RtUqDGcJvW8m+X3U6qBjnpceWcgjtpr1jELj9Qu1VCbt8wc3Y7
hcEgrfPM/1iXJiyM3BlkkeBbYDse3XnWo+OdufN/nM5wDWsFLrNH575xJqUTTOcgsG7+1THpEYiG
blpJHgBFnTRSe0sJR9Zz0ZZ59Ll6oi5+qsQyRdecUqrFNISnnSHJzlXZ7MT+OsHPlJCBzVUIOs5v
izaeyniU5v82yjfNnVWmWXMWlNC8P9t5iVDYak5crsEqbah9ZcYnjsSfCzKhAUJJBd0J6EQx6vV9
L63hQ8lzPfu3xkbejJ5hKVf3kOjSIdWniSRXsD/z0cXolcfcEpDrAZbMlKiJTCSuX46Mt1UAAhK3
yCvc88LeDw61Ad8lpy7a3C3CWeBdDamQj/7jG8bVE/TPGVYI+RgHYAS4NxYDXY1kohp67InrB7TB
8vdUEj//nBhprSazr2al2Ntx01stIicrXAlaHRFGO1aiSYz+EhkXtIIGg90RGskNbk1x5G3/0Sma
aRWUFuWzKPR5yk4N2G0e2/CIcE+TeIuqcm7p6/XcXv8GRiLV6Ndw3EtqqpcWQWqIVbXvOb6DJtzl
5NOxh0nB/EvTlnBu8BUrMhmxbndgqQDO+jOI36mzZiZbo8b/72K5XMy6w2EXE96ynvmwggXh2Dh3
w69fn2qGfmtNy8LQtphsJXuW5lxsPIoP9JMcuofT7NqR6S5fkBWBdCe171h7x/0BeP4LOCdLQcOg
3CJgS9rDZmIYA2VAy6SJtgRb+x2q0uzHovPDYJkEWA4qJOCa7AdLR+gwzlgDXNSXITL1WR7PDvsJ
TST1MzysfhwVX0ZmRkBQMBQQ0m5C2G0noa7IqHuDVpTqvoLhTXrNvxKBDRwjIm6icDNwp9e14CHx
RV7tnua5fe+SRNgC5W1UBPT6O/wqawiTDrQ+47gtC0GtVJwvB9h4XvyWyfg8THOLkA5S1LhGBVyb
1qQN6hZo/27Mx3qiRx0QA9KedUjg0VgIcGlvxQs3N5Z7yXsTRImEAL4V31UFMfGnl8BSaUAGeINO
pf1l+tQ1yOPvKR9ExfJ3KfJek9qbX/x5GBpcr/2/5tRXiwYrdQ7s8kug39BGpv9yJPNoePEffLDK
H48MYsCCRLbQhXpod4RoezvMRBZ98kNjCpNATEdknZnJY7JyprP112/0C6SsDsvEjcdOhudap4Yy
R/qJ5ajUkGPVH4fepiEfnYpYNSlyGMiXj17RKDT5cFnuKOAkQelJa8UpmxMSPBxpge4JSF6Bjvkn
cjmo2hi3pat17x9uWtmIrllRtet6KUmQ/COrlF4l6GE037xO6eDfd/RsGA9kZH8H7Uxt38aPTnoy
d3Y2cJs7IvTyp3V7f0UDhJU7c4+E/XZkB8Fg0Mm8LOmPS9aolve8s+7KV89m5QAmcV1KBrcO76Tj
TNe6PZhFmKB3IJdAmZArDfxn2p3RT7ZbDGgLq8MtVDzEpSkogCFtsgBUmhLgZ7IugxqgkJrUiJyF
EPcsTnFXQn6luPxq1CdWqZ42z60R+Pbd22+A1eDFbThTUBIbOpBBBAIqRGtXqyifD5y1gYQN6OCJ
/KxWHOegciEZwga3xsbP9bSvnV4v7SzCE29wyc/CALW0/nE1B7OyK/svCH2TOp95zb1xaT09ewnA
vzjHmzlmdRRQNM77AuZwC+UBWmvR2h6+OaooIXflyc88JhbjDSKmFgH/DFF9kS9ZQqhNhRfuBWhP
KSUIhLGknFZs0n/88BEmAnFezCzA3ItkfGuZs6FYrAWbEMk3twJZF2fZ26+BVJzVSRQ4q+nci1qG
/qUiKuGv7z9Mn2NIqtcx1slhRJ1W1+MUY6FCC/eHmf/EgiZKA0hdINWGXd1N+2XGcO2c6vbRZ1+g
a2YFMvxOGhE62XdPdP5YCnT4JtDdd1wG1lB4WLthMRUy0HbmD+GfXBZYGpCuo6Q7zNa27gWbnMYE
AKHAIkNUOgd2SmMO80FUTbtb/Uffcdvg+lq39kjeAIbD+08ycQ9miSHV5sB1+OaS+ZzBmmh9ZErU
FEAZccDrQD1fwULe9Ln916oYzIz56/U0b2GNNgqu6XCh9UW+L16J4x5bNIQfD95CoaX4MYh2dA09
zJpDh8ABfQLnKuz3FneOIzzuPjCk6nOepLiaTSArQbHUAZSZnWVZZ15xek/YKWZyregXzAM28Wad
JhWO2Hetx6WoYrN/Xjx+9hFW4kZGSn0ibUsnASM80FbOc6D2AT4agBQ2JxriGQzLq94t60OpvTyz
BG/iZHcVyhyuKodUKOJezVBSjtPTyP7TNJXbuB4TGyBQy0vjSbHvW0qu/GVwCzoQSlmei41NTgdW
nuv6r/uc2mr0yTrDbmA139k4r3xebALxjRWDxK62X8Bq2G98h/84W/DxNFgxFsveEyteVgiVf2Hq
pGa2TqyQwK+LWLAMjr8p8fdDfkpr1PcGdp992z+nysxLE3/dFe1zpP9olxtmRBkSTpy+BolCgRd/
9yVtmY8aQt8NzPRvkXb+kzKt6MHW33qFhI2IkmW0nc3L00UXtLuKQc+96+gbQRTE2sIc2B8R5vDd
1+9hBrVSH1kTX/xGrdC2yjKDpIBC0tzv5zT6a7h3QGjKDXWqV5Nge+iWRs7O7oWB3jRJ8kUQjgOp
Z0nKaCAaVFr37fwhz/9IkkFXc9Z9f+o+chJdoR3w3ObbhYcIHXySd4QWzslsF+l3/ot40njtGT8R
bfTahXAnN1Icht/3edQD0SlNH1p2WVwbegvGiS5fLe96dRGxULHg/Ar9FuJX/TqACQwS9WSJjMiy
DitiOftzdWMKigoM1MT9NjrIQEO/mliQ0cfRGGyiS114ruQdAPaBFjG11ZcsuO/EuB9JpmbgNA9T
WUwmQxjBN7lIjULHAl8rp3kfFaQE+HPPKJQdg4RPYsww59hwPDuqbndFR5V5DQ48tLcOfaZU4yDm
jN0xxswo3tTjPyI5ZLPUyR7KOdFW/ozsLiDv/Opb7qZ8q3vYPl/tOnV5WjYvpbcy6/YaUERIa372
1cvYUyYQrcmJ/QxJGFfgRTPXBewURMjs40mxErM+/BIS29EoJzaLWDueqda+brJlK+PeZ5IyqrCw
ufcSL86P3lAmpv4IUUy7c5Oqy7apEuiwYjhmT1Z0+7DVEgAvLP6vCnP6zXFRn2e+shUC4RJ7f8y0
wDIccqlOF7LP7mtORlkjFPd/dXPRd5ZZVtoTa+vLwQqj7hLvgCT+X8wZ3DUCBFHBWQvhFoqPrWJ8
KnIugM/dscZEfwy2LCxLkAiKSfhZBnW2XXVwbAQ6PFkw45DpBmnLIfkTwR93HJKE+VaGaOg/mOTD
eoWwTc4yz8aZSojVUKKOj3CZzQhQUnUpXiEDYMkaCEK8sVDHVLip9noNtKZjm+ETt7mqNEVSy6d0
6RyC9sCN4OiAFdsFRN7Q4VletvQYdtvjrobZ1tzQa6SUdwFYoLF70EzOf7hEq5w+7oVLOcI/gpIo
khv4ApeI9XStxyuI6QuAkSb1qh/rWFcx4GF4LKCB8vgWYUWu0PKUre8Sf1WYZHAOA9e3uS/2Xxbb
8ct6+uyBmmJweQK7Q+6f5SdLE/XhYn6ZCio3kgUBXObPu2KejV4Kf7OBEIctWBxu/rfNMQHOG0cp
KjZgcWv8Z4Ovwca949WE7FtfJPr/PCRGTKiwj62VM4ZvhfQQU28Ngw5r9I2kbw4jIfkB57MdINMQ
lJEpu+UXM0Lsgng4kKkiH7BRxdbPBni3MxJ5XorHBhbL/yYoGRUSUpL18YFPbs7kk098JcO3uAq7
XArAwCoN2SJqUSD43TY3/JcX9GziL40oQdbQpH4BkEuKKCLeB8syRNzTQ41fF0/ztfhfZP1flVK1
OF0CYG4mlZHzJuKYkOze4/9OWG2kNOszmL+0T8XkTsSZKTbFMdAG7rJ/g9aIAFxOcOWxWUE39fpG
zKtBWG5++JD4By8znkSdc6eJqWhETlACPutmGZJmNO5eZPdxIkFcCejMBk5gVnjnj8dy+N2h+fsy
GucvstOsPYcOF9TkfxBDEd8Gn+Gv7LjYZm56jm0b6RCVPgHCxLvmk+ZMtqlaUfHrsxPIpgPcJnno
UuQ++QZgS5MP9AlKs//XK1jCXzmcPip/ZTyscoBJnBK00HIVL25IXGuqy1gQt9NIM++OcBNsnaw7
B1eUCvRF1XIxkfxcb76oX8Dep0/rzPOhKo0lB2M3Cfl3kVsEBZlw2XHq+m4obxBWfpM6ueSSUpqP
Tg5yOyLx0d+7OqoOKauhqOjHUcZFgHpVlaCw24TTvdTRgm242FAOD36/O4lFb3fiN5g3IJ0kXuzW
usJCao4qfUWzL7E+JWQCgWW9s/0Hx42FjN3Pf9tecjCDaLj4fvqz20llL+HsegV9OYjO32nap/1K
HKjWTSh4xtjJ1Q4b5kP5pRiUGF/opHQHQ796I2UkIks9Ma+C0gzlAt/R7AhWvdndRxyeNJqPCtT1
KffjVh8297ZE34qJ2plhOEAjqWHSooyJhc5j0GaS0ntb8c1628USNBz/A43/KYp44VDuzZMeDQvW
iogOWxhb4RE20JB9vLW70qjO7AmTXkssZvl0+BlCtNFL4DWpVObkPVvxXWAhsv8ouRbWExoWE7NI
TTEbkNTuFuo27fW8LKmjD/7xUdqOknB1vvarfD4n+abINJZ9Wydo6JPnBbPQ6F12UD0WyZbGA0Uw
nD/ZfKCgTA/Lz/ZjyQxjjWFL254p/5MGmmujc5aZA9dadmFAkY2zGQG2fgx2h327kGJYCtXQnIQJ
+w2cAPsb1n5XMJwtzbtJp2vqXav2rdqdKWVrnIRWIfEFzOrlLJLEEo/cRbamgzfky/2w+CAxS/Nt
bClgz4XA3pzG4W0YzO+Kpt/sGIyfU73uTSMGCgVQ0YMNZg+CD+4n1U41J/GLszVXRdMy6kz7/PpM
yyzi3tzIUp0jHNBbrjqTbL+IfsefEa5Ml/yQ0up1e4ZY2lsacDaNsMM0umYXHQgIEI6uADXH5cXa
EulvC6k3w5ElxQgRoBAlWc/1F8DFAr4BuukOkGqCoc/hCZ6lzDgoAdkQjJkJP5oCoay7OJdloSOY
UO6XFh2X9ytd5OeYJgMKY+nHtIeRUYhnqHCZb95N2f3IA2FM1vb+FF7a25VZEsE6vCGoZG1Gya8P
VFc8SgE/8zfrDc5FClLmZTbjv4ZXpIWuTXCfAtdA+kAHwGJYzHtSh+Oho9htlHeUB8HIUGiHB0hI
n6MjCD6lvoBEPI188YC/97rYtJEI4FPJI/2yqHBQ2tTX+di0kGjiqVW/KJA5EQ72f6DiX0WKPhpZ
duA360bUtfFpjnj4PRP67WVr1cz0xUNw1TBCaJyW6wjYMp12aQh3OV9PsJuFkj05r7qQ8iRY3hMX
R70ripdAERmWQOw59E5HkMCkCowxviF0oXjBTwpbId9yc35983qZaAzOP/w6JX3TV8bdM7PUcq7e
w+fc7nbif+EJqcT/QJYkqrdlbXm86aBeIKNiCIGjDGoexA48wEO/atz62jqh0bE6HrcjC19tyVq4
uYz7jgJpFQGzZTGxmWdb8HZcb02F3UvWEcu6SljojO0HruNGJTBY6d2JW2cqFMknG7U/tCXr91in
AqK201VR+CM1GojhUI6Vv63tLtmJT1byl3iGY8n2GQSXJKUo3iXF4Lob3UfM6260+VCGNEILJypX
op5QXEDJkfkvgmET8/XKCEP1pkilROz8d643R7nA/H52Xf6GYMkfuQ2oMK2vxD6zCvswGkJJhn7O
oJKO+uqXlpBDHw1laycD3zxa/PTefDEYE24aICDo3v7hv/IYo63OXchvZ4AKY5c1yrtqkSJk8iyF
NiPk6SPuN9ynDVeLDVjY25XWWPVE5x0xBCMw3la71g5raiBEygaFKO8ujuHRNvwAWadhji7REfMQ
CROyCF/tP/P+CZL5ODOxVD04IS8zGBvDpIAODCyaX4MPlIwLR38av5BouD+JAjXU8t9cGjUz9qYv
kTC0UIEyaJZxQYZU7RB9YXFKdFtYsh4SQEExp+R908NFNhFUeMh14WA2Q/HYUPc/hHo92UC4tS/U
YP0PQRvADj0gxcvQvoNRG/ioBjz67WiFDSxwno45tOkfQzdyL3A0e5GIoJaA9G680ngvoLmGd4Sw
PMGXmvs7hvjnbWGq+vOi4UTU+dRLy5z1tDQPukUKLVpZukqAnuRsQGTYF0nxI8J+z0/DWsIpdMKn
SGTnwPOVPhVXwxhXsKJ+NKTY3he/SoEhyrfx/WWun8B992FdchtMhedKBmIXLQByiAW9o+KuSukv
Nwp0wtc9ChpMGKzlfEqKns5DNG+LqkP5zkn67PiHeXAzvfsr6HGqJMjmVOQ5L8g6MoESQJjBXrPB
6jLrAHuCbU4oqiZm7LcDZiMcRefzbdf4EsxfohzR6sSfWZcdaV71Eo0jT1rdR0SVHdw69RW3rL8n
g3I4gK1rkoWPyGaX1H8x3mA6xjj0lfxTlnCvHwc2MQJmhAq5LrlrMLoYQGZ64Qhy5RENfqwXNcuy
pJRF4urforIPeoCv5VdfaBVR+XgCmuuEACwjB7zFnVBFRlPt7lKd3KA4lWjPDiF0vTyPsuS3Zg52
RNBl8XKNEKrfC22Zb3XhTEZDSMzv9Gcz6AHR4NHf4fuz2+POK9p3fqeUJ/k9CEICpjK37B1nvhMT
po/LfJxqMMCf97Sm9Jd/nEReaUNmC2MRDajRbDaTUg1D9zWRnjS7l1Tqb4ykvW9tkTr8Dd41F/VB
i0sRi3jbUA7dbgoRI37T4ozF/DbCpmFzwkfggDBAWUpUHlNWNJJho3BprykyKZRp9iiIhLVRJb55
ZWq1FtuX3yDbOYz+dR1Xy7PaQvwoKFBrH5ff9IRVeJv92oOVeBOiWmNiuJY6T07LETpu7fxEZe6J
B0Z9z7BZ8DGmrkBr3aS+fNO1RW5q0/SLKMiPpvBAPKfkbdcHfrC2PL7IK7n0pU6pNIfHICCjGz/k
r7IviJ5OAUsa8+9W7zYEAzuJ6MASFzvTVJVjZyn4ioVJUZVypSrYoAyQFF3InfD00r1fnZiqdT/t
IsKkSjo2pD36K02YhiSTeUmNpUyqCvvzUMLWsgTA76RBkFGElfYcEaF2riY39uywJfFx0EH9iwwE
dkvhn7HjcmsjDcS74JPIhJHzMVZAgFD+XE/4sAEUn+mi3ZINUYkVk0HSBSn8+G9ozcq0REjOzMc1
fF6T07K7yPVZ9X9JcEpzwqnEQ6/6Vbb9JDCxGcc9m1M1qcVdlmQrKt+H9ca3ER3H3DLdiuCpwyEe
HTZ3V4ILNA+w+jWHpDu9sLOsB2mZiUlYc+PZKFQxP6Nx+mC78YKFPrDZiHDfgIXpW3taLYdHZ3Vd
CIHYZTVF1Az120bPvKPjABqry0T7hPOCuqP3oHNDTdGqkx9hOW4/N+8inr7byT2X9jRNJkMt/t13
BcKm9pCDukdcXb3N2lV53rkyNir5tOo0bKIlyPYWDOk9SRGKftVdrJl3tQaEYyEhvmb6N/lWZCXU
L7vCGX5bktemjDky8zM/XQIxJqRz+NqS6lkIFzo+l7Bh95T17YFCYtpJhKuTeLNPXlZlaZYlifQ2
p33h9Tx2CIdpiDMlnYNkPyZBZNCsb2ptVlaeVOe5YljGhB/6/6WHTkJEBckAD6dWpIGYwp7hcFFZ
xu8brLPll/ThfowxKG3T53a23rakIaFGfTy8kgmBGaJ8rvgGwmsIEmFBGZuQ1Pps7BzrotOUy5oJ
jHcmnxhfFAjzmU0ZJsN3MPpcRovC/Ggd9o5hNVub+pk5lzp/vQPMINFJikEF8sgv66AhHHKcKgcC
DlMKw/QfWpwvGl5sA0SZ1RZfpbez92xMhz1TEtTzww3d+L6kHI24eRR67efO95opJ3XuyLiVNmUM
C6i650WhqmSwS6gD1S6GHLkqECUO4KAnSeEd1M9gC4rzHccZdA8Le+RCy54xb/4HVWiRFHvFaHzG
KWo41ajhjPGCgfyvQmpLyZ44As/xU9kEQ6mr+XnvVS/h+ocCgbnnvWoTOJewR+iS8xVP/yINEO3X
Jp+7NgDrw8iimg0LPqcN2H+BGxN4CZOMT/4JiGAJeUtyYxM8zb5tLpdnQhYBhTWWsmuPF0+qsEHr
kXEvvcLy6l5NQMjZeuMDCvQIQJIOFn1NFk2YB/ohmiXcAwf72IvN83Pe7C+syuUfUjg+c582pyt+
AeuXYaOxWhN+7Cy1A3++Nxl4RfReU8nGD2+YCyEK/4UsxOMOdeNCCSItzDVgqj6FLYxL6q989ssh
4LBab9g9Zc7JgunAZbNtcPztSMT98vcFGyWiY7SHRzAvzvsPGkHKn8SBPSh2y8TlIzy2Bd2NYHyD
nNJQYcoXf1GXcDCpN0+2zB8Qo1QZ9ZbIt17iszE7Tym38RI+/A0/1gPLY/WcH2nrrkFZSoSbptVA
naxBHC2IGrNTem39MnJqG4jEs//KqF4+3XKbsA2ertW17nCryXWpGvbu3SigcCO41CiXG6dlnT3x
dvQjb+IHbAQ9ACV2YancW/RzewDwKOhKZ9p8wGYgQdw8ieUPAcsgBb1UXmkx+HCDWP3fLeMlkrsA
JvFnN4tsNcijb7zisYqT3CT7h53HGFGdnW7rlKvxG3uslvTjCq4+MY1CIttIfA6o+O9jEURv1hie
aMUEhEEkdm/q/dNSLtmHAzjiY/UCMvawXfEdtj9ezz1x2hVWwt5ss4qY12Gfi6w0Bb1Q3NOrwCec
BZrXjgJUm7XIWfkjU3DuTfZldFGxv+Zu3/tqd2WfugHxsMsZ/IgKtLLfFVLdaS9ZG3OgyIkSO4Cj
/Y0QWEjED90GxRxSqd8DmmkR07n3wVGWvLTEVCHmhbW3gbJnMkpnE0NEX9TFE5UpaFRHG5a+OcB7
PmlU51P9ZgTHPs1RvV5HSxG5GXI14hHBmhz2nW35x7p+fF9eqyfRTYAU1t+tX91ihnoZysM/zpPp
/H5AVtv/58JZcrDGZzIKjCXfvUpQLafEC3RXECQiD+q9UDQ9qtIO+CUQHaONJwgjTEKlBHZl9rA/
B9Auxk5HjViAVQzwhk5udMrdXsKMrdc6P8c2J2/T1U7nEQ3hL5ZD+XbaY6tmrp1X9Wa7t4GOmtGj
fjUpCDz1gKtSP0ug8IL7+hRMoKEW2o0VsdmoSDLsBlxEqmUL8YvkK3Iclyh7fKHt1d4qLMx53ouS
iBfYm9CLTDAuWVlNGQAT8I7wzz2xhGuSW05E6XfDpSwesEIf6atFvRxiiv06PnULThUn6Yxc2CDx
QEt5tc12riE66VZNhNMi5VmdQZZqloBOL5O5v3IK2HstWyKBTSf37Lx4aUnLpvjvh5Jrek93JTxQ
ezJCgrRuAa+6vRNNDgO6l/DxqKpCBIG9iToAPA2APfizjccoivKs9cCzqWZKyU9sfcHbWiBabk0+
yNloVsg7w8moeE7Q0X89zvEockzYgFwUMcrwHsJTwOhfRiwvr1faZGSZzmFXhgcS42nyuGlP++LO
LFQ3S7cbeHbvmVz4jFYle/sD1zdjT/b8yJUhY0UKyAvi3k0Ih7Yx4276ent3DKx5W7gUygG2eCJ8
Bv2ychYlBx8WnbjK79b+P/csqPi15PbyMchz8MjYDjG1gxErQtPQcRoTCCdmN2TGDbvOOUWxxf1K
heaL8PnMatlf741AaLsJbi7dPqzIi5c51eKIyyj5hr6nUi2K9fS5ehAf1u6mzX37AtLvC+rqkdlx
Cz578IYNYSANfYjErm/V55Ylr4HdbLYYc56crgJqgWVrlxbPGBTfjh+HlikM0YQnY+6jqVK/9omf
K0vNbN+r47c6jsmuhIJxg2ojWZVrecfpVP0ztRG+J3wxQCgsS8pWe/Kaa8BSgjNlkxw+mSG2n9yL
rRU9cjoy9CiJKHV5BQuEAgLCfztIRUcq3X97OW6kVornZDHTvsU+RKvUrd1CizXQycoe5ln/wfX1
TonEEU+dhXqfVrko/sAePXJzUxV2rlC5gxENtsMqUhPizh8be0v9yqRzXwIkxy5VS655b0+5oS6b
mDWyCtmaVB6zjjf6jDNfqNJLO4UL3k6io2WsxZtX4eOoZhDSBZ/sWf4qXIqqnpkSQ0oME+hbh0Bd
eONMBGEPszFpC3KPj+1gWBp7q/JTH+mwk0UbNNbZTHQFi8xEscTexFKIRoZ7DoJSj+35ESBdNkHK
kXeuJII1o8ztCkBc8j+Hs6VMk9UHNcifLuIUBhZEOfO9ZRiSWgPVwkSxJ3F/a+EuT/CG5zNVQMZt
4wcOoSucFA12KnjzzCDN+1+JJxq66vUK7WRVTHaPlDUN/mx0EJmXXhc9/+NcFvGcyYCoYlOGQB1K
1t9g4gqOiW5BBX1y8EB/Yib/c3B2q4y7Hufc1uKrDaRAETq0bAY7rVZvi4x1bco3CGg2bMRWQnNW
Ovcru+OJTw6mU8lAdVpZjP0Nn9iqaWrs64owvg3CGnSHugvrvY4eM+gxRBSbuESUKD7eaqIJLVEU
Fn6B5SdWTLsw4/hGIwYjkV3iujKG4I/qM6oqTLnPlnT+t0f5Zo1LbLxpGaM2D/e1NlupnJO3oUoU
C5brho5lepDWVIrHH4/DTS0rysu12vjsNeniMaxXCKTMgCdNpomAIm4tNU7dw05fsw9QDqMhJSzJ
WrFDBNuzMPsPikXcstyEN36dRcH4V/Ex1Lz2mhZLOO/698IQMBES8Xcqb9DTfIiG+KlMUqJbbuGg
mxMckjCASu9xaydlD57Eowfp1oGkFdGHW+VULCDmQDdd4XtlF4rvXz7NJSyH1ZUs7LqDeQ4ylcwm
jJmWX7aDmPq8gyXgNr5BkLwkntpctxS124O+HUFczAILWldFLKN3SDvBeyc3TIfqqqdftuVq4IqG
bLjRe+NKwMYwFJzI7l6w+pVW2CV2q4DDC1cIFJVSL8Irmk4FDnzVjNifJ70TB9yWq5mWYoyGba73
RUnJHOuYySnx7R63iToPAzscm07Z5FJAeQRZwK502zBCrzaMGC7xg6pbmGK6OLVKPiRgE9G9X+t/
6XLfYkf2p7L86aa0ZLce6k229VW3lKWeg62MLdvFA5Z+w+VQW8MyrGo2GsoTTB674JLIfBRcPvqZ
6sEhyvNU777Z3CIF4OFT64ySCGVPP6UEZVF0m8o5PN4P8wPU86VbNNcOapGGM7Hc0VSF8XOf5hT0
jnukV3s2c/yAvli+gfcq2NhSBSd9tTtMQBTQtsjzS4yA2DRU1BfqHXyxdnFuwNBrQHu1wsV8CXvO
X9FLosnaoXYUG1dAXjkwly541HxYokxmAmFzmjwcIUpK1bv7wP8QookVgauY/wwuYpjaNLKiEafp
2snBtCw8ZTvb170tspfcgH74ALH8yZFmHZ0eNBk5eQ5S0cV0cCI/G2TIs/GptduOKcer64NM/NRx
EIxR+RiEkTlPuMNNUherlrvnEfeyl+3zWs+nN5c2c3evSCE85HQC6Q5YBFyfE2MeU1+D6fAXKWvq
HXL0gadpkyQ4GTqP2ZvxHNSTl/yiEBGewiSNy3F2Q5Js6qRJQQK9+KHa3hxRXf8blfuUnQNTxHVg
Dp+/6MbyXbkK6ZeMc5ZrCRLzMzyhzJkqHmKrkSvRQr2+BNkkumiaHTJUodyCWDdrwITVz3m+DsC+
G1QJi/GmJFoygjaQzumU67CwF4hsbpLcCh+izUmC8QDjKwuJJhpmXQj2nINp3OUCkSBUe//FuTVT
lttJx00aXAjgX/hdZkFbR0tdyuUc1u65Yoz1U78clu/9VfCfxKfYkcrvL2i1JD8HWL1mm0GwC02n
aOhwPiLaqosEuPzIEx/G6c0/ddoW0hhmHX0PtZY2YgCF0RlnD/gs+/7C3zlFimxPkvkpgagKHXaO
mxiI6l4UcOW0Mqwp8w7H9RBmXHmWvwis3Qa64iKWN61ssgfwDypWM3U/xARXdKgYVj/E5+5inhF7
3fI5XhB8JbKL8VZZ7sbYv8LB1Ecx/DkWxB9fRL1yLeMjJjEWMiRjJ8jje3dHun9LU6Jq5mAJ+pkK
nUprMIwmAyEHX1iTSV3X401Z+A2kQqe+5NpMQchp+2r73ACDtT0WQEQWxBgzbF/rQ5rOYQTOczBu
dIS8FxjjD3F1/pg/9wgnGx5EOCbZoKCZOwxhdP3eikZImXgsZ0xu7IFYDsMwCK1OaYX5e9kXj7+v
pV1v6cKXx2eOs/AS1C0dju6pd8j/Tcxq25CAY9jQjpEou9ESwCyGln1Pcvmh21sj7yS3iquciuhl
FiRSFc+MFhAlN+rAEc0AQluA9ZWxHkFanwAW4lsPFN02h1OruMHMajJLe+DVAODzDEa6wmTBWn05
qVgP4VxTtTwwIlP9qNjP/TAKQpTHd2NC8z8f5SE0KWE6HwSRRbuvixo5hQYNsHp43AxZ2lLRfXZ3
8eCLlkCt7OGFLhKQj0qzOcjzK6sKPh6obLFsIJ7+wZ55v/dzWoECPuOUS28uOm5s4YXAkkZITnB/
zZpAqLxO/311lppeKnXVroRfs4Ok5w+6TSNw8Ng5kbDOHAm6XRTzG+oHXX4soOt2ARnIx8WTBeHt
BOzTuLuE5boqFoaFYLz9gu02Z3f0JljAl004micMBH3MEURR2bilKpD4TMOzY28j0hjXjyiLpdD+
dsevrH8TGJ6tSk8PxKUl9qkzmvUBwVzsTsj4eCurfCY1pV7w2hl8oRD+/y5VGkxCW9a+E5l2jBEI
7XLx/LBFwptwVgWICRCmdUHdVLP1eKBxG7AzqyAj52R7RDwkNbcPxSNtIjy00VS7FKux3ryYvFSE
aeuxQeNoYmBLmyLGYD2oDtMUiaR9W0U3DaxIUW6Qkmo0WVyWk8O/6idYhROpLoeq0I8pSd2bpsKY
JJy/BRbGBxGNHxrFLjs6TT2DE76CVUEG33G9R2FA5oKK8jzwavcYYtfsioKbjkZekomcE1gmztgs
5e+a0dX+71g4UUUPFHKGkHyV2Nx9VKJW42Kci31Hn6hujM75Orgcc1a3gix9otHN2SLAzusY+pAh
Ej8GQ/Z2lptIZH0LhGQRPzwi6JKiNXZ878o0xdNWLKcjRpH3MHjWYLIEYCJkSfJWi8QmuqlGXc/U
+5lZjPHq03AhYaXvm1Ip5+RYELUKwthl+0nhoAOBXKmnO8APidU9wDK4ZBLdzfqU3HWZWMvbPd4X
tvBfx4TVENfyj63/inJxKFIOM1rG1EnYSGxYID9oq/0e13ov4pn/3ZryktfEZtqwuTTJI3TEJcad
r7FalfropJJVFyDaNVReKArCySY56bPqJpGyOsbG1277T2fK3PuW2ZDiQgpO2cWkmi3Dz/kh4W5x
H8zCBw9sPjeGMOLHC06zgeNeeT1TufCY8bOQZl3IZiW9g/hAGl9kvwf0vDam0XV38qvmQQWEfxTC
fVXFi0MYznfNg/JO5nREUM1kRoS4Jm6qq4oJEoKOk6lH74kTdS9CGIfZvQc4jhBactgYuR0Ji2l2
DthB9xrc4ecy5rxyULSQ5U4w6GEyqubFNbUxC9HNR2+7JFqoF2bbZTcEShenhVgu5gr8NxSuAtTF
9G5He9mbGaai1AoVaPN2QNDkPP6/M7OQxArfQibvjxq1mUA9wWuIjA0cPxJADwkflkmSLHoySQ8F
sJJBMHOweFZKNME514gqA+0+ExLtJBJWLL4+nJC1fyaB1Lu8we0t7jjhZ1+LJbImyssc7nNAZRKI
b0t8iPz660tOTtK2ZOvkPtUGsdTVenTQ8/hDwZQtLcF584QvlQzl6kmeoLS/aJD87mOQ2NZl7jDx
4vdUI8/xnhlMJPOWHqHz83DLSMlZsD6foh7UXD4eOTa3Sd5GvoqG1h2JHPvTVcjPE8OIFIYC6DL6
KzpcxJ6Ghk4Z5oDiLWpFibVY2OJ7PWzv2g/wy1jHrCHNgCUpH2SnnjPRiP1F7y7E3LyAmW+e37KI
EIcYYhBzb6ioMY4KfXjX2kmY2nmwzf9dW5e3Z4S1gpWajaO8bBxy3by4bMfV17IQQRJisNaPQKGE
F6IsPKsf5WQ4dDamCJGI0EcA7fZ1QQRxHlOUrLLm9M9van2NfnOUJOv6ikX3WQWRiq5k5JqrIB/0
/KE0V6i75SZni/Clc3eSsEC4hEKskpB+6YbDxfAmswhss0xSj5Rr3qEj8XDUa1o5XAhT5OaTS0Ht
Bn8hN9TJrbiNPiXlusR+eaNJfzHDh5bYB+FcI5v6tqzsMrH2iRIkHCqH7Ks/hROYBOj/AAIrylg2
Oluo71sBNjkp68S4l+O6qPu0G/FRWTYo8wj0LYZQcIFMDjJ2pOuupBc90pzzNunyvNOmaHQra/3n
ClPUATs7fv4zLM7v+Ywnb4L3faZfqtPbP9+ru8v8XOtd/YB9IolEP0Kofesa47jcPyBNsQ7Lyiz5
zMj2qfnomxX6dW3U+ev2YHaJ/oUGy6OZQ1cNgt2FDjxF6TIg4n08k/rGtmfjpKT8h2CTf39UhX3L
szA0RhibDItWvKuEqdz5KYDJwI8sclfKJSZ2inOKnQzuH8D5yyHRb3OrAR3vOyOfdYmkk5DRtchd
+sYpWdaeDQymKbL0aBH1DT/bXiZt/Fv6asv7QKd1QkFqoFuyWScb6GXgAidf4WXxfYuKaagilZWZ
RtWMSGVr7UVHg546voCZ0rRPuopD0Jq8/P8/IEBzWJmTaDdOHAMeRF6zoN8Y3XrMK/JAqgeC28wr
ssE1ep363h7UGVu7VjxMUljvNcMJNp5VlcxXQrKcalN2M0kHbwxmmZpOQQgc0m5NA03UcHaLQyfT
VZTb45/loIv03/PU8ZGNyao7ksoEja6MNlfXu+3jNoF+84keHFIrfY2mBYxCbHD99nh1qySItuRa
7pUyiQXnAULlJzdA3cSN/HSrkt2YoDyDDjXAvwhBFFJU4R56VSj9i66WM36afYKWz31p/GwA2IhP
+/SBF8InXyAjqcJmOQZ7hdyye6yXQZa15tQJkIMORNT7g9HVhT3M82XXcl7p+BrRyCEUY4WmBPi3
soKinyBHERd6iOK4r3BTZYUXkNOCNd0Z1Nz2TNkhDByUxRDRpG3qwYlgw6jxsnPVMR05EEY0KZvi
eU/51ntcmOQRzVao3Y2lsRADoPo9nMkG/j9RT0Me58MvpymV8Mnp5qlNPjIL8ZNy/xwkyFAkWFGU
e0liH1/I2wlpgffAQbde0WwS7k+j5e8DRyhL3FxCL1RHumbdQZJlP+5Iq85RsQx4juAIssDAVt5p
w0rVBQkjhEJxbyhh0Nx3CvOELk/b5A1bKgCxd6zYZH+cznrklvF5QzCqYn2s2T4C3CGpuIS/u2PC
0OHhQQqg8B0T/2DrFfLw6gOKl6Rvade1lcmetIDZSEyXRThNs6ESB918qSQRBka3HQqStUrIstqP
0Q+gT9jRBvA3/MkJJDmd2zWFfjVTR0QCniSafqFBovZ47ZsS6NXcVY9NrEAqPY85IoPcsdrbD8V8
rwm+lrVvmfgnVPdimaHbGhbl69jJoA0tXSeVY05PEtuGwfvQYjy3zwnNXt51UNAkyJIIPsoHCemq
Ran2lWmP2muFP41uXJyYwZg4SfZxFNmeOCXl3QT9S3NsooEuYXalfJ4xJwvciKlmoaxfP2/0bK8O
nkuGhfkmUwPr76f037T+I/6plgcnHR0g//iyTJ/WUAhYT8LD7m8iVU/ZKva5tGLy+Xx9TyArKlq4
j8qf7Ug6FkVvmfdf4jjRyi15qWegwT9J6tW2hXXGsTm9m6v3lJKiaR1fokCDROUIM+Z2Dni+mO52
dGNj0QcSycbaVUZG89AxqYhNo3lG7XxS7VKmvXjiulbTsbUnQEVoApoELjEVEK28ZuAkrfXXSX8s
Kb99tGatm9foKeEup2r82Hj0e7A1RO3qB+JIq2E1fOSGj4y4Sux2pXxEDTHjPboRzN9Sch1UPBMf
bqZRYaLLjevRvCsw81Rbb96zxzwc+9B2rlu38BNSmilroa0/7O/nfAgDqlmb2VACRrCET2KRbB7x
re/ab7eODWf31tozZ8IyN8UqmmLGPQQfLuSFvO6XdaeHU9olT7hIxAsgHZ5tHcDj6Nli2I2hNdb9
7ZlPko2Ef3JAzj3bnPG5o3Xf75+lPvm+RuEbR99NolfYBEirihvGuX+wVN4cfpdbsvOYOX2d3eVs
C4kSy8d6YbB2H901R1pFAZKvgwlLds5Zbe0M5lob9fIZJhq3f7HHaIOJueL3W7A0+BUUdC2nTdwa
GG/t7PTl0lteVfgdWFzsDR+f/mN4JRMXwhd70ilMDCyOCS/mtR6bDtVm0c79NPvMXSySCfuEFIO/
TTdbRYDEGRfInf0dtZKArlpnGUYjNgdUxXeyJjSG7Ax1zTXvoDMe/WXWy5oC60E6LI6gtuL1cfTw
rrwZRObei5xB9gdLlh3612Lm/riIprOSTYTwBX1BfXDqb6HtxRNUOljyuDrsdgHPOi2RGOE7hDTE
BVv/GJhmCIXDGLRcxFayLg4vYKJ+02sZVLjnKTdR3IeEh4oqsJomLvPqLYD8zR3uTs9DRr6BlE4J
T4UuravhJQn2IGbfGHffdkuyNySwBIJUJWpZMKa+6DsfHQ6qYwxnwOy5ZD4AhsYgU1xsLsBWJfFc
zNFIwskT+xAA0SShlci0tEkthWKjLg7nbBBfYOwMPARMVqD1hVvh/Xl/+GGw62jaCBjyfkaUw2jY
/tpGw/Gefs5xozFIi2GrH50EwQLgsIjJgfK2xsHuAwFipHpzI7zVIibWLCFi04XTDTdGYjAbvLmz
G6NYvbK28pnXEhXQDIe2WUJJKV27Ilep/ZhHvCmJeAdEsnp/phExOH2jPyUL3Lpjod0al51U4EGs
abYmg0hdDK2eMGEjc/9OLrOOG5Sb+byZ54BjMFXRXCcJG/AhfPdf7ASLIR7OX4sAplV3iwG+yF3I
vww5lmynckI6qt+ElT47mlPsxpd4sotA74giaSsFnhEA4HNb4C9mleqcuRYrUshuGqov+DF6WO15
isIXrP6ZfyAOZr1HfH5gAJGcIIq/muDuhYbxjFc7CqfE9XONm8YBY3UKIc9KYZPWqH3qxp20xkVr
F3eBCHTgJSjEX7XRflT0Ig5XUhmKV9PdIouo2AX+hk0geZy5AuNwkIgQ2iHWWG6/97CUdb48OBgi
f/65VhsFYRIIzZYf8dOBiMVfB1St5pF3tfPXUyhjjJxBkv6jaVnGDxML6cfqYlfkU/zQK/6zrsZU
Yye/sQCJnR20F1ckmYEy88vW8HHK+EiFoJR/ggcpmv3Kb127E/nH6Tc7sz2FqzATwzK00AdlJ3eY
AMu+FvyFLP1fwK7TKcns3SsP3O2ZIeaLNpiaZ8PQzvQ1s2C452CDwYAjIMX3mcbAAPmus/7QDE4n
MjAChAB8lacuykdM9gFEfQ2IYu3D9W4Ce2m+advGLGplMNR5WEaOJ50wLC+8EI/xbvMGSbDyZk7r
50C12AolHS3XRtBFvL2PV18GznUDtgO7tOhjhPOVkxd+9TYGm4Ku6vtHT9Wie8rT/XLx00Zl9jtL
5htxMv6FmJsch1UOY2Pbfq21RgksMJB+8elJChHizUh2D9XWWLr2jNwFa2MCMVeC6SlhiljdoQ8H
JLuYrriBUGULVnSQQ2JsQJ5qHh9FToy/Q5hvQiKTG3QRhK0RC0Bp/lxCIlDkBD1KVy/+ijk4CUb+
Sr+siOkX61pToqzQU/vz7HmO875FmzseZl6Qou1rdUnVPuqfaVubqJOa/CzI14/emuQiM1H4OHVg
X9G5Db1IZOcO+iiv0HVgOz808OnbiC4e/eWFNUIw2B5pPbVeVb45rEwDTK9F90usfGGjdGRLZEvU
lpepetz0EDEF9zsTh1VNT+dG0kqtlGAOjo8n4rhyqkkfVzFBbFlwO2wuF2KouS9rzygkTED0VO1g
A5XHmVtYR79zag2cHxBN4p9TEDHOiLLPUhiXQZm2LVS4WcRrFLteO6eP+lHyyBdiPnLCk8oYxh11
ZWkZss4agtVUy74r7aS5mUbHk62V90pmkQ7si1Kd5ZB0SMTSYQWJEWyVvwPRoCjgQlpe3RmOhXDy
4GRa7mkB4dofTp66aGUh7GsJXNWFtFfI2a061iTmYYJ436jm5C6WZfYMHAAai41ZOORzuwDm+nW6
hmL6bJc0Rd4qhTGd5KIuIZhi2TQF1b2VTgfd3Y1PgBBfBxCVawvq9NCI/pDPExS38b2ow03lREHw
FfLXUgc2SHRDoMB9StqBaH9XQIgWixn21mTeJLP24uKwfffvEkMZMAyIPpsuRMpjuoH/c+vpTjzm
FAdUH68kwvTXAnYjRm0lKeF1lDkkRBYfzHXRJrTe6tNbgjYe9kTctzQuQXV0Sq1LuoNatlVefaUS
pTXfyubjK/dutQAT0ibE7t8TO26lYqtLA8H0OCZRrOOOz2NC+32/hKVjNtknVF5UYqO2QpTbW5Bw
yeXhsS0/nxmgd5RTnl6zzk5vGrTLig5zWYFwa83dHJoBvWeyLREmfRMVfatFxNxquaZWY1TeTtsU
FJygDyTAJZvRef+sLH82D+Q7E0r00ILP+fD8zvDtn0umCLqanra6RskEVc+ELnn0FzUtxiVP2wzz
kai6UuD03GYYZVXP0gpDKphgB5PMkczcq6WUZEtLszvpbNY2lnF356Vk/jxFuSMq3LensR9jiMz9
N4KV8KFwlFu4PIb7K3hUy+InU78zFvMhPj5MeWRmtYkzwD34znxRkNAsMi+g9Acl9Mqkg/PlTAFY
mBENPemJ41qr75jNEy1yddREpz7HTY/9KRDNqqnfEBaWu32UsmFFxbLUiGSncKzf325JtevxVfP5
srRyKUvI6Gwe29EqUDEydIsSfNF4sQvuwxo+osJjvRdXOa4MgX9ONUdXiR3fyww0wGGaCpYnN3MR
S91y6aBlbpaHc2fB03U9IyuIxW04xGLJkx7J8bb8+dv3G+TO6gXUM7hfZltv6z92mwugPinHynZi
I9pMmqzRZQ8neAau9LvOjbZlai1YXPdyMALilCSEtbhIRuVlA8xrmrZ0W/0Jc2OUrz02IIdSL2kl
tr+nj9tKc+ElZWsAAR4XqoXvdTJd9nsIPBdauCTvqjYki5WlttiFJeN6raIa12sC2WTUX6nuHC8P
dJ+uPFqv7wWzhcukwgMlIBl+VOEDw5NhvZ57HhJp4YBA87ICNUB754KWLEHCmgRg5miQ4VARRRkN
NZbgfT2CmQ9WrvQMX4Y1DHr6aHZQARcI6E/RGnA7VsQdBSFHKBrf6mGRl9d8PINVhcHNPgG7vfnb
E3afyEr4h70I/3s/YfLuIiNJnkE4nbG8ii/bsow6f+Y08anpODezDDYm6uTWlK47wQhC4ZvNxtT+
R2eLWAjRzifvuhRLg06md5MZ/WWnH8G8UPYyff0zOLwuVArXwfHohH4jc9XLdnoA/SSVy+zKDUpH
ixHHiFdH+QYiTZQ0JoLIPcAkT7TlNKFy3A8/lLEDDEaazPMs4R4DsW1oYiKU1AD5jd9DC3oNI2rs
Bk30oc7biBZsyDYIAcX+IFQXGhkmKU9N5prTbjNddkFxy5AyE4z5I/oU7CDmb2qcGh+drJRrrhwN
0fT/9gPCBffvdOk0YtEgpEFriNy7yyW3MWk+jLNCVYIIkNnfM5GP9OBpaZ6qVczEBKN/183t8VuX
KAZH1qBK2EFuPD9/XRl0+rNqm07M7Ot5HPA2+39sshevm/MGAZa4t0LeBovpPIzc1dr2GmXq9597
TbyWZOPXhDjX68bSKBQF5RtmWzc+ZNYq1+xxs1eKH8f0JlS8YfgWWEfoOFZ8DQOA3sr62NxqhMAO
Taae5q4M3CtDjk24FJnpES66Ydo0Q4wkT81yc0eV62dawepLIcLTQV7A8xrBqrJYQIg5Tb3hau2M
JZump0m8owZ11YPHWWci44ZKeFrO6yd4LPaFIESt4VYIb1aqoS1GiN2WEqkHTufmefttMTTqj/jV
YqOI30Y2LKbo3bOFmHWFWTtBhh2oXXEqyGCRlzKKKEP7TIAGyJ31skkeCPw4tq+DrBwUS2ixcuLI
sP3GY4kecWbm0HqSr6XVGhiaRx1GpM5sRbIUyfPxtD1hgZUFuu1tX8g0Safn8W92oN+FzVD55oQZ
U5ku45hRW6a4U1vaaueKLNVpVepycxz/7X/aIj86c5lEXOnlzr517HVrPtg2stFWMgpcBjTXrh3d
/s1BCv6WXHA/kAAldPD8WsGTP6NxLOYoeyFQcziWAPzXCFjwDQYKxml69zcBnKWn78i6u32Hwvbz
NUphO+ndwVS7Iz4xaGzWTBTYYSZvBVFbeVaq2wi6cs2wANiJF/kYKas0JBFw9Jk9tR0EYFl20jQL
gF3gDd4Sfx0YzrJ5zaeYzV1Ukg/Gss7q+L4eoS0Vxo31NQDEnx0cfrU5Oy5F1lLudHzzJSLtIBob
NAISF/n/XzyS2Fl11pWrKCthikhHqPcVYZwe2P2BJsGemfS7iyysmOcOlR9V6EcR0GiTc2zhJjzM
ZpEKb5fCwD5V7D0xmuSOzN552+xM51n4ErUoUDmKE6jVMI7TuJoV5a7IlEI+AbLgFVW+aeAcj6Us
Kd1uPK6SkK5mKVflAPvk7kQK0r3tv0aXDy+Q7OmPDtbnSCLg8NavLAwA6V+UsRkTq6CgeQElzqbR
nA8S70x7ex0v0A5yCiH12P1tYpcKYAZYzqDJ0bUKYN9UyCIn9CMKrRXazKf6yPQXBCkqC4sP/DBN
4SfxSZlj+NdV7N1u9WArUodHFi+l9vkZ2BoM9KoPEAv5/yJsD8GIIM1I5pJu3Shvg89hN4xC3k50
pMsb8AZhfCtYISnHzVVa+M7T9XQx+DnAcn8pyWohsn1dtccF2fWU91vDm8C9dO4wCbRgif891KDV
j3x9pV1cnvMyDSmZRJv80cWNBjAvI2Wa9ckXsTLBclPRcc91Qlxu6NgJxEjc6z8f6gnNYhMlgOvq
VrpYGoPQNa2MjKltm5NXRcsPshQFycbuElm+HwRy+BNUku5Uknx/ASn3r17MSWfNW5n5viI+Do9v
LgyZ802g32R99b/PeCroj80kme3FLi3SYVHfhxPcSMaf2NKA2nU3yO+tXnGkj0ebBAqszOyBJo5v
W3A6nc9C1HERIT6Xxn8pE+HwUr7UlHEK89rX7qFosOIbvtGHUhBhhFZtjhljJZS+FwRQpLPy08ip
nrD3abTzETFiMYZ6A76TujCq/TxTLgS4nXBK7TT3cZ2Aeqb3S9gDlcfYT7kjZ39LLByyX6nMaVi5
7Hc8lvbKr4ecI6UI9I4uOmr0qZEUsmd+OulKS2WDUvLHTGITLjixQ3Rc+zQeRDgv0n/KW1nyz3F+
0sh6+9qMLQgo+7u0y2rqCHES4jyTsJwy+OSM50GForTWViyRoO3zKqIcbYt+YILXsnvOBabZVAkB
8EsL5hnUdaK4XpEMk73F/8O8rVGgTfWoM87yzvGwOBYMJOuBqwGlphzxoQ3e9HEl9f/aA+m00EdK
DjD3+3Z6VgOuHydqze6SNo8Egg+9C/SSe+XemeAMNEn+Ne1GH993IbPceVD+9wjFdNMqsAr3ACmi
5FPkuL12A8oQkGvAR6XVSrRzzLrPtQWsfsRBg4RUXmoW7iO6F/CUqrtX0YEGMtlZxaBXes0uJVlf
29MU8/f0v5GolSKe9OESd+OKbrbQxsOp4xFWqkFLdwWyjgGxekBXYNmia4bl7HjaLi1w0VrcCeR8
X1Y69Yz3ZaEecHkGXMDNzMge72raVMFPWkxX3IzPBCHRZqE6K3luemkIjg4iB8vrsHWqWAuxFJU8
/Av6uha03ai+J46ZkmfoRJBEhM8P9pW2LZk72vgoFPbekyceNKc2ZqRm5HVA/CEiTx+opxditu6D
/RSuQQFxLrL5tkVQsV/TAI8B66uXhv8zmaa65cy2oO57ruuxfC6pBtFf78z9wxSR9VOyQkgPXM1g
JoN8Zzhocbhxpdj6t2UN1SPhuMptsP7d8hdzA6UZLUV9+W2gBiTIKZsw5k7jrK/9hlAcUJKoVnTJ
IGBVuZFnmm2jHZ2aYf/ohI1EKeH9DFrsEIJsd6XYN46mN/jLsIEkAIBebOcpDyOa3uraOAGsJB4L
QNQUTv92RvUG0GvMZRhZrcml3tGV0iOxLUP2+jpVPhdgm/qSDIFj/7CZ3KERP3bSX1p4mQmlvWv5
Q38PvEGWCm3rBHCTLpNiHs0PTDb9VIEGsBxrsvi5sdvIcycCt5HSlJoFrVhpN16DbTbmYYp6ZBv+
QBTEL7Gd7Lej/299GOPDBq00lLFHS2TYskoJjBtmvGNceIBwM4z0i1curJy6bt12SIIMMvR2o/hL
Q8cIz+elPEWfq9Un5X03Qnl5QM9NJTpd41lCMDdamCn6I4lFp8QZ+tkHC0cLcbt4boBM+nR22vlc
4Qmy+pamI31dP3/SDgqErDN13zK2ay+L/fICEsMmYHJPgkK0btRxXLtFi6SYCulJN7tbKLpWAKxB
x/iw83oVbAAltv3a26aqYRybt/RjydbYxgvWDpn/1rKtC5rrEIvM12pTx/rtjPE8ckdY9un/yhAU
ekE7YAicfUJClIT8GDtBCXT8aoKW7MzHB7y3vu6Tb8LIBCKKE0DsdAxskoo9qAW8em2tkIxDuxB9
hlbg0+2MLhl4oDqKcKlQUd+6N6GSrKAXSAmCIjtDPHXrrOV5bVCacXalVslWoEeiNnGnXshsEW9r
KSndfgKT9HBXtnTTM9yz/iR6dYdfmjzgY8NChVpkIzH9o+9py/W83SL2Wq4ITonqwwQKKpCXeWdb
rwwUVwfQ3bfATdJPHbuFnyT8nzPo6U7i2Fma4N6643fE9ZfuHxhUmCJVi+IaE/AY/ng1tB6zbSbA
h+dTnv1rq2F6GM823zztRpzZK1P4dr8SZCiWkUlWYesyMnpwAf5dYtH3yvkLoFmjf+RD3XF8RGjy
OcUm0hOFz1j54s519S6Ss9QaGmsw4KkdFC5D7pzGyKtymXSle6t5o5UHUxYbCR0M3gEPntz2S6iB
6qM2bBcJL4ywhBFQ6QcjGPf5erRa4zJtVUiM88J4Buqr4sUa0pv4dVAVwratZ6jHR47MSQXvZpYg
BWZfMU5m/mv+Qc2ba5gduUXXICN5EpVK4mrn4v4WTQsbnJ0WjA7AWhcpEFR1PyPptAhFotO8usxP
Dmj89vCoZL4uvzDWecYCtv3YfTiDsc4OsiXh3OQDPdXKy74Dk05Sf5fR2tXSBKPTN5o7YSsLp/2l
hmkno2Fk+0G3f8LvMfT9CyAjQ7SjjdjIIm2OYpa7MyO/rL1jzgt6XtjZBRSY2qwuhNbakjSWFUIY
M8fqP/aPadVKQkXaPHy8nDzphMf/dveei958QY9xYFlVCw40ZmS/yH4nrNKevIxpmK+nvbmKq7Yd
GRSP5Ji5P8pBalLR/MDQu+TETly1YXEjWZEHUPq6hH4haUQNKCHwgFTIIGOndd4cxgaFLNdnDMok
00PeElcgjxnlnvcJKSILbrKmCl2SSWnRYG+DG30AVaJtPjXFnw3iv9CdL2n/fhiezM/tlfWtOraL
i5OnnEdNMtkPbNckSaXWkIcLq6WNiP0wlg/qyCB4dIhjF132r/5VWIRUPlEEi3pjh/9Tmgm2hLE8
YVfpFHsSrr2CDFjdwKp27RvN1K3XGMC0uXNsfvmFbLTZbo9bjdEv9yMxKd09TZBGK+kL5wAqVrnl
B5V7fcgirgHpjVqI3W5HwHEcRS9q6IZkyT0HOwLe741bZS6T0CB0lKtdHWG4l1kqrT+NCYuU8PL6
lneIpeqcYxpkADiRWxCGT6G77m/sQeaWjGkRMEpj+9NCM8n7Gk72Zsb3ci93QI3mCkPVk18SBxH8
+oplcIJxFTCOKqL5Vm1juvUrTJzy9qFKyrmfGOdd0sfTsL5kqBqOc4t1bnlvFjjmvtH3R1GR9Uv8
yppMy5dlxI8R+yIPdtjRX3J78gJ/w/ATCVSDxilroxwai42Aqc97WIZFJjt90Evb73rrY0CUDVbw
L1+KP4JRJ7N/vCvqd4zvTVBrD76LHhO4oaMkWdSNtNozfoDhqdEMQqCqQVgTNwkANYEa2ELpUdSG
2/lRvP5p+wFm20Z5PB8Wx5tyYBMIpYQXPnvME9+vlGnoi0DuvcgoMDEhP9akkdPeb1kaRk9phfUb
+kLSeU7bETKxfLkQiWt9stG4+trqW5r0TwxMiXrmcmuFToFp/YfE9SxtaUigBjzHkbSx9C3NnaqD
X5zR56OIWOImBXzqQks70aKQja+j59yYR0cxdNC9pEiioOBRtSFaNvtHGwscvrAkYxuf5amchbsI
eU3F7JfGiYqyq2kKfhxufGVwy3tgdMA7kalLXYmdow8obu06guGXk2WywvGAf724lOMrogLDaJ8S
cCq7p5vXN5hQifBeRONU1i1JF2WChEDdPtFoCcw5Ct3hAuKGvu1/u4+LA5VfcS0jG6pEMHFvk4H0
kHbpCBFWVzcd0kruwjU11m+nJC52okMaZRJAnkqIJXFRtPgqIzcf9qvObMF8fkDMNEib4GW8bbpq
f2xuPDx3+owpwBT5hcboXQw3ecdKVTmqiROJtaRu2X/+OzEf+UqFxe0Ho/cdr/HnRyW1LZzKWrnw
4nvYeaVb3VCDNkdt3EZnR2NcZl+RMn59yvroQtKWUEg98BI65a7Sk73/eFXa1SXyMbNzdAW269Ll
3OpC3eNsKGTjDQmcfaPzpJ3oUK28/0KY1X1wqqtG6LiYCBauYpNvArqX+OWkFt7YZqTe6+/xjx71
T6MM7K9og0pX4pLUPWnxcETVCF8E5epS/ZmtncW23dsNJt30UWHbPCldicwsdc+gi4eGc6e0p5vd
ZXh2y4Y/xAIMFt5uvRduCqrVJJV3ghPQ2Wufurci86uv9Rw4BcSrU9TNaygUxV2iTQZHT3EfCAqc
IUtTfmLs0+kAptd/yGJ1pljWuje4CL8q6Jz37UF0HBfmQaqD69ew4xrztDMyoBHDZk1kDsT80k1M
oYIfMxQT/+3tCDSFuHS01LFIeXihdWoFGErHvcHwnSTSiPutQVrRZeANjAaDBXUaPUt4e+n7fg9S
vhoq0p2d6jMQNOY0hshKPAgrK5TjoUIPp8mfF51i3qKptC2X9YdZRlzk/+i5qk6HzHYzjGOY/wqr
Z6QUhHQFSshjHQjxf8x6rwEezb3OgmQ+5/jcsLsPaV4hZkjnFYjequuq64CNtWoghDvoGaqL7PMD
FVoNGikrhTWCxhM9wyPDemc+3OHTTJ+mmpa3FF37lzRNrtuNGkg0x55zpsA8A6yVNeOZhmOdFMWS
Mh/0suOUPE73fATdRADz9jtlYUkidztZRdW2n85eMmo30wcs1kP6kyaXs0oogZYMGlMKEnPMmXxh
1297XaY3/K2cPvvGfdWkY1xJVWHHJyPzbz7QC/+NVMOXXtn6RG4hBSbFfXygU1c6pIkTo3KOCF+w
ex3kYOqSRu6htdyuXNEQEYNgGBAgFYB9RxcnE/AIJXKXoC2KhJ0Lk9Bs5SPPx1Ee5eC/rOPdo6Dn
yMEh4etb53iYBlBtwZ8tPCO2wOMoU4uRKa3CgK6QYW1vjr2msgQSHv6WHZDGgNt2D1NhePsbZ37R
CX/l65oyVsHaT4hx3Ib1j8I/LwJ6Ebao3GrQj+IfAmLLTKB2/6a/7vHMo23QHnXQmoTTleSKxkz3
x7dg4wpZh8PsjrApgsWFaH6gtdvQ+GCgY1lAINIBWUfOczgSZ/ypNTi7j8aAQg9w4B9LofGRP5mI
G9rgHWGBRdY0fvnKGipPrpR5RKW2V5CdBFiAs+raJCOvH1SbjylPtqm27/CZmzbEr0JCXQqewOa8
BpbxEP02AAMSO75mQE8JzS1vqZjX2/XCM4u4ViPefutyY/2BvsMUd1TKUtnopwD/pEfVAfz/Q+pt
H9ReyYFuYbJJCMqcWraN38bh5xLhs0mLxZNk6rkG11DFZAVmtNda1GOYwuVzQjlt0nhc1wtDjSvm
GUygnPyeHd/o3fF/FPsugW9Okp3+PJ+n4EXkfUb6VCvK57UTP0+C3czr06T9v+IOf75iM0qUCc8c
WYYW1i51e0UzIH+TP6PXExEgdbhu6tgMJbnBhA4TPBORzb2RzFL+dQwRdaoZjSdGvRSoe1fVcctq
N7DjgeTytA5SzECm7wdQhBscqOt95iOLLJIWU/0RMEJkmOOdCnPtS57BCaqHOrsbFBbjm52K9oyr
QlcrV0AMn2AsNucSEOvqMxBRl59iJ+hWTpXiR0Mha2oWq3ZiLCFyCE7ab6KV/RgbO9Gos8KK3As5
jz15t7W09WJzKnb4vnaQHmjowGKAgsPYkcNO5FUuUPRTzcUSjK1q+7HgCq2c1TUji1xVceoZLY39
/REQnb2CKW2NzPFm+4Jrfn56tECkjYZ2yutp76w+hZ4FU9oqe5+JnOB9hrQ/pZQBVp5rwreFgA71
jLZHICOjSFfs/JHEnVGEwc7IjxzujqF+HWwb5LFsvhPpii9/B0tG/vCC8kYTcCpwpf/k6iHF+goK
aKemZKRGnAcwdUEsFNsjCegdOPGWBLL8cvV9ZC+jsyOfbkHhlBHxv2pIBFoVihh0XNmhyLT4JLwK
AFmZ/zl5ov+p60EWrxDS0jBfb+bTnC2OTMWw0/B/2gsO1S2tW9kqzovRl2o7/Xdx9UuXfmHQ0UAy
dsLEnp44tZ/UFEnbRzQWlU8GTBwGHzVmpmOr0JjWEsj3AYASU3gAi1srZnKAgOlOMr5z56nQWnDp
7Y0wSa/GczDLtReQvKqMmzsdyrVlwSynzwKIMnAxgL2WmHIKO3S8+n1k8R3fHIxn91IlezfZ42BB
an+3d2DJ5KcPD07Kc9pvRDds3SG9Oy8taLFwWhMMoYexxACgFZGFodzGDhA+kZmpvpYQsEg5W+ub
89j9fgd0EPf3lfLmOIHXNrCxgXlw2daIMw7Ib3RCNldcPBdS5NZqnnJSnN2ZxIHRJ0MWn7E2bSBK
WApkaXHud0c6hwno+WeC5sip/nFkRg79Wb6/lALEN0MTGKHdeWSigMFtRMz2eY2T9XSvjpJlNMcR
OiK0I9YoPCHK99LH21wO1uW8lfrYZI2WIaMGkQRqlfiRYruhJxXhb02yMrM05INqGzKc3OgEMLHa
G5l/1Aw+2d5mWacNDb+x+evl5Cxt0fRG/XY3HyEZHhHwLpqakwdk/giJ8dhailbVD6RZUrV17Y6h
+5dud/HgiipTGWscvmii0PJebUI2G+1z0sAEB32uxywQTjgq6+MaR3ez06wQR+4BzudmW7V1O3+5
i4GovvTi0/jf32oI3haTRaofmnjyuJ46ncRQLGAPekGYpdF0xj28IzlHKF3H7EANOG+MGBJRmM2/
SKEUF4wslC5gYfa2zJ+eJDHSYuUCTY4QxEFgXCNfdEyGZhg9AweNaJLKagDprXrVqJdc4vgNKO7o
cQsjyHLOfx3ck39pkNS0StUUgXmQ4nzSNfZfLaHLafc3ZnTxLnoRDtRehaQQRuBEsS/m/RlPPP4e
LSxWe1JC4vUIskllOD96R4TkdvZ0w5SmSFtBEXizv+C6seSGQsoH/uZQwqb+zNt0wqkZRlzVm1/X
n4xrFNDDRrIDL4az+qzlWS1adewjUdYo1Lt7TPztyMNaAaHMjJXN7pILOMTGOP8+IhUv5652xqf2
sBQwQRc/W278Gp6Q0knp6D9PcRrzxyKZ8QArut+ztRWFXr/y/IolLiRknm6UvQBDZJmf48JpbMAo
K699z4l1KHZR6Dtne0bBjVWlMHMza6LHa5H52uvd02+jZcGpwCUX/Gp0cPDxvUiKOwOXkJp5mrj6
Ksc4KLqT4Uc0zHQ4+JBRSmWJRZsv/niCsL0qMMzbHXIs1wwMeBOD53wOuP+O/Pr3ja7Q6dOeCZfg
bDf8/u/l1SUiceOEo0qTrA8GP3OjY5QDlQU5wVujOAOC9q5E23UzFRdWXW7Nn5bKvjRuHLHsqyZH
kcCnkxBCf7GUMp/ZexPx03UQVqmxAqylm1tfeWDHCkLfbPIG0bPvkwcp6Q1Knf06q0oYrSSdIPy3
c+0aJHQ8Fcrmxinkb9s/VPfYdauPkTE1vYkVAV0A5DeGYf+MGzrHib9zvmln4DIMot8yggqOzKDY
9p6FtfC88MU9hipvwaFcrgzexK30nEnWW2chf4k0GpwZN4n3Spci5XZkIceYmD6fgbI8n5fG8Zys
tT3Mp/Am1Mo7iKAIKd2jJtYG/+shiSOjlcnlMcPBZK+90d08Ox+GDr5nLZbu50E56JsdyOgWX9Tl
zh1rcrUaV6OYNWPXMbaOQX+LgYQp6IvoEi7nkTGHmXf7nCM5acYmd63U7Undk9rHxpTeqDzkJczx
Q9T8cDNeAjRAF7d1amehdx4zG+O8dSfO3YH13K87FXVggJPbBeqo2RkjDHb5b0lNJIsfL8P1xf+0
y4SSWkIO647D1Fy07XSrzDHaTAdsxQjCQKHO+ipJm7oaiIoYxLDATBUiMQlgkbQtFXeu4H0/Qvxf
N8yGrS43SnHmXkknGyvz9eAkWGHuE4XtSapETrm5ON6e5V5qXog9Z12hzR5hj6zE41t8Nfqgl2Ig
30tTeqCn+TzagnCYIEDXYKjUKQO2JqWH+nSwKUuVziw7dJSX3YVrmxxW9UYQ+jOawRelFqmu4S9J
k/XQOO69aFE/J9lDpWUGe5xNZTs7WPxEmw2kzSUbgtnea7L711DP9qif5TkV5AsU/0cKolB6R8Wh
H/gdwR2TkZ2VN75t39pjJ9rkTcC3PEvISHW6WwYCXAcS7QMdAp2ubKaKUffp/om3+brEpK5qeP7n
NO5ppv4q88ilvevYJyLYXJrnYq7Pedx9We3O8rBmF6C/McoKHGPCfJmXeItrLv2sr5sMPmXZkpRG
5V9pGfyiNddXjo30N5HHhMytH3H68QlYsbkT0Fqjlpu6ytLM8qLYeE/CIYRyLDblDT7ON2UtE4SW
BLtIubjkOFLEO0h8+wCNdVaCA7apkzRRe75etWquKImAeDbpkerennNReyqJ0DyOW//ELJ50VQZz
6mCJy2lKEX1C60KVAuiW5+9ZmgbnCTuN+B97v5yygsXDR3jc7OJUJlD9O6AlaUAy5M5dnO4EXxDG
7YrfKJI6QXq3oXlWH1qqN/ATi0nCzo8lkqbVxTiBBa64KWsrEQGShbmRtmP9SmAmtaQ6odq57pcr
Cq4b4n9Zm7Wfwqjsw7OYCX6laXqMzzKaU9Vtv7tjktNTzyFxuFjwNBVPZztoG0UYCI8r2gRUsbdb
MsZWHdiIstRWZypICSJQZfJX7kKCjCC5A+mI31uvEOEv4tTpnKWmfKs+kcPLdZQ7atVRjmS9/qk6
oxIG5b021SzQV+qfU8zsrjDyj93sjK/ZbxZ6mPWUsQK64o7O+Pt+JYsP+0t9TRTxhBYpHU9ms/4G
wyC67LlSKiiEbVjJLlJRjp03QN5RwBW8cfmfshqe/4IHt3hXwJy/gaURNGHx6BJu/bJ4BERhH5Rr
am+GWxYqeC5mZSEPqJZLCxsIQT/vw9JUF1PXZOxVVtOqbGdn9RFThHyq9ZCZMQAZ2asgiFg/BaNM
5Abdqtfmi1762qw7amoOzVjVlClAtAfo4945mgt6B1w9QQf10VFYMUWK9QIlVjwcqx7YmXjW4I7j
O+UFzA9l3Rx448XUpX+Rnjq/dfiC4NAr+H0vojEKnQGZDQ26DwtcTbmSpwmd1w6AbxMzEsE2KxfZ
I74TMHIZ+Ij1TdNnR3iTrKY2kEioTDLkeEUbXUBz73rrYtB1Siw7WOZTXHFot3m+dwcpk6c032q/
2/b4oOxX3rUtMgTJgMdGcK29N5fRd2PC7GdJMFHlLf3HPfTzy1aqKExW7u1v69iy9E8HoW/AQZo/
WzJRzUiyHhcOx66BlxRf4flqPcbx6hCRh/Lz7hCwWLjeuOWod8Fmm/NIizlx/G38K/oRP2keMFEG
RXx3Gr6bka03sBeGveDIHuHz0pWbZ1qTeDWVokELV/YAoRVv0ljku0AjjqLQxw2pjLg9LpUIUstf
djDpDeslnW3BGMjRmfJDeiiBKWdelco1xjSi4xZ7UL6tqqJk8wBJ0SgaxPDnNyr3AywISzZ9a9dD
TCsQVuTchrmf6nuhWkyGvtUzgwNveXQmVnH3jOArkpT+yPTxWMjMynKbrf1E8DT/ivITE4o5IQ1p
zm8RSInGDr3UnrSlDaooMGeltmhHK97M308KeoA2rO2w64W6ZCVCNOc4sjd5Xu3P0iyyu1VHX+eM
ibM8+bbRAt1+yN6OZaWIGgRoY3YnFKsaWn2cP/GS/1tHtyb5K6mt8xEKNBa4KXVGq63GZXkh6JaJ
TAnaeZkgtU2sRyteoELauiFoxFWX9rHkiJ/rRbElYvcKD5g5fgUNi2bIX0bu4fPq0wYlyQL/E3P+
Wo9tHZoS3NOY0EXLexj42nQihUJcMsHPF/p0JdAFZsIVuwKxfUO4p7GFj+7ZywSjeSErfY1Ef6ku
1KDkma9hI4WHZp0Qb7cC4CucQRaOVHCh3cdzhGLJbJp9BqQhNxJV73LqN62gUz2MMwyX45cVltFk
8kH+ciNdVEF2RtoT13GstnD78vRJ26NE6r2vWs5EG+InDvNZjAJRkOdaPSYE92NJmEFIfy2a7KLO
Cvg981ybDeVsNhWmMhXgfebwm4FJa43ZFGabuoCgTbTNyX46o0MYG9xokdWrvBHY+arAvyWINlkx
/4h5PbY+35cm3VY+Je2HEBCCjutKlzOF0/PkrsHGgw1CckDgwqOrTQKShXFJOZZ54OgRtLjLk7dX
/8mi+jgJnJ/EtkUK/yplmaw+CR0SyADWhpMu3oeCFZZeVYSvaTvsVCb4n/bTzJ7tEEHwEpbXmlfO
bo3Iv342oVF5M16U2MYp6eANlklnpplgc5m5YoMcWNrEL1dGDC9prL5WkVQyMK2BUBDFdSGheUf5
F0TXLCF1NQwtB1pjx/JSU4gD7UDe091lSWlX5IrFtGYjTnfUVHNAtyZtnS8PfuRo+Xa0R4N6N+wG
svLAsZj42lAWOM67yWz0sF+eNz+3e53i2M7/eO0pt+cgGt+R7YCQtpfO/r6sYZlkaeO5AcCFsaVG
vgxQ8Cj8fYs5wDbSRZQKc3P35qSolrdxH4uxc8NXuX5doyuyIr78fc4TDt13B2fOOBllz4FtfkWD
qixVz/j92zNscHaen0MEQQ/EQWPDy/pzyah8ny0uUfAoJrGTMU1sS8N9AEL4K81wDxNJzRPhyJDp
TiCVEGhuL1yfrf3PVMtjq24BMsQCOSr07b3DPic9th/HG8AXBic0hap3hfRSzIrCPCewsQox+gsP
U0V5drlHlCZ0slF/ta4RlN4Tr5g4hL/j3vSGjor1SidNBaYbNNHozRLDu3yn53DKoT5FSEB3nsc0
Ny4SEAMO+OtargEarA2B3VDt+HwbP0gYnfQwrzBuo656jakyQgaL8LLPsiEC4IQw0oslTdSeaaQr
d28cPWvm0k/oWGZVTjjQAifBf6mnkd+xMD+mCak8CBaNRFsP9zGkYfXisIhQLfLNVeoDPfyefxmt
CqaTPswKCgPBHykxBKjnyCHtGHgsYRYqD8ighHPbDt4KTxTpfW4Tn74P9VLu1NC4dtoGDVaQFq+k
WSDA+daESHcLznlpiNFdj5KBDmxcXq+ymxDGVKyUOe7BVjFRgw7raO01jqEtdH0v20DY2d0qyB0D
bV4paSqerjOLN2Ay/z6snc8vFZr4hRPGG2SihcROLdD5i/PCkDYwv0yuITxRVyK/n1xsVddFGWVO
0hoVmLudIj6FF/QEarQKAIvEMUErUVbaRxBP2tZGUBf8wwkpyOHnh8ZNojwdECToR6dXSgXUMblL
YnPXvS5eRuo2pnp4mnfjt+y4iK+5TD/Lg2SOWdLbsiQlQGeIXSglSZwDr+ShbSF2zvsZBZqP9hdx
Q/EgausDUmq2bxRn5iICvwoXgs9XsFQSNvWqdS+ILFBGXwO8O0D3YcdoSV6H/cAvNJ4Oqwkt5f+T
gPEf9qpzwMaNXtuAQObgvipawRN6ZBMGNW46mAknUdWIa9zhHp2tI/M1rEoC0X4bs/Hwh5KoFrYw
DMVNcpH2v5mCy2uIM/HcgobN0IdlRnks9OJ1h19nZGunwnmfMGtM9XUk8Jk5JTdXdgp2Jzm+A7ma
jX/zwaE/eC4GCAuMA0AtX7iseOYtf5o9drB64feWHffGSHcLnQ23LrkeWKcz1pt84/z40OpAlHfW
oebvoIbcgnruJ5xsjyMBvi4WmKTGHzpqJ7bKl5s13HuElkXZqjv5C8ybm8vkWWaafYlELkXZ/73S
MDUqMDOGcEoXA+DH5rCERpC7TcS2919hP4RzOer/VyKFt5BcoW8nKdFdmNKOlq++wY3HFna62nA9
FxUmXp8zeBmETTKq+17SS2XlMo/JTCDKzIKcecPscGoUF90Zvqq/AhU4EMW1dJ0ekHB2RUUeirLd
n0gueYQtgCPWuOXKDcwyNvYHB8itDALg1anhXO2Rx9yBnlFu089GPaQnFJvq0ASTPBF+ORpAq8a4
OHlnDbpO0EFavsW4GJ4oYJNfOo65/M+2V0IeVVwnDe9WrhLzEGg5h+zPZAuEe3gxHvb2wXxdGT9J
wPBiGY59IaU37nzVaxvNgY5yjrR+rWvYiNxUGMUcB3Z4MGQPX8ie8yAmncR0CeszolZzj0t1uCNk
Yx5Vg6nRut5kdf3LJdSopXehFOScD5NaOeHRCJjgdyS9opXafhah4wAJAlDIpAtK0bCiVlQS1EqI
Quib1k4JH5kLIYlMFPgOPyiXssLrb3POdqBlZh6A/b+z9YSCvCQpy/6z/a3+wS8wrhX0lQLj7PEr
c/0xUamwUWLWluFFr0FcPFxJCS50s0MUToJYrttD8EeYXTrSyCkEFKYIB+k1QeiwPPCv7ozm6IDd
bSMyN2sQlm++XuL4z4WJBEimrmMpE7VVm0eXoen3IygEZj/ashdjZ47OykYgFeHNfB+0kJma1r2x
5hIjlgcI9vO7cHnUtVzcEQ4UeUfLqC9+Dfak6FVaSQpkmcqPKRU4v64Rw/WZlgrQfLyW1xWvuMk8
yyd9uz+CZhce9dt9seKwTSsPV1SGNR0mTMf+aDvw9KIfwrI9+gDHkzawTrjAXqbvF7DkXTaCEMQ6
JBf0uBXuFtNxc7nSigepR90+bkJMI4LeKUNQNrK2DzboPD1tzNcP38eL0nrshjuj7cfHVP5/VzhB
6cRolbUbA2wBkMbZjgJxLtdheUDLJvjxbEajAKVRTRgK9ciR0g0WguZjtxI0fYneQ9NETybfPifq
gn/b4bmEJMIqKMTJEucKiSdbFjRr6IzUWu0ZA2mBhK/OdOP7fgK+1A6b96z8tU44CIao2nTa9iDw
Mtmb/NVlj4eULjbfUJi7+jB1pFmq6X4/rhLMIq9WVcPw4XijUy79QDF1B/261oTQwyGUy5UNgcg/
B6xz54IT5gVhEZcELEV/RI71I1pzdQ4TrW6sSDFX9UmXP1lH4DyUu5YDDt1Grh2miMyBLkbIc+O3
+5aBmZJ1V+0p+LOgv7ddnormmiX1wqHAPbsCqJoFQcSQr0YMzocE30ZRr7SI9Gkl72Wr35+Q+sV6
lIzBUVsNBgw61tYZHOnl+eVd61pLGGvwXabgB7qye4ZnuJuPzKbbHRqfGP8hWK8XHsSNZdf2FaLK
viM9G4GyWYmF5bYoSqawEYoKG0t5ymkFTZDTWbBsaUXmCWkxqbH1OhOkvSRRefk5hE0W5fC2x6eY
1R4N3Yj8vk+ntrxACnC3Q68uXMS0YVD8gueiMcsIkqNkGSmp9hnM2NkZGP2hk2YfL3cDJ19fYr6F
5B+2A5yjl44iWy8dxj1KOJXUwzp3lpoAPpdF6HUEKpi7uOUQpmDYgkNeaYznUd3lDU4Nz0h4HfsL
3ybxrqfnkYfjLDP8e1LXDo4xI+VIYw5ahmyawovBQtHIvYrqhYHdQN74U5H1Lh19g5oy+HUafkWY
9htny1uoDvkO8N6YAre/kv2fTKeC/S0JlHtWoWRkSq+PQBv8r4ZIu0WarhB6MaaNF0mGHOoiYelH
6v3YLHEKRA/ykFJVdlmXfH489NTf1cx10QdBHqqrDAzkujSmQ+gjOzk54KLJApOqxR0R6l9hSQN5
U84BJkBcuY0bJXqu2BVXc9dY4lVx9HtmPp3a+VylF+67/R6ZftIeu4F70hXfqwPixGwRt6PG/vx2
jM5E1uMwXz8MFcv9HF2mG/l4WdX05PgE2xheONJBFt9CuUa6WBujMMc7WOUzz/+El6sjfPg65Wki
kJQH0CdQ4TtDj5MkY4s0hqc+vcVdF2GgCFwI2sjo74mMUAit3OAqh++454PaPVRoUXYPRsgOPte9
RPlBpS/5SBT4LZPT21p0phcsutMQkbVcQHCUdGO6LSPt8nCcln24M+HaJwH6imm+eD+LokrJmSrk
Rl4T92q8RHNIjU2gjXotrN2KK3j89/+a7Ndiukr/s61YJihCUl0yH1iE+/9CDal6x97B5qeNlMYt
wl8iOIochy0zA+vN77ZVbYgeu9/Nrg/uck7qv26vZc1HBrZPp9dYUgDmhGhOQl+sgd8HIyEwcop8
TYfHYRfIht/pVQtFcC47UjyhZwG9jn7g+iu9pnNHB5+u/h46jyhtEEWN7eh+Ck+MwHdzqnDzUbYf
8SPzf5GXgstyI2lv4IhNupMDstmaMoK5/JaW6/4TotGX25cfbpOQ8VZZF+1cvAvyl1BlGQVteA+7
CAxmZGWflNdt90Gg9RslxutidwFDDArhVNdaXUkRzrp9hgigd2o2oEUg3E+f/hDphc2XZn5Rw3Cz
SAZh5sIYuvj3tfxX76XRszG0cajnq1WsUtG7b0tbj4/OOKO77duWKNOXJWqIrWciI0Cg8sUnXBSB
ShzspQONlfTH1GES2E/MdvGw0kiggpJLuPl0dlprxR4EH78lDeKF6BhFSQtZsuPqj9OhfWcUCMiO
ObY10eaHUSEfjC/uPO8XV8pJAVTxkeLVhExyGkQlXwT/zTzA+9PbMa6J6h5MsSO3XpkVG0LXjjRp
NLnsGo3uwc5wgYmQqwx+NuYr2JtKLuDkv6FB62mEz05H/yG3EEZ8NbsXwpkSCwud5OFE0+/uCcHl
jRqypzGp/lugQUYkgIOe15TTDtBymr3WCfBz7tVAf7goeMPlrWhrnKlyyqh/4oE7XjeqasrODDj1
8L5v3WW4RBejjKOjVfkCnUfkFSP9wHZtRSQZQK1vaR6In9PK8WQi1c7xn8o6mU45JX96esSqfDnQ
ubd9g9nu1qLAv84V/c5u1GjFLDbDyvc0FUppPnTQlLulGujAj14c1rX/cISTuu06j1iQiZvG5Gej
kUHyl1AnkK5FzHI28W25KrC1l2u9JD6fwj0QQCwpLOHqipeVKCr9l+2C+Y1hmmRR3RB15hOENbsW
vQzDKj7iZgsqXENcOanBooqJoKx2gNNKEig3s+zEc7YUisX13ygL8M26XsAu5aYIDHMrNCQKXWWy
LjbODbM04c6jIsg42zu9D7wKvIEwgcGcu6ELxmtrkxlu/poR5KcJH0Earva13Q+ae3LL5VnuAOvE
QQBsbn81pUhPqBkz0VPpzFclSR3y3XlHvdFvohXt9k6m7Ivch3Z+YExHndT7dEEh39MJogChgwsU
Kpe7W/KNyOHU/DEsw4AR4rhTUAN+xjgFklWnpsNquPN6rZPlHA8ZI8/3gYJyIXkZdxsc6YAMcbbd
OpkmcaBx6P3notmM27juFHAmER9PE5WBwcdp1nBXXTqJ0hdjGXFNIh0bnf0WZlUAT4f/CyOcXY3X
MVuKiU4CEHeXQ86N9sVXhjtA1lmOzQXSwVja3ONaYDVrv7yjx/CjBirpIMfIObhc4cMbKhjzVY+O
hLa7INfO5vzJjGywnSj9q+RgsB7VIBI5PwDYFtS3CL26hm0pwRPZS57V5CpThtovd6SPjtqqxvKl
8Kuo3CtkoCYW1gBU4dPavlF3vFcUvQ5O3qeOp4kPx/5zQfz9KjMIHHJeKG7tWFC8bqPlQeQKNHgR
cawRU4g+vUBA4LVRBNbrGJYZ3dLDh9dF1TaPSMbASH0Q/ivSU00SsjDoJWo2iVB6lYdq1tOpF6lm
eoWJxnDZcmCmU7wK/AOnj4gLx1cU1OjOUhFmLfIrof2xdhYajr4KIY/FfGC4cOiW9OY+jkVKyeBJ
l0mSL0VuhewCqufuVYB794l1Ri+xq0vKcjnbW76cexZFEVaes6RQ/H8A/JcyPqcvM/vGZZ4v4RMA
dojB8DoAANjFMxbD/sRiA4MOp6YRNVzqqAiwHeUBmSyV3zAWMa2GTsMW3Spxcbh0xk2DyKe0dYng
xEiTjcfLD3qK1Smj23pG4TsF4UlCDHx07JRbjST9QY/KNYpiL5zEYeHT1+NaBa0rKm2f2IWrZwat
vXt9m3fYQHsAqxsu350OC+Epunl5rAGr47Qbf3Cuk8z+Ikdl56HNIO5QVV8I+tQjqgp+6eFUsG1u
EHRvI1tb+WAZ8yQvNhmdvj1JathKhYpZOoVDxx2iWH150dgju1LZVr8+hIovddAdr2LcVx2fDWbT
mq2aUMhxae1tb8HRbH9cJ9Pz5m4Ma4GQRmhvjy9x7Eu4MSzgXGkDC6ali9iagUqz/Tw579YCZiUi
HotJxpKdYGt/aoDXGxWSm6RRJ33oK2A/Ry9WqlaPSukK0lMB72CID4O1zQfQvdgHcWVX73vnwcSP
q6O9h4st4qkuuCmpf39u5IVPWeVuqXG9T4JFtYBeWmASIXJEyAfviMdT2fpzzyi6PWrKOkR5F2mE
t0+YHiWk7hVbgCJ3W+G6+TAgiOd9RP/NLnual6QWsSuUgcmSULZIWVtbaG1xbpOTpCh+/gjKDwnY
RIyWM526QRARZqzuKVcMQ/NpSdoeN9uOn8UxdTvYiDpBFjc59ZDmPpZNil97hh0hMjaE9ZFzKoe0
Hg1fE9AekvwMXLQw60Nw4KSnrt4B5hnJMCSBNJq11yo+7zyPFMSmlARLoWaKf3Dysk5w06j/6CuT
HV6pAOwxkAvg1Hfb/aigmPtXi3z4il48Y+32GfHFscAorIJSgLuC4US7vjU6rn+80YyO9w21OT5g
7xoXjVxCboPBv4tjVN5etkOVBDS7JzeO8oEGbRr+T/cJWuHgCcqcgX+wKMSDDIlD3UlTBZWrJzwI
5qU7wbAKTYlIl29GPHM7WhsL11/Mm5c8zuhK4mncWfVzA6ihlpApXvwAhs3MLGYmIs/0N99UzZcM
fZsXsE4c0W4i41aAg4WDv7PRfGtBBk1BOjIpKRVMNizmlyfwD6fNgpz8+OgnJxmpoPQR3BrUyH0b
dAfXk0tNdXLfjWZlzpg0yaboNGycGDSrS09Xe7wFDyIcaFNgZXrJ7goXwOLEh54a0FrwOP3EfaVc
y6W4D8UyHhXmZpJE4+TXHCy8Ybv9OmJTkikPdu7WMbPkNIW06MAuLj/HGavZsgshXdt68c+Q6YXk
6WP2xmkzzTGgR/oTpysiYh2BxpLFxNNhL9/ttkRlTVUXYjrpUApdqfl4XAh4oSitlhXcjeHOaQXa
AsQ6ouAqNzDkLqvkhRf315B2jF2hE9KjJ5UwPsHl3lai+6yWU1swvJ0cj1iyx0lXt30jVCJnAON4
46FYLUJPs9AZU8Jj0p0aSE9+R/fJR/ib+O2gEKVaZjqucvPQhxF0mgcA6BQTztl+Q2Rcuw/GtDhz
d4opoMIlsArSBxu7WgC518ciei02vGte6B48w9Mn7m7cMaEPYEJ27wkcof3abrjztRwGqeqqPAxk
nYOXO6kdk7gzp5DAV8ZTSNtZ6mMrUpIsoZIP4sDCathseVZHVd1Yzq3LxhewNCSJTIBAfR67Zwk3
IouZId4XW5K1fvBz4W3U1DHNBigNX+zZ01pfgqcE5xzHeM+T4g9CJujgzgg4iSSRsEysVrtUTymv
BRpnw5u0xoh2V9UM5zQPerJph0pAEz1eiqeGS+vTq3h+Kq+QJ/FbPNtVvg9flSV4CAIgYypyetDV
MZJCQQVcwWaukFJb3aVq3/mDB+pgG4I7g99DluflgySlPdJrTk3WIsUikBf+g+im02qJZZlSewmI
ImClsGuQ5zJM6Ao6L42YE4H7/nEsrGKWUgAk9h8KWgnWXRcWucj+Dwr7lfaNXK8uUU77GBq8uN3R
mmZ+kmymJBx5sospVtCF+sSKhqYm6XaB6SNNLbiREn7ZUcmZOJ2MJSwmdPF2tnoKJi1dl1LGzcDI
GhaqxoLgLBiiPm0qRrqGopvLZJTIEMiRqIoWf6QGm0zaoE1RoEbWleS5Kb2l6D9n48AEJRFaoK9M
Uabx2hPVeKAnZ9VPQcfQUYLN4DR5I7t5ZGnrkIl3E4NgXAlIDMCEpdoi60BtPhe1uOhbvQq0+c01
BzqGf4L3lLISsjyc/+D3S3S98Noce2Nd79IcKQ+4QdArFWzu3o8YEQ/uyAc94+ScwiP1wbQTuyk/
cr/HvAzCmqneQeplyc4zvSXAIB2J7Rf70/QFaeMPWa11yvbZbarjnzL0ekcB6YAPKkRiaFuzwM3+
oiagW13wg28RvYM0ltZYkRosZ5F1vAKWOiYAOojK7jmFPa3eWkmZpZJUjefE8k6TT8HYW2dGEDO/
hpX+M06lOnobo78dTKB6NXmfZ9Mov0jSr093PIXxTxX/NkzcoDao8yJ3EGvGINldq9SwZ5wZcB/n
J5qwe/rSrFlPpR6R4MzKlLb7NnmMlQWp/r/tcAseZn9SAPSmNUGZ7s1UmTBsrVZ3Nke0a1M3jv35
Xb0K8W9eKZKHnwjcxgnuDAkz1KNqEJO77ZvWWezun3HI8wbtlvZ0PS2UVaqThqxyG1Ocxvsko3oS
Z7G+rrMasJ0jI/1EJLhe63iypChATwZ9MF+3ggiBgPi2cEruhS+iafmVnE16XZBeK1gxDZnpmzpk
FFjPGCtXdxrl+N/eye+g3Sloc8Onsq/W4YHyqM/U4yzi502NJ/VGGnEL0jcZewvzEDPia3TgZCMj
ozW3Od0um4MqCRffYNrJ5IkexSLTgAjCepUbuVmsbLWfgzijH+B106Kze/sqDLNsACv78FcaFN9N
WqMTFcd/3/pAgg4VS0lJbUKDfS7GfzuIMN59D13yVC6zpEU5nkDdN4q7uDriVv+F3kFxBRum34Fd
hpM/5tdQL+IypfIr7WHAJER0yrPYU9XHCb/7gWxoPQAWN77jlB4ubKDrKWmHARHD8EXuf2nHRoY1
iyjmkAABGHWFHnFbEhbiMTnah3ag0uxsy/oD95OKQ07gBN60tYyA0XcJGL67PWRTFPNG9zX7AKrC
mDRMEfIYDAxwqu9TuMGw9c1NedexmPjHguViOB229tV0MPwKZcpf6wkxy8nI5B7m63GH7+CdlSWn
al1dd4Upn3d637lAy6FLE7lisdpYKR3BNaf7agJIqK97EnybXmCiliO2AygG9a7nVRAAAa5POxuW
9By3fTOKZFaNheuqe0O4fkw8/A78Gx5G+cl9gb53WaniRPS9Bl+UBeihD646owcF6eGboo5og8SZ
XXU0F7sIJmnr4t7WnOEnwsqMRoPQbAJ0m5AvoyFABoyWocNMFC21QWoMTT/z14qHGq23zGmvETwA
nVbd6r32ay66G/6fUAKuelbxEkIOC7afaoI0afHfVkeDK4u4X4WmVuEIj3q/4+L9XXUNIj67u5O7
XpdpkK9cvqPYglGAos0l8H7UEQn5DmZpPxo1ddOtwIJHFepejD96e5xdK3uza3rcMWATnjFzzQ18
5Zmv+IyOyflCR0bWrBQPcGXFxdfdAufHLOixu6XjRDgdqgj93peLv70BDThp+ChFU47f9KaVlo9U
03QiBrh+xj5gPfy+8NlF6LbFqi05PanKmoujM8I8rH94NShgnvhSzIH/9/S5/0PZzTmkoP/YnYDA
wVOWZJGvfFpwzseehPFEO4+MaDs5DtycKOWk7hh1GWHjrdn4C3E7l3/67Svto9sMQQCjqyRY06lD
8RencBysBZ06b44YkBAOkQ1epUCTCHZivqC5MYQZN9vRiH95Rlfau8EpvOCsdSYNtc2shOkmgMZb
H578268fPVKWdzEN4xAjMiSK/A2Z0Zyoe7WTDbeqryTaJUk3n8dgOBVE52NB1fk2371yIaH75q+J
nWAVyqodnVzmHWtdW2b7phZ5Sm2xFsX33YSGIuyNOtDmSBeehHpcG6qX3SgLKbqTiNhUjwajMwlX
kNmvBYcZTwpO4HUBl2RLnAT7ebKws1E3HcyHWtPr0gX3cEhk9rzbpeoWbQJvOU26prIlii83TmK8
4vtoYY66ygyD35QCI5XJDPF9EcbNl690d3AlXKPEbGQ5p8Rjzbex6Lsz7MiEl/9hjSabxpYme6ln
ZCBH+cMBOJVzoJxE0eJf3HwuutaHQgQHPLf0HHLZ4dkW24H60FrvgiYOt4eZ7ynTeh6XhUbj8tSe
fG3UCCxh+iCCuUDjsLtW+Y9GEImkk8iI/94WC5w4GffyIK8tjpJV7skLQIjgNkxjbF/gOFGT4ReF
k7ysQOu1FuFi96OsP/KjTzuike92WrqyScpvxA2EfX8kxoRuXNr53+6NzCEURXqLkG0pbhrNI8g2
/9hUtgRbNAocadDf6+BUpT219hu+Ykz0d3LS1Yfk12xEzCKHWzonRW/VIcW2X+pG908FYNaUQElS
Q6Bd71hIpFcDokCA137E1MJITIF/BFt1STKE+nHHroq9wO+mKGDGCKmxVVuKMX45fjTZGOkGu0nk
+hdv0sshbzQrXXoNZpF5LYDeoxVDhNaI0u2J4GfCElbLBqAD/K/nOCNg8hH4N4pMoX27HAcMJoLO
uQqbxAXcIib01Z1zBdnxhBaQ2CQ+BXKcZ7PY3K5cOJ1JjVfNvyBqW6MBxFRL+80CYmptO1Y9hwqs
tjKJFsQ8uAUasYkIUKmaxkOhpOhYbkyouMrm9XxI6+w2M8V3AAUDIo/CZ9Qlj2ACQof52o3lOaFZ
7OS46gVcSRJ/Eh+MalA6un6e8SLOF+ewnmpsoBOKTLXYTpfchxq5hiwNnfxt2KFGrRQhFnuQ+y+Z
zRd0Ezkegbdf4JJoHZjr/kkwZ6xEfePjG5y4mKopyBXLaQfFOTmbBPplmx75qMzQAvNTJ5DW+LvK
+dPjTuEFwAmrpvuzg2PNKNbPcY7HuuhP5F5bpbdk0hu4moTxiUHAbc/wS/hAgnqMEzUT6xoA8tF+
GLKTYL8vjcpY8jmUtY14gaoW0waxW1ajZwFXQ6ar+oowqObd3buYRDhl9W91S5gu6OmJD+880kFY
GHgxbBMSCq0iQhULgchrflYrlvO2ZJzEMyAE1MntfkOrJugeh2lIhJR5fIj/Azzh9rBItbeIeIR6
czJpHJWzSn0sWKxjA85H9qWCCV4MLV7612bHzK57FYJHVCL5gVBXXYzQXNYHOzXbRrNzx839X6le
1KdLo5tdcsGAPggZrz/mQdMvl+6Z2xjYlPZmEHM9OQXJ+5LaqWk/Ajh0xjnJWjS3ZQ1vES1NCFFN
v7Yhw0ZHNnq3r0ShqcJOUbCPqHLzU9iLJT0ufqsXnWvnevrjuwXV1a41ffM1kAv/71miypjGEdmF
YxdT4J5Gy7saAKaheqIaHe4ur1M7ccqyAwtjIaDaqyk+4PHGpCyZ0cDQ+rtcokUamwcVuTwel/3J
SEU+s8kCfBIyp3Yztu5zPE2tDU42bcoOtofIgJj/9n+F5lL0+d17LVKGV2iksE+GGv/9LHPRcI1D
oKe3QHRiWGq7nPNwzQNgd+8kH4Pa1+hosVGneHEL4L401i7S55dMbrT0nJ+oNeuTLtEHMf5LD9ri
ahhkKzaGIcAh1J1AGfeqvTCFwSijZk6HP0PKZCZT+/Dh95DpPaPcMMAv32BcR8y93+bnTetP5Hd8
vz4D3a1t8zBod/jPe2CQdOlQPFeRKmDFJwFIow0q7p+pWntf5zbyrlaunTk/A/8jky6i86WKEcOe
EdChXOs5CTc3BvWsuOavvWXOqslLboevdwpTnRIwTh1bFVKefdE4LchASQg9uZlt0RyNsm8GY+g6
U+dAX0RHmeFaNqGx+Ef7+XLON9HfEImMu+q9hMCW3hN1GqgvFO1eEwav4wYffecXkg3OrJQCe4xK
61dltR1QC642BKNlyWWiWxCxzu+w0UQAzlXLbM1zUQLLXLz9qhSGP2X9YvLUlK7DnaeCw6D+2ymt
zeuTBA4ZtNGZB5GufChRZoeWWdi6XcJ30sbGBqilMKl/Dwd5XTn5hFrAU7gfwNyYLSFthw8VWF76
4dmci9ZBSaqFb+KY95tl7rrBe88lWbMo1pYrTfiBEw7fDWax8NWNh1WVLsfp0NKYgpY39XJx6HM+
y3QjEJXwU2dLxG6388aJDHLtj6hx1KzL638wUFK+2lttMqECb2QaqTAMpAoPJr7Gz+C9zX5Cd5E2
q/ucsSLKjmEW/96/yl43aDdmoueExDfMBnyZXW47AJe93ZjLxzaKZh6zUVBC01Zdn8zyA5UIxxBq
pJrLAKdBIK+a+E+zUoWkeSai+YHab+GhBxAAx0jOSl0tt4LnRV266GfMS1VVJbra5cbE8t2dYWez
y7hgVmgzKW0wodfox/fT2I/JwlkIR57rd/ARbCwZX1xy07N53XWvggwWMU1a6WZ0hRgoQ4k4ui2m
5khu8ODBX8bgcJuiKWQ3H7+26HBX12gd0YNCzG+u63uG9zdGG2PdIp1dzc/BvfHHdtrZ0VOTe5Oi
r4K3f931Vn08nXi/X9DXMYo304l4HkwvF+pV5zT2tPOgqHRpLot+hvcToGDRGHwnR+x2+MCndnRo
5AyjC11FobIFWzG5Iftb7OkEP+2pTHMRjrrhAbopdM4n04lriVWM401r6ilxzE9nnTEo14KZh+z3
1cN7yGV8Qu6vJo7tPHAfIdDE9ERi2BOtEKBMLicyuZbb2xR0PnAaeWYwly6LGXvdAnx4837ApvNI
3px6yvlcGndagMdUTSVLrwtrLvazYceQ0qXVq9SKjsLsIqLk8aHqD189OxLvLNJ8fZHN5v5GidwL
0tgSCZ95B0yybUGzVpCyV6USMPNdHE1cfyImybZQVuYfp2Qz9G+z0/k+UmPBmz8Dn3NQ6NOfX9mx
jgTenxZhn/EqBgU10cZS8yTZK9t7LLWa1XerbpF8FTdIgI2nnpeVXGBAq41zvd21U0Cvp+tmP7Xk
8aqEYyCi1MhqeoojpRc2PYsBAM6jpZT5cpSupoqp17T0CTwICBEhnchQziR/2ynORfxiA5R4aR+2
Da15sZsXMYgE/LZEOQ8QOlBKCi87W9qbKY4rrhirwRichnBebJZpU5xw630WWeGH7xkeilsferKa
8cNceYrlVfRksziOhOVhBXvbW3B1C+NRldROFL+9PnYw60XfSSI0DaDkpw3fZCPGkCYus1ZB0qSt
78r1Ae82XGYtDLOsGKJSkSqXEu9Lr3/Q8iOAKdxtCsRyYpSomzsjHywdEkUXNIq6iMnE23ybSy67
0IcNMkG6G+Pp8P/ADmaQZpldqbUXhuLyKc/cUVAtsPbFb6uTg6sL8+3rq2UM4dAQzqeCtshTVZaH
dDUzzhNXKJUrwsJm5mhgTfrsMczKqqTJ4xwztGuMVIFVZ3v6M6NNMgUl+jSQxzYoS7HR/NUq7HHj
kjg+8lnPn53BPmj6hPOmhUtjlJehR9MKIsvYc4RHc2HTVkZ8MTN1wfAVz0aqj7DkyylcM/oTuqiK
HylZMkNRMjgRqtshMxQ272TZugFGqm3fi+z/dVQ5Uy2vOwzyC5QSnJxoXbGEu7AqqnHaZRf0FzlI
ngunYNMZE6pPDLxycT4GnbnG2pcOjzecoXHdMc65HL4UU8yxLBY2pjRnY6Ri+JSJLqLfaT6Qee+Z
DmSCdPiVD1IiZMr7CobAalmKAVkwj1o7eMuFNi/K8GPvl8rxnZo3SCKPs+SV/lmeYaG+mzZaL1rQ
2eNcjmXINVCyV48zqjrzVJ13Pq1sVqS4yrRsAgY4uasX64pXgQzz7doU3shkYajQpMzk1s6NA+pJ
DHi3krwF66iAa7VhlrTqu9jJK7eKMLBrN4T2I2o0n5Q17Kn6HBGd+go=
`pragma protect end_protected
