`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3152)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qMfody8nr5xJtxmeslkpjbcyQ93f/MlF9rFqP6+2wAV+CyrXaEH6OT44
absZMXt9Ydz5aOf6Lt56VB5Yyt3x3Xo6ce+4Vm3ZgnmT9uXqBk+MP72amt5sCX1bEcJjA/bX/jxw
6bLJkw03ahWkyP//igi5gnRA6yIKuxaHW6dPdXKsVB444KyjSIu794Gba2JmBLRwaUMIYl4HKQW9
M9nji6HmIQnlF9E4TyY9RJq4LwnC3vUUvkhgMBI2Z0EcGDj3ZDAl8WWujBufqWrI2NT7QCBvfcNk
C/no8e1uMo129iWd9a8JWQYx+bMsGnMBrc7AvfNEw9BIbwzsaYoQp/xUVWkF/rBSJ4iPIX/fLemn
3rw8uAd33jDy0vk/9b8gKQE/JBqNqZUnd4PyCGidWp1b/nTmU/vNcMFCuSY/+XTFzO7kfnj1Zr4V
oMhNhGmm6x9T2iWH3fJ/avn7lArmC+0AOd/eMhzlIiHQlhya4zONn+Ud7BfDE+Z2ZbHbSeBCiNE+
Jab2jcP8VahB+yKojmp5FWFkjruq66YkKrzpAFelxtDv/v8zZva/NYx/hNGZ3hlQGiGRnf0qThCy
/Cb88Qe4vfqoCOJssSttV5e4FO5KuGWUu2OCHoTqr5PbLkt9Zm722QmQMbiKgSNtkojNcvCv+Sn0
274u2+6mDCKm7eAIZtPv5i8M4hzDABLReCEkDtGzNqZO7HImAzfvR3hnYaMZZvBkBINYCgw1ypsR
iDCXhwBx2SjYKHWrvKwQFEJBJNuPIL9KpTtCgRp7rvVMhONBr6XafxOJNXisas9ryVLyUXf3mRkM
eXVigu/zidkwOrVRH24oyyIPeCGhunXMHVTnDgQl8rzrgkZk8gPgIfawfF1ucUzDOo/ni5ogrGGu
LT0EFrAITHNP+UiQtuWMsFyAT6eu6I2bWq5ZUmGLOlgoO6CjDJdFXYhv4s07jISyxTVRq9gMIx1D
gqhDvzsGDBjN0xpGVj2EyMFQZsnRnfShf4EVVCE+uFabq3Uosqc0uIKwGzhZedzbTBEhHCxHmKi3
n9NXCTNpgxjm3+rT2uiMZxcTHrc9suo5MmdmC3mBoBNd0wMgbWHsrlZMgmjn5q8bB1CgEFDod12o
6dgjH3mcNkQ2cSpvB8fOmrD/Vb2ekFXU6PKN8b66O/tiQ0Ilk1SZdy7wtiT54scdiFTYufzK0Vme
9BERXuOp0dd4vv8Qt9ZAsE1ygYalpIdtEalmqCgZrNz4x3WiicaCzIlfC1T+AN/i7jZ+g0bymOut
py/PJXQJpP3IJpmuvRvKwHvbcDR39l4/uyoQ/hh58OSSkCjNSdHedUIqOVinGIqisErC7vRkH8DE
al8pN0mC+IL9T+aIo+hkVNUSyCJ04v5aCUHjNhVJWLAjyNwsH3pwLwWN2a3gIHrP6z75sFg8X0ka
f1f0GX7Tu0FvqV+1uHo7W+UsQHctYEd1/oFhNiLaF3D0VmAEsjZo62CA45KuMvYkfD6PzhO8joHZ
sAzXoEUyscFSiSuwVnwaeDbJFTEOEMRgwiqw0dJaV/OCILLSJmJt+Ta+zaiuuca0YMz4LnQk4XMx
44GeveX3YL6rqpXI6Wbz5OoM6Au/dvNBR7uhpigrxoIB9pKN25wuypJakQCMxUYhfVBnMtWZPomJ
4j/GVQaEtprEQDDdk2g557BDbtdTs3UwOs5pUSNUqBdgQ0q6q9HEDI0dm3LufpjI2i7flJxoPH0S
PGv5gQQkCJ+IOXUyrg+Zi74ZYvc9tZ4foJXrSMrb5lPMis3G0vNI3TLKfK5yyLIq7S4BFWMOVXrB
BlAUhxTborF5/a2ZEohzkRDYBsOh0rkMN/aqA6mkhwVcypTxn7c5AfmU1N8+ZAyklVXegXYcAH9I
yB1G09QyfpvBkuJc7G1n2Ks+uIwkGDe21VjdZU0xbtg3qBIUGDWqYmaiA1abh2+bRKrztnFMWZrr
YiSNeLe/zs56DcUUWC+4pjVWCeRHl0LLcQm49D0y38bXE73yRVFB+99CR9mjuHNhhEGpHVzSx/40
WRM6G+ZXDvjoY288gJstK6I23WYWpe/euh3WCDnHQgKRy3Z4xuiHyr2J/ZCHnJbqFu3YrE/XKDZj
MZqgBoD4MYOR3ah0u2Ts0sRc3o4gXL422q3EN+8xZ1mcU607nYzMtIoqxduzudd9MDD7KCDEkRiO
DSw3NZfgmIWXv+HuSeaFnllgO1xiGf//q1/4op3hVntm9UuicdaNRvJ3MvNuuRvJPNZE7BLhqpC4
5oxWMmRYKoyllvbAZa9aIwCe4b468F5MUHv3wmWjTXkij/HkA/PHel38LTSFXmarvIqWE4oEhrL4
GBYGcDtZyi4bUKYsunVsaMTm29i70lQVfmPI9VBqM0MLJpuTp37P8x+WRj8Bmi3Vp9JoGLUZ8VRt
XCFZewoB+PbBpUrYPt2BJZtDnLRHIBjhsILilDw0QJrs+MDsKPcw2YtID86IA1FPRcansylHHRPq
z6GhrEMFmQ1ShqrxH4YCIGOxa+yul2Y+85Lvt7dFDS6PsQh3uUDEA9T7hjmNKD/tBagPXP8Xn2Fb
YKbZslbE35UqBVmYqVQotN3X8P6+rXlyDcGxzaSxI2mtJ5tpa8eDEkHfLRUL1DKexDZCQrtm32E3
PrscVCSmgb2j5HCu3X2BOpdOvCqHAsf2Z5c9Pd0qbuiYrgPd8Ve8A/TBTapEQblRYha+gAiLbEi8
PCwQtN115g3i5rF+/cD+tk+805W8ZFtxedcyM4+Q9HJKan4kqT3/10K0bVokydbRa/1kCAtzdE2I
othbdkJFTLK5r6QdVZuEsgDqc6HoSozAYxQ61iGWEj6FmHOawzUtSB+fWvczRp/wGhfX+iMGNuCi
3JAVD22I9WFcokJvZMfNMdoZIwiCWCcMUqbs5pYIwZ9XhRu2e3JysbW6Ht4zmcpDpSeHAEMMfAT+
3zuRVd7LwAcyEcHzkk/SxMYuBNmNt3cEqI21EWmKt7+1ubKftr/1xPtjkw0Lfjp2psTCen/ulu0b
WLCjhJprM0tu1CSNxMQ5ONWLpFR5GolQFJJkVc0qZSMPIMc2+qJh+RdkbrIRp6yiWKdz2TDS408u
5XOmWhppdj4b+Dd1g9LwLvcFTUMkeMNuHrQrhK6oubvJ6Wn6wjhmQ6t1zcsZAZHxJObQA+1Txeib
wkwJv5ezfNMHCV04X3EL3ssVPC7UlRATrmWY8pr6tLZWHd0cqeP3caQZU4Ok4HGIE3vhh26bsO1X
dO+I+cmSiolIeX/mzHFxqjFIyesfhG97vHCOP7DYYIoD2UBin3ZyQ4HUC00kMGsVPTmMjBcHlBzO
YsqCQoKLGJbRIK/x1ywOFYkihzIbFZsrEYg+iFEZ1+eTqiXcn/EpJB0vovNk1L1T6QxkTnR3K/Do
B3Eq2g9bhqtUnuQiPT3Cgt47+pp/aPCJU9GmZYgVNLam8zZVChr+6tuQrF8Cqfato9QVS2iB9nqG
gh8Iq7OkPkN5/orY3mVLy7PJec63iiPYuA9Z+NuBOlvUQOIvxdVxMdDd7WzABi//Fi4914lmM/Zw
VYH/OobRi5N28RhvN7bF+LVBuFQ4suV3EPgQy3vbP+5/zE0dy9bYsPhguS3WHrl0C7g2HLDV4Nhd
wJWgQ796t07CgLx0yM6n+Ln26fFeRonKRou8eFwTC0HzQKgPgiuVsQ3nKLxmA/W/Yzykz4VPM9LB
E4cer0pPw/Ea56XZhwjhZg4bTg4hukJbM9wEcjdsxzZ4l8UpnvsyNDMjdjO1eCK17Ds1d7eNOH3F
o9ZPj6mJlj4Ywbqb75MnHyum/ZmE6W5ZJ1ZfT/9+F4v/NpUBgOKHjLH1eLzDJwBltZOk2h0RBV/i
nSo4EzPTmftRbmAxYLvNF2+mwFVtxMbcC9/K/Dt3VZXzCsQ4bZR07xAOs1aOc5EyNKVJIq1nwNzG
0yiKe7Eep8PM03MAtOX5149zN2L/qFiGULqcpIbu0CCJx5c8VG/TWPL3eH99pDnhl00dcPPZMim1
Bhf5r1IWKxSedPf05Zg12LWaAwFFT/4l8G4qTAANg/PSirddU2e5lY/zkFAfXCpoGsjaodeaHFgB
S1VlVLktsxbs+SAB9aLpNnaA6Kgy4zWH++CazCDzIXNNOENVfUNjK6Uo++WkdHaTxC88ZKN0e6d+
Rj/9NXbtWC4MPJt/0KS5ebY=
`pragma protect end_protected
