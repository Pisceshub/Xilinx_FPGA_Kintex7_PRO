`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16992)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9MVAJWDJHNzPOTKFbvhWRW30e/Hobgd6wCu0QIypve1yV87QmtGExzBA
PSA9vB1o/Vu75Q7nhs4U6VHe6gDjDxPWUzzeeE5+dd3fTpPNe4LZBdL0HQt2DMpC0yVoEgjjTX7q
c0fJDftyKrz78+yTtH9kDoEyVLi+RQrYD90nZOoiDaf7ZgY9o2NgPmoN6ETsB6KHz80U2SfqAFih
E4C+uQI85oPX1A/UZTR6qEqbMFQRPSpRv62/pKmL2o71SSt1wjLSBMkMirZ0hepKKMsuzp81vAcd
eQJ0oC6WAWLqjVyhH/jB3XvOKxjWj0ZUgwsfCObYVo6KViz08hJLwZpGZMaTKeV3TvvlgDItzz2x
oYZ7JcBkW+RnC5T1o+p/TIzJhH/nbF0+ozYfMnJeiqVb83pn30lFs3qZYWgheL9RK/Yy7Pg3yoqi
nmXKvRBd7avQwFuI+TcUWdRqNOYJvH8M+YKxt5AJ6NfuIePK9cd/pnDEv8qsSDK91UzeFDodo07B
lB2xndkZ/CeRJ1zKBdZtiArhnUJcavE/y4Zee9aW3FSAUPmOsulPv3rdLMKCsEtKwIaXSNI+6tC2
45GwbbP7uZ+qb9vTFpLtFQJOlmGiytXaknuzlh0tgujd2LeRsOpYl5M27QYRd8Q+FatbDnVBl4X6
9HhMwA8st0Im7Zx0FNHFF/OFPp6Cjerm7U09xw++WxBenPIeeZufWrAFeMYUTg7zlfHN7+gj8Fef
JX7ob2dtqKmqaaD+IYgogce++KDaeZH+4LDSOxEjz3MvW3IFTHapTDoIJopvJPEFfC9kdgrtKRR6
emeZZoS3iDk/v01IyKL8L61PLCZ93ZoJ7FNuccnKRGaxP6wEedQarMAuKrmErTJ/fr5SsEs+pSFS
yLJMJ0d7oJtfbcFHLITUwn0H7JrnY0foxKV+VEZjRobKdjTE14nOkp6r58z4yTDjAn+NzRWXZLUa
+MVz1xNAfJi56qRw6xpOoeX5Tg7vpKl2vgUszWrHordHCUY4n9lOvzlAwmymT2wIldkIn+dRyt+Q
lObuRle2F6AMCmQyk2oaMSokLWaGFZWQkTyI803MefKhvYjv2B2wgTpGRZMIlmbGyx0U/uMOkav4
xltRgcDK5UyfNvnRm8sU7hSD/U9SswVf/M/0r/KyaNmdhc4LoJBKSBe6fP5H83tfIhws5X+Os6Hy
5sLsDi8kJtO4el3oVwdKOrhQjA7tCMZxMuQ/97sU3xEJq4s7zZfHDJKeUDTxLYsDvVIgYuRhN/Sm
7AGjtMtstgeqGyguEg+25VwjOOg6Jk8Dq6505VYY8O23lQBhudyZqSLXBqNhmAHDlyfUUFdXfPUB
CWq+2RX0DwSlyoZhQo//KNh/1kpM//Rl/C4zJv5qpLgiEYaZXcewS2mkGa1X4hfcCzxiIK1CCm1U
fVJgEh15NzQhDSR7Y5v2BeIDxDT1AaOh2ogPuysBUOlhbimHLGVRvin6v0z7+uTWBmmZz9jQmmVQ
KccRNjkFsSbgwkj64RRrcdzDT7vi7C5b5v/XrkeIQeK2VM7wBdXTKF0dUuRThCUrX6xzF1s+ZP8w
wehZyuwKfCYI0Y9/MeQwTnd2htUwY8rvraCu59IJXst3ajouer0FCyw1CM9YoEV3snc3GtCJSSLl
wLJPufTXRwSKBlje1ZDEJpcJ8pDaLqRJpfbBkEMcUNbzx+8/YHogsZqPTwz1Lyv4WAKTBLaDW1cV
n1bSsq4vNLkfR0Onh2ZyhFtRdOIJPFCz7p+4OGssl4M3aCyY9cgZ2ChH5NwGUB28qKdmLCST0znT
v9oYHEZtXoQtt2Gk4f3n710nk4Gqykbz0T39t1Nw2zqegk9PPBe6WZmzIbRAp0orD8js3gikPcUl
lM9eMxiqlQfr79l/KnI2sbcbmt4ooNx5C8RSsB0SonXNG08bvPnqQpWrE4YE1DQ4lLW7czD+KwYG
VXSDtoSic5PnJ/TwRjA8yIX5jHjaHGO6JjLad3t7lAcvYCZVUAW1+VXaXBXuiXoMNc45p0mZy5es
UME3HONNMAZrlbtfssDxfWlnnfWHvvd8tMkx5oNSUnK205+FTYbLAoKke7/UP3saE5kcIkklerRX
/RZAUoIBbkz6BbH/LSwdZy81suoFngXUa9kdp6dKHC9rCT5pgToNLk2IvkwxVirXMkafkYNP7qcP
PBP+/bd7F2IbHemoSivbAftV/PNoA5i+jNtFyXoYT8nx1v2VxvxnELZSaEJdTXktzXpj8WLRfEJ5
u913ZHFebmodrXQcL+stMHXRn7W+UIWL7i60ugGsDOZYOLsqoyNEriaB2hoRhFKvyA1qKviAPPr6
OOhnLNZMnghLAXnG1Z32dLPVS4U2hkuTyCyKg9VQ7HMY+3A/8gqn0ryItQkGUFdrAWP8pDofpuyk
2OwGFJ84JAnNsTlkZtRUX509p8sCyNrtuuLox+n/mlD8y58UQT291bcd9WyQ5Mo17Gk6l/FFi/It
NgMW9Ik91Lug/wR1OhcNasiun0opbySDdgOmUeYk1TwGodJPBRYIY2BTporupfeTwa5OTELLhVhZ
zNJN/fg9gRWhYmjd+szRZQOSIxS6M1SVo28nh4SmxJ/wduaMLdf6OOKpauoFqiNgb2HOp4WWrJaP
byQ4ln2QsBP/FWfGuLP4GqZ6J1MsEKmax/dxdQ3x2hEaXnihdfM0ByHCS7Xa66D/mYNmCBGZLbWK
IQ2LZP57CQDvFJcY56walRa7r1LCbs3I7FliG5XBut+LzK3QnxSQYXWwSRhfCZg6XLlPtx7v3pDZ
GNJyPoBltIomrWsoXtWbwsiEX9x6LRan3HaW/l5qPRbeHpq+cVZHFjxRhT6/930a7ex471Ab9eod
Wv2xr1gqcmjDDncDeuQPu8cxxEn6gycXVpQEdfeEGfX1wmLZaEZFVhtX8L06gkBuND3fPURTORlu
j4BNN+RuQZ+nmrBjdK2f7KDlf9E9rL3bYv/6XqiTa28XfSG6aJlbJ92iBWW1W5QZxZi0HqHOVXVE
Sn9nRhah82Oxgtw6Cg3gpiliPF5QiuxlFee0S92DV0IhJzGzlOzS+Ax667bxf2leUZ9RXay0pB4V
hET0fHpWYMTp8bnpTmgx671jP8t8mgeFslUuslsUnzjm3OlGnfOAtCjRl15YYJ4eUNHQZXPyj63T
g5n32BYGlP1UZmTWG9cPlyt2HdkgbLvmBrhShWZxKP6QVouTHW1B7nnEU65zhqFM+MncmGYL5gZP
glWCFH14M+9SNqEgnJn9AQxDWwEnUgqhCmrwJkxUrJnitzi9/yCEn/APf6RRCTWdIQEYLEH3De+y
xX6x7QKdywFzZ92/miphgQvzkttjNPUSZAKTkX/wZ+7HmHy4L86MwfsvkYfPZnp/X9yxbaa2w9y6
1HhHcRHPP+MCMKga7vsPWD0lReBzW6YPu3TzPtDBracoaO8Ez7jDUlDDO1vVTbiY0abGaNbFBkOg
klPs6fKSB9QMOEMB5iGssNm9dg54nBjdewZQ7Fs7lXlrdltqb+C/b1Ol6DgYZPqdU2mp5orFFmkr
AqX/bJGxaZDPcDG+t9McWDo/2Oe/lpdoVz+WW2r39I9tyag2FZPCaMhcYUiHpb3Yc43sJn7YdTXS
+AHoQ6iYl7nhyW/NDQe9IEPv7hdTnx5liB/9dOY/iCNpBvYLkF3mgdbh9zIE8WNpjBvAMfNPHGPR
fkIwP1kMBJX8lMgYsEBipV9SUiTuJYXaV0C2yWSevGJ0B0wPkGXX1u20zQfldc0wv5dTx7Jf4cWv
jPhXxu84C+tUSnLgGaKMxM5DtnQKmk/6zRHOeq3F+NDiwe0yBbG+MvnZGUp7oMOZdBsg8SxTRO44
BVYzNLLlUJJRM//3pkMfVa2oDhgQlzFD43B2mw90wZWJHXxDg0hl3kGh6kQBaEjg6uEZBfU5xRhY
PMl61lQnI0EupNMgKdO6rd67EgnAbiGNuJf671rvCRKqLtfnQBFSNGEOxK658fQ1L2VwZQ0ueTab
Pa/cS8TeNuefJazMRxLQGUcBePGWT5LiJlp/yo3CaQXKNisaH23hRujdQOwMMkC2T+laIw1rZKui
5VxjUG3lRypJ5z0+5PsC8HZ58alzMK4a7uMCY0b7dW+zFqLDDr3bdjPCRIwa0pTRcyawhHdDAMtT
kr2+Zr0EnmS97NeVtDD+DExm+9B4IVt5Bk2PsGvCPWZ5NrzASgzE6pCI/dMbcIXZcTm/AT+k9jxj
lBf39GLi7I9EfRbC1kFg0wji1uPkjwIQhhAEKtjGp7aj7EjLaTh+bGXC6xj5itwV+XqWM73c23eI
4AAa6YQ9dJj3zawUoWvQl5yWNFF9aU8KmLjq8gVOYDIkMIInY72onEDfPNjpG5h3Smc/mKbfT72/
T1Z6bmMQUjaOHzAL74XZDSkPYmIHPy+zkScyxxJrw3lwly5Fs0sFS5tYOKghGTGcDw8dXEhg8HAM
/PSbBEGenzZyEturQ6muqotEy/+jpiqazwfAOowigBGXq7IPN7VzuKOC7SEXQJ5CZTeS5YQMIzeT
0AuT+0QGZF8oOt84n2T6G8xuaXflL6Xi5MpLSdqsTRW+/RBeUMc5kVXf4+s9UnQhXz4osvIoF03p
xkhNpA4C+fX+iwNOhYWVAk7bKoZVXKA333FyYvsLoLrN9j1Vn3JsHizX2o8LcpfIKD5SqwOTqY0G
KOP7He1KepMBxihzea2vvMm4lPpIvjOw23VvU8QYsjfCRV2Dmo902PEDyvnLUsVWt/qg1dGUifRs
fyHb7qSSF/KQDE03k2NuMJ9A5Lh4WZphwgS3P0+8/Y9DAXd56BD+yopwSNpS5Q+pi/Tx3sRRzyI7
5q+t8xE+z2jrpDFOVgI8nAjwiacrITIrxyLuyA+nNociAwqZf0p983F33+xZPF//5iwuwBTXse10
s1lvzLi4kAgZzCa9EKMNLiAw6l9eWSANht8qroMaP50bnsUCiW2+wuN79uc4T6oahGBpn8miiXw3
yExsNEGrszoiuczwe1Y/Or6AS1TVPWpP5AfqxKPjXbY+dEBTCzQ2O68MwQHzl+u8AS01Q2knu+IR
opZgbyW6edJ8wWa5VVwzd/3Bkj2P1iZfdYIhK5yy3nnxLZDoWWtJ/+zoCRVqNYABqtKssA086+HU
8uwJFRvKfhP+9279yipLxpVecUTx84w5ws584EvckoIqZ6FtRONYhiv2IKmjzQgju7jUPZp+nSsM
szXeP2idg+MEZ6R91NL9jNcgLb157DUBhu28xXB24eBSJ0MEy2XJRAqH5/nq3/06sxc0LkJBNLNN
rPWUPEkq6sEZ/f1qKXgYshFCN3cRn7KFrPVqlhEiuLL0jtv3Q3ZR+BoywiHC6yXxKgxe1ruFG7gd
K9gKa4/vx/gNega0MTPkzEkfcz26NxbSvDQFcoyGbm66VmVpZ8zdH1sz8F1BeIOZTENIqoAcgjRC
sWv5a1OMRKoUTvEGRI0oIYBJEg6y4dE+12I0e+tBVu3R+geym0UpiFfFTtq0rf2fJjgDwQTHn42A
mEp0lDniTTtbBW+nLIItF3MKwSrfbjJHKpm4rAczWv2RiwK8aAXJksjZcwoNtNiC82HiFbPJKv26
02Qp1xEOObDOh0+ujlFwN7TUXK97HSFJ+D3FY8xK/dXUZZaOuEsxsV6FNAGr9Wo2tF3UEfL9JytY
zaihXhJjZAxY44BGIFEdJ4J/4REZh1s9jb9CS/6t80pLslLJK2HGIFl3M5ejh4UW4lEqY5aAisMG
TkDBqsqW8jow9bzG35em2+IAvAthP9j+TVJG1X8U2FQYm4zH6+3W6vIBykJmjqBXuW8J9CmF4qda
pOyw8wDIZZk07JWEGa0ZQHOHLByurvuTVKWbzr85cjvwGUREpBl6Jxv191a04/91p5L+V63nZgWU
DBojzkYWmDmqSe7daIysK0UyCLVqv6JTfPxtmbj6JF8aSyDQvgFX8P8OHBcXK0eSP255hkmwXUHm
sXFjtZlLoYkreLLFGf+co2q0gRG3CQHiS6C4g1H7jGFV38wKUrI50ReWUriJ9SPkM5/L9gOF/KA6
RAM8IcAndhpIubxZ5LlzqdvjvibF99vmtJuHKwl0rz3ewlfNB/wZhKZHSc+IrD9RObLME7kjuU/j
OfKaXa0QDWCKQ9NmRUC3o/qxbqAHZ4JbMLPqMxqr6aPtIHS4uxD6Y3WSG9CAdQqy6SOmJKq+as2a
/6uWRhtENEHwew+Vlq0hSAPR356wb9x7wN3HECMoSGImR0dvRr0/A42O8lSTI7oVDbpmVLlhJuq1
IDrUfIas3/F4xurBf8r9mTa52euabATjb6hy14lGFinS1A1oIjiDR0fu2QhtJ98W4jvdC2/z6/0i
w5aADI2kr5qC9JFpuUvOjVF0xjf/r0Y9IzIrLZ+ZI0CkQyPvUzNweR2GpAUl2iW79mP49eI9snnQ
+sDCC8Rh3LhKq7SxtGnvakcTUCpLHds164i6rmNmOi2Is7l5m/QBNk/Oi3AvSIBGrGFQS7YUxdhw
2Qcq+0GC6n8DYsbqJ7QGn5vPIJXiPMCo9AmjBasM3e7jY/0ArgC+GNBti8d1NwjI74lIWRrosU95
zJqr6KoxzlTJZEcznw6JDvX6MqkxLxNm7hLu8Jx2DHv1rXQzkqjoMHjm5pmwxZPylu+xkGxOLI04
7TwFCJHyJYPRRyiizT1D570MllJrO3VM9eu1k9GI1rzOrrLAVK0jXxkFkId1si8LIIu0HPbTLf6A
Qk2h32/MZdcP3SaccvQCCDJTbEo7H8VszZdmf99rRUesKcQhapyqgOFIMObVQHAsaykDB81cj4+P
hheUaiWKt09g5gtsUDKKNmgw1sxuhpfjdA2TgUJmgg2ZFfwGZNhMM/8LUR5q8DaeOdYb7hrJiWW2
+xO2q1Y0Wz8S/HhSWR3uor3TENwUD4dD07c9cF2j0EE0WPHD1B4K5jV5/fQb/1BAlmG5hVpi/4eQ
0vHNG5m94oSb6y8cbzChpBwnXZQI5kbaRXE7gE/fkZe7mXGd3fspHKhoH+B9UQ/77aqfdCW1tQKi
rwiNvm/iKyozvb1hKXYOwfE53Uw/Ra6viKbcjIXHnww1/DQWHB4JS4ew1tl3xSwRajZKLa2pTVui
CrlywG3QjRaSStiLnbrwErGFrXU/ygizRshgNiZI7TCvzW2xL9Fg9V0+vd3c4VybWEWiw/G+tN48
RNpPogzlw6ZUqYWWwnyASS+zVq5xgFIR2KT7o+V79DBOwJUEGdIVvLmHzD1+mER6a887XyE3JEro
ppg1vTSzeUcgjh1IkXK46Si0tgxwraV+z4/8uhtTBFRzeMY9cRn6XADeXGlhYe2SGgZyTCL177Zt
BzkAmEsJn8rOG5NDVSM025RYoREed3HtOoJfEgqwDxHZhdN2fw0p+jHyn6lp1FEo5z5UnAUR16rh
eDYD0hWg8UQShHGitfUPbU3zUmgIuVe9x7pj0hS2GPCMGg3v4xZNuZFeRI+2IDW3Vo5h3/MOir4v
2tpqjgiLwHCPZPxHENzieDZ4rEA2UBbnOlXPKA4eUDu/LRgtrwzj+mKun1zE0+cwsxUcMnwowxVs
/2brSz3ntsAEOx6+/i9Jr048G8FWnsZDBPRl8qy4hHXppWrswrUZOwnUziQsxwpbnOSvrhCO2JNA
xe3AFfeOX2FkmneE/fBeuQi1tCQvocnTdET6yD/L9rIbL1HJ3YhrpVD70MXbu40jwrpsiMDqi/Vn
3/cwyMa3exs1C/bSRMwQ/QupbKLvTq7khTKmQdxsmv2qVokGVO+RmW4s60YC9LNvUDeV6iWdknTw
rrFbU2UuLM1JWC3e2QEY/Cp98vDF79EDNiMp2KuNr5hQlji/cfrDRa2geBTlK2r4iCgKS/eaIZye
Lwmwl9la5Xf12MpI3UIcy9tkKTXyM3+FcSkfi6hT0BGI+e4VAXrNGZFdfkhHdiyTrLNnN8Nu09Ns
uC4h6MVrRmej8dE6f2RSKvdtRLCSDjVbBj2M22zJ/ALqclnoksiieIBZDcNaNkTMJAyEy9yi0S7k
tr57x6TnoPGeKhz3EoeKVmaFPP4CIV3/lmNA9msbxFfiBLMdMIwIJb6JolWIzzjEDWT9x3ygmmRh
PLm259S1zSTpjyNBPlguHn9FMf+NJajQLYVRZq+mI/5YTm4Pz7EjuMBbCJ/4/f21nKXqV7gY2fM4
sDcLFst7sLHrRyKnbvvCYeqjKw4h0MsKR4PHjss/TnaDu1/NDHTxP7STDSpAsVFC6esvcHb+5Hd0
VSKOH3dMZ+DG7i1h8Lyp011HNky1PfPj5NKeqO5FBDu2EsRi7rozIkUO2M/BLNxaK9aVyXlmu7qK
bkvsyK6Rhw9rNl1B+gSBzKmW06/vz5ysamXq2lcG380ub3H0S/+eEVH2F7V5XJkq83OucxiOrU42
WswKYbSsbD8I9oYDzQ5epzkQbUE0kIRhqx4k8jJYv34TSEaCZ0/XWoE4htvMQsMyueMPUHC2dlXt
NNf6Krkzzt+/TuIh88w1scSoS14giuS4lVvMfzk3ynyt3JcEgejfOC9ndbC5RLcUSWRXb6uJQbIm
TXLWfrZ+8+YlCv1lXVTJEzi7tez1FKP6GjswUZ7y2wtsU217dK0sqCr6e3PSxPRKfVHa07i62UYQ
6EXjM8/RFi55j/g536V1//F24EC3veSmTZIh1fIqyfZce6Q6yzsdPPtaFFTQBvahWwFvcgtvGI9d
Cu+EQ8guhCvfMHSd/eCeptWQddEsNpkvAc01kAvEbs7YWgkva3ttq3MCrQVAXZ358vGfmLDBZXjo
XJbC4l6j6tTK5UDEhSd7WXvpvJCqQPKDn/g477l6YOZf68n6rLyKKTcEVs3oiV3HkhTx8qPvyI0Z
yn+BSzXgpiSxoAREaNe5cyNLQvHNYW2gZaD9x1T0BMF/ZlDEG3Cu4RF0muNnFnmuN0cSjWFqhp00
zVqijgZkbKqlG+ak4+xKbovnrjfJf1Q/mFcAlOiuF5j13WEDA/1z7XfPoJ9+vfjs+JVXR5Fijbi6
j3MNesKoYB0eZliRUifDytZTPduc8PBmj3sLPG0gTDO2pos8kWJqjsdjrm7zBkTDxzmeBsQxsD9c
DyK/m1XURNLZApGNAZ6yLdQ7WgWDPh+L5Js2M3ipb6xaK6ZDr+u4PmAZnxh9o8SOdQ+ncdZB3xSI
pf7XDHocQLuAaIdUxWUwTIG4UfSvnfAtQCfzpPwOUHx+vPxUwbJ/+wq2Qa4cbhDQwgaApZtvHMMv
J6O/HTsAaiFlMMtNDyWEnQytSD+H/ULsEExZVBpqJD8eAl8fawS/Sn/dWb74kgVdVdWS/ECDAyjA
KreH+AHYrx+Dj7+iOtIeNF3M5Dw+eAfZH8GXixcL4mFCgvvUE1VV1H8FPYvwuQqLfVGFwvRwwgbi
iDtc6iUWhs2DqOTXmhGYzDwSw3MNw37+TGUF9dTrf6gfUVaLbofhRKIO8NSrzB3H9VQ0qcrg9WFC
3pi7ech5mqVUfLcId741xcIytKubhMieC1cTTgQru5hLvruIWJqKNCSJBGcXnczsSE8JXmO75AVY
Ocdnsve/ZE2QL3KOJcSIvMerKRauibSNqX8q4wb3fTJpSVM0xNTKW4AWWVD6VgoQnbfC6uOncr1v
2b+0umArohi7y1nLgCCSxnNewL3HsGdWFCTM9JRwj0cPr3+MESGdhI1ZA9cz/NyPcBrtDxcguU/W
b81ZQzL1c67ZRt5EIsTF4gBI8KgQWNhBlgvv5W4ndqq/AAZc7c9vfmyHNEXYd9PUF3aldm70jccv
m4ivvusYgdFNLJLK86c22EFV/WxeRKPtmpuh/ShBW7wylUE1oGIOCEN2v5nZ6wxazIcq5Wyeaco4
VZzVf44Sw2jB2/5DhPdGbfKJbHfvfaLenRNk1uPjlGXyw8z7PTDypUW9KI9DY24RGJ8v2H956/Wr
JN+0Q27m3pUoAdHC0bdwo/ClJtwyYZcHoKwBfWUVW2afnQYUG6qe8S2umjTP7TPEaQwoJVZz55y+
Q2MP3IZkaAbix0Cvn2Mb2VuQ7Vh/i0e20RCwxpWX0yXgtI6yBfR88eqa1w7dAcmQAGsR2sbCGpKu
OHZYuK+WVXPWx4uaXnWIEn88AtI6CXcS0J6ufmifj1Ql/GlQUwM6ov4vwC0vrOpB6x6gnpG6Hapn
RXl0NwDemc/PGdA9TU2mm3TSmSmiEWhttpu2kB9c5lwMO68IqFWsPj6ECtmU+8k1yKWGlrv0mbYi
O6n0Jzn/NtuW6CdbFHGdUNMDf+40RCfNyZwV27SLpr513E0i4Xd93Ew+YQUbYmxjVxWmoPTxx2C9
5qeuq5Lh6ikZO0wTTaDx/sJwQ9fgTt4/5wubD/MsnkJ6HYs89YtgBCgdodoLZtpE4QhaXTPeKr7a
NbQL0kwOo6xps3hYTRnMxV5QfWqD1Z1ZGumxLXWBdgQ3ejRV2oumjOKsStOMkWQv7avozGQYKvEs
cHrLBIbn8nWra4UW1y958Uc669PREIRwr4YPCqRxf6PNDjKaBFokiwc3r3vob7j/P37eqsCwfck/
BN2D5xkxW0qPuYi9DiHuMQRHTdvI3rv2SmWc0r3pOLPrC4M4n3ovYle/K6RyH5LKJa7hJZIhFdAe
UUSCOSFqkOc9w5zsKan5doz8qfD2lr6I0a0oGgKfl2s9O/yHCazOgjC4jUZe1P0CjOASmwgDZmx+
8APRnsqxIamHJpDU25Bz99prtJUqsDJBq5ArIcjffhi2iInlmhy+b5h4aVSZHPakHE1crRR0QCTl
k/eKRD+qkjaLKAa8p7sv6WJF+jwz7sAsAD14sRNE1UngIkebCPW6gBuPeOyfwm4wrkPjSNc2JHZH
aAs6UCxdYx89BHcuRUy/qaCh0g3ynoNbOWQSJg6tHk8mhrJCYue3WsDXwi0S7dXHU2eQ3TNRYqP7
Olby0FL88/P7HgqcOfy6S53C3QdOKkHKlmMbwDuOMF1cexv/ghZbBWnAwSMYF2UoE5U6581OS/sI
8MwQ9RtBAfUlPZFwKjRtw0PcY7j94kRDN9iR3+HH5WL4iHPE7VM2tdZaan9SoISFaxOJm28pGAkb
zKADcrUlh9wCZ//j0AXk+VQE8ul0zWgkYquS9lIi7yDB+ha9wtkd3R1VgcBITo/VTsuyO3iQyI29
TFZfOrOzQLqoiImspFxOEHEfmpgkSEE9dbgQuwGCsSqnrLW3zK2l1IawT1JA5aBZUjwjD5foOcii
UkeiZWFZxDMHKKiXxQQK0Nk1EU2e62e7pM2m1PZpGn/keT5w/iAM/ERoVZG13fmYUig/ojzrkSSS
u3J6QFQ7lD5vgKMxtazoGTZ1NlKgDmR+p8ef/toNm5TonWWg/usD68j7i+WOO5IxlfWqfSzHANUn
hOqq9EwAtF+ofcGJTto3F0Qli+PueemCtyfH16Czw/r8KFmoaKtr20MMnJ8UwgEY13Dnp54eeida
pNhMpPwLIVErAR0YQUrUvYI7ZOdXb85dV/ZDppU+f6Y4Ju0woNUZTsYLXVQ18kMJxJGKgcxIAKd3
ifpz0sXx2LzAh9vsTYJipCD/DVZKNRDpy6c+HdFhIv2sK+958ieXtLO71RZ7a1Kq4WPACgGVWw43
keRZyl8p2+At0eq3GlVnuuCoAuBezBSQETPafiz5T2evj/b6BE+7IatcQM+onp/5NAvu8hVFJhJ9
6WaaCquCM0WmL4Nxss8p7jBIiWTmo6hCU2UwGduQnDCBcpQcQ0zYJf6ZULc/quj5/ZCpvoTEuhgR
PGL30LxG7VPwg6wStwsnVpIXHhUr83qQuDOyW/CRYhlUiXwPnQc+Exg4C+s5oGWcWayI+xz8NDES
J+MTZFK9eUfdF8RiTpk5QrfeCi3f8obo9kh38GSjhohJfUCQvmhYuf0fWluIfdX/LiRHGhWZLZ5i
HqfAilqd2Mo1NUzje8xe2x0zfakf+fKvTfpgPEhfzMxtD/phRveoETsGR+NVpDp1OeSVjoL29FQQ
UNFIlQkTqxdDfs9qHgPb0K+u/2DzMN3kKkMxObQAR9r8sfPjibCAEhHsr3JqwUXe/4Nf0JLHTWmn
zKHZau0USpX6O0IEA01UJHdP/FMmo6eoTF4t9S4eeQ1nM3EpKuoPV0ExvcogLsnuAU1XkRwEJdM7
Jza5WO2ZtVOWM6BLEcMKSX6OhtCMxNG4qUieWc74qxWe3k1ixu5gYvQrypnoJhQF6SGWUrT6e2Re
B1Cs2dKMBzF7oDMOcIpjXZRPUKrN5Lw+0D5VseHkN0JZBoOc+G4zeb41ZOTlxJTReLSWgjPQ3Rqh
GfsKPpgtVWkxygnARMEeqNvSMmw9/16BF02JjTK8R1MhSyRlU8AyzKv9+ga41xm7TghCzw2fFkJL
ZD7z4VtogRsV3fNJKoFj1HKIGJ2dLlI2arzYH7L3Zl9rf57lUQDkIhiNDdYAS3yC2hzTaCWbgzp8
b61Tr7Wi9efaopvUmaHm6IS55xZB/RYdwHi3WYYK9dp77hyK8cDwFPYD/3M+rNDuCEPkaUeZSKyc
Uk37jYrzCszz9Fd6Gjl35GvCEMJopFsw7GnsCfMvZt8lqhsUKWz27ifkvPBnYktAnLho0Gs3oLqg
SME4ceEwB8ZFIvj0j28QkgIDxv3+1tmezSshXtlNjSdLpA+DyUPVlqqDgBNJsyESYh53ywYZg9RP
paYyv9NYbdQawF/bt52ld9KqbYtTwCRW4tkILFU1ou1RWu5s2oX29GeCVJTqW7O+jDx2calmYJ+I
J/grUS9QiFIyc10GkQHrkRaXjxbOmoe44MMBmz8BaOsSUO9iwU/AqgCcFpFk0en478XT07tiJPRD
w0v4PFXOZBrb5zwauzXvgdbpag6oF77pxAyACCHvKqtBOfkZrjOTps0E9QmbfUOeGu0aUjgTwxZC
Sf6nfoUlsXwKnNe+a7qVtD7Oogynt2UA5l9XE+XkVTgwumW2d4X9o7Bu6ybgJUPmdevi+eJ7iKyv
dWzuOgaxLBmAMV3WawW+X3wbFWRtt3gqISwkLg65ep7dexzr98/uHnmBsQ90qXgAiGWbtqWUKMzF
vbFzNgufUC56l+LDIkWPuWUSBOK/2P7YvXDOFLjD2t13kUsMukSueSp3zDWL+O7IBbgWrv0R0m+m
iB/fwSixvmQQkKdlLG3qd3Gm60XoCoXj+zufRUS0iOBdCvK8XiWTZSNLYOxli6h45wf71C9nzdrl
Ttesm/1Pd3KPMVz7HwRfZyn8Ub5dzU/V07mdOkGH8ExY8kCG+AATfM47ecba2ouIER5Ygwc8ryeA
78SjsJrL7RuOZZ3in4lqQ6aFSLn5dyOCK9l9uyG91azHUDM2nfuTu8gZJDepN6BHBegT2gYNo+T5
hkktHiehIIPF+giQ+tg+t8njISgTgcT3xTNH/AMjLLTDufv44mzdNdxR88qwDxiBLXVdNb+gGWAV
ba1N91GPrjrOIsg7FSa1Gss4142lFKA7XddUbkQGrOC83cXRGh/qPk9xYgHZyqVcRAD8wJAfJLCu
d5UzQ7Q3CClwqh3WnYdxdJSLGVnEqobdsfjw6Y+uATsPKTJnpEmBUcA/3PA9BInsqrk00yOglTba
K/fQ6m3RbIux5lTetLGhLadMJLLSATmxq8lR3FsXNKzN5hSZNk+dIMqUqVJrIJWPR1NNfaPbLjuK
JOMWdYWyZ/LWUOD+JC2MzPH2KyDlUTb3GGRhHDC/R2hDAm04ncu9+c8i03/zsW6txxzBjBAxXjVN
sDKEGlf6ssQPxtT5VW8d+VHMCyKEULHDzG1aReyk4aBct0CkKRFZrkSH49otauZZZX+4+vjOixCN
caDLM8jO6Ov+fwasqZaQm6NucAULwkenU4zumgw/TL8fysZ+CMeVcjdYbz/84WEnYHYZqnDcyhBq
kGOzeng7An8CFs5JOLMH9MMr5vF0Rz5zTNsBiG7y8pEuzRLU391RgLIFz84r4e21r5Jfbi/OKEUB
9tu/MxTwkSrayKx23rrgox0bT73bN1KsZ4miIC53RodC0jcfuvR3su0kosnCuMYIrVb8gnw/SmKH
ICpqseX5oDB7jB/zimIaTEOlRi6bfz+AP8bE9L5bEquWZpumm9Tzl1SB7bVEQOSj8FKHLHm+8xQY
87LIf9GMT0CB80Y003kbt7M1OooltO3j94XlGFpuB9jWjNe1Jmap86dbNVDZEJv7dWx/rRMJIWwm
2KfMGcsGFUFYzOIhFnW68JNWdE2T8q2iYLfidbHEQfmGD3YuxzysHoYGzTDj7reYncWMgY20dD4F
oHQVpKZgQ8FG5pXrT2PahRu+/lgMNYVwm05tCOMk6uH8xSsXXIECjcEeaBdZXW+UtS/7qL+yv5WO
0dAdF36UjEnzPdC8PrglWzokryetqK5iUYC4qAPRyYo4bz5VliFctKRBVcFoWxr9NcTZBU/uGmHW
jDuPA2TybR7vKlU2fEEzE3MlEqnzVFICYCSOf+ii3+W8mI4G0qeAWErWhIe6bkqI3XOAnWD05jdd
0hCWgacezNzDxJz5R4oLC0vrOjr20mv2wE8BRHuXg4F7UeS4uhARIn0xibOeE0X1QSeqZFIPI0M8
705XamKu9aofqU8ezbB79U2yd0HnkFvkSSpoQZS/ZKwKkEJW31qev73QnQoBDo7ezYR64A7zHXqS
V1l4KBlU2m6hZIv88xqwvb8G40lGa5v4yD7ts0zBQKLozp7Qy58bbf/aoES7yBha25qWFPTzY1Kr
EkHHDFQF2sEau6JDhwJej7vYFJY79DeoVIi1i1H6SizOhbdOgHASSDYmHOFtdOsb40HFyt4eUzzC
txPkRh3qnd5GOOTgN/m7SGNk/zICSNGX3llsWELqzLM+1jkh1IPFUJgMfvYEzqmR5UDaeQ1i121Q
Xa+U7Yaj4Gk2Q9SMk3nVVjaZtAoJXDuAbfnYLyhXl25cL2YJhI3OwmX5xbkHrat0IzFrFtJqZcFX
iwKJkUBirvOxf0nRr38ym3cjqpvRSmh/i0IxZHO/r7pNXNcF4oMrDcWnRTHjAnn5QTitOEsQK+vc
47+EDVMB+MAYzxUz28WXkzRQnAltqUjLWbhYtUpa1dABReL+vMCPNtzl+j1Ugh4kQ3us4oa75NP8
1zW6Hbg1O2fi+CTlb9/HdFeg4D8tJYf48JwZwXYhmH4nVPt/08Uu8YdjAfZP48IdwKjm7+hZHqfk
AMIvrNR3zgQA9lJCud4ILsHnnndtLDu5ScHBtYOL9ZPD9V0z4O3+gtPHN5PO8cyu8mYUb8liXfpM
+qFJmR62Lb/l/MNXfN9oFGF0ogm9bjhYyaZcLld47xqnnJbb0Yv0B36gi+U/tMQuiamHfYSOVAvX
0zb1P5mx6NUSLU237afZ9hunOW+5zh23EhnVwQuB/j9rIR6DE5YNiIh5euShBZWF7njO1VsDcgsh
QR9hTIkpLHMk9Q/yvqaWC6uMp2i9f4AoqP0ze95Yg9S2TRpAol0I9535mENCESEKieRE4rNBHpjo
x3v4SL01Ke1VA5AQ7hTffmskwWhg1tfjGDiuoQB91PkUCYiLmhOvkrRawHORXymGtfyQAzCaEpiT
EV8bOxPFggiSY+H3ZT5CBZJDlpWzcSg09dlrD99nPY0JV5uILB69ORjKCdDJm/gqwZAd31XcKHkJ
//2FncUslV7qg5zMIPl25NQ5L1TKa2DqSlX1CIHf5f9GkIoyK0f8JAcHZUDHkH9TcNtLQ9UNScob
27lOQgon42LZ4NYLvM30Io29kEI3ykdRdGP5TvYaLZO7r8AhaRB452CWCQH2xGAOuYL7enn8vqlO
xeJ2KT5X0bVH8VpPKxBMLvjmH11rYwI7x2znMI9SiZWdSYfnJdkyglA/asybDOo9VFdwDlgtl6uj
IsWnqXRU2TQdulxNf7H0ptgt7zH0ADM2EhZkDSxzAiYkRo0sSGzhJcut4DpzGo3TNuS0o+5monXV
dkTJ5kQm4+j1hw/NYlG+kHs+mFV9vQVyAuxrYt2KooMDzr7AvMlj1Joz5Oc77TK32gV3BBlTUybE
qbRQxuww5uh2i6522lfgoe155BOSOT7jVN/XEerVTmYjUlN6WOOEup4CX0NpjyTH8kW/5aFYNoLB
HiRfwVDQaQMnh7OY1VN+xJH+I4ZBqh8u4kBNS4rVjCk3ZcbCkW9K3z/Ks9J2mS3deyz3i4XdPnki
MR2rs8+rSPUWWJnug4AH1G1PZatOXwGIPgoFTk0GzVwPSbU0cZsQwupQqm1hv3v+Zy9QATX7Ztqz
p2lTByqU+OJ/EruAvTJ4rxzuPqbvjEGOmwgfCLNzfINRa3hqIFQiek6f++ubvLRv7bM/KuT6p/ck
N/C4bFLvegD96eO+0LyRS305o9qxn+khv/9x1mSN/BWDqWB67jfSTANs35bLyNjIgScQB6V5IBbt
fnt0EYsyIFO9h8Z4d9Fdzeqv2mtOJ8avUSG16MINFRse3iWL+6X0r/wtFKla5LMaPLvXPn5MYHrb
VqPf6J3q5SndmzWOmtP4jlrnjjPdwUejDvpn/1+1vWR8SHgZroPUcbfM0ANXoVtzojBYiV0YOvvP
sP+91fZ3PFVZjVQYSKJJ7cpEml/qGNDGjkAY6rsbniB+Xjdx7Qm0ve3pat6OdwLavOIl+jSzbW80
ANBU8eZJ4Tjk9Whm7JZH5Ta/sGdcqdvc0aYhTe2L1Xf1rWquCtGqMi14SYj3ILXF0r+LqvIGaki5
cd0gMNb+GXBZ8T+wXsmkZ17rt6/L8YnbWL4jdfCBLy6XmInICyKideNFcUxyIHhpJkPNKqNHE+FO
ppmO7AhpGqfXAO0o3g7YzXCTN2s32wbeCqtntZGB//wP+xUIj6XD31TXlYsPGGAAuUV77RqWNBrR
fGxs7tdWbRcPm6/XZN7ljj7jji89UNT+wJASfAM78i0XqufeoWxETAu8eKSyv7+HIMz2IduCH9UA
Keg/vSCLp17jHpQgLqFXJc60HHCVYu+csVj1QEgKP0AwLmmr9oJVuoExY3g97LIwNlrHoQjoAntM
7v9AQ3yYCfHE9XBtna36c26S4qoeG+9a/FZD0Oe5Cr8cbdCUCJAz2vAld2/6vF+toTfDwFdwnpRS
3WKY7Sd07pByXxO0DBblErAPllU1oUkaDVZhTZmWYQCWvdSEJO6NY92fRAbEn00p4vj10EIjTMCU
CQQmgvi2W4s+QdLC30UAtYnsj3d+XTdrPbqrVdKF3N1hLEf8UgffxP5ZEVwr38YDZzla45/j7FCq
lSaK+0UsakO89MnrSD3srL1JZjko316H8Z3cjrLGzQI1PYgFnD+42RuGlTvGltNs9uKwAiZ+E6A1
FMyclkGHR9sW1+Zhs2aK/tqPwMgG3l7OHUPjPD6xd4T8qODJ8qWQbemQ0pgGj/0H2iKSdca1ooG3
CovInP1RSkLHsATKqu75c8CODwHu6CH7e4OTqNUZoNSQB+FnXyyYBBgCehgq9MEWf3gmahzLOL2c
ZK6SPB1+bt2JfbQFAAuXALsVOJUjIYXAJgFAySVcTQtZDAhg1/WMW3mp43TJ+Qh6jA9m3Ug63Dx8
FCFm/tTb2tQdYaWPfiDHVKl3WfvMVOTNbfvtcaH0p7pwY7rHgqa/N25LNryl/R/Dn+FTeGDkwC/S
+ZTID7h9AnFUOqrcW69kO4sJTae0Ariv0+8cHjkc5p7OfJvsf3aSAXHN+joV1We4XlNVKPZIA+rr
g8s6d5RGz1zwAz0Z/KZcQOxsWOmtL8+yYkfO7XiMnSHVw6w8rBl4P+J6OpmTVl9jhWo4PKTYr4kn
hQQA0mgtgG/OkCf7WNXDtIhMMPElEoNPKzWY7c/gMHprjgu5Py2F+dtKUIz4sHjDTEKpxkr+TQJf
8K47w5rXJh4macdGVP8SbA3jIOC6AuPlI69jDhRrHhmMcv9zzwcU+1st7YIUcq3Zn/tAjDIMvmWH
c4C+Hhzs05PgbFjUOHg+jMYXRyUpeRW4Sy7UXDGPhU9hhlofDCnnTlHjy/tm/qHLlh6L0r8eCCwS
8/L8M52KLo0pCPQtfD2n2uHSf9x9W/rr6iNd5aNh8pNQkf8ivBQIBQKgJCaSRWhr3KpP9rdRGtfg
UN4K4nG8hRlYmoEhoXlevPaSsbWMlwGD4UHrpAD5DM3yfh18dEwIqy+cSVm5+beEKT+QWFgGxlG9
H8j7rT7lPTF8invdg0SNHJ9fgBuTCc4gHsXMNDmUp08EcWsUdmBambuMH7P+AVhP71VR0j6Ez0VQ
oOHIPcoj6sQLc4AahCD3iVqb5knvsaY+b89WkVvcBCaRnXMdiUN2rJhlxlrwrnPK+1nngVi4OAQU
596T8OSNgmEnGlG07im9zVjL4+7LZdxLnEQUQJUhDgNsDFdiGZp+s4LLwzkhSlXcRe0HeA2IP1qw
UjyCM2Q7UQzMU3MiQ+HCe2F2L5Qtbqf5qYgbYnB3lFWlXHp6AvRxMrfpCIZJ05/CEZJMhxKf4ek7
cPvzYTlt7yHWYIRRQ4jarIk24eBOGt8mNB2Tn8Z8T+TUtqQ2m6pLFxpv0wMuX91h7+xTwcXLnPfu
/YJ3uGp7eGStiuPgcDsoUv9GlXt0cwuUVu8pmyr567YC0qW978fYKzfQOkabv3iiCyr6UmLVOW45
9ytO+Ljm7RJ6e4DfBADeizgdgll++v1tZFs2q1/tE8+xJEDix1MCs0D/+fOvyOZiWaip/mEKq9mk
qWNio1rq0tx27MrmO64b5L1Lu7J5atNsjtLhe/HyIx9ulpSMuS2wZYcBlnRzQEU/GBaT/nXjsfA+
YUCvra1LGf5MzO6kBod6MyuqplOeEbeKkYr7+KoT1IGPM2q6sk1uHcZTMc11N5xN8Qlxw/o9cXUD
WnC6a/wYdTs6dbNEmmHajqVLxp0UiMfT1yRwxgBI0i93GkDtpmukJHhfUDYZHjJL2tc8d6KRHN3i
JLhZGEnBk7Duw/7sjPAyYj/ADXMvH6kPL6DM4t/SSS/7NKL/roOuaJLAo16MbQ5aB3JULHARiDz1
dhHUwvESFJh8Ij5V8tV87K9wwyFFo6lyQbKScG4vGR9sJWrxUC6P0LEt/OfQCOTQPKzHpM3MBFa3
aqORLS5ejX/tSTEtPuSboWD3QKhAgAnJu78J+5uc7d0ByiovCtJicq4IcnejdfaHF0X2na3htyO5
RNJF61G8Fmf/Gi704/u45ijQ6UNpZGp11M+MUSGRB3XB/2iXPKWcwOOGhJl25lfM6bOL4CAQxFyH
Rt/J3wxzGy2mgRZLsreN1grngA7GpsbplnVDZxm+Ro8hLsCAU69S8qQhRsg5c8VYGKgaKUDQrFCk
a4DMfwzh9y40binKjnBdgoy9RkPEgLlCSCn6EHWfnERQ6uiiPkLP/kllwbOAWp94wy9HFtRk2hr8
qkoYe73o0ASp5WZAy10hjo3XdmW5qxegDBJp7XhhkT8mQix5FgjnXeVBq3OP1wBlyP/7M7VFRq61
SQ5UqYSKBm1kp0PdgDyBJ0ywEdJ94+Ots7zUyXMZVSNtye18pSQUM8W8yicOwmQXvIIY7hWQjcYO
RQa0fsHV682fWuMxRf3zyKDaUVqbfGxz+/5kvhEff190XvXmYvGLuJCEWEkDQw0B7mm7fqHH4gsC
4iq/S7wxrvd25i1WBU3muH2QaIMhfrm295J58k2gt4NXFdUEvJdDNW2aH8O8a+ULDE3XCymVrQWi
Tx74D5T7MA6bcntKfLZNM87gUOPJX/QIXSRsb5xW+O0A2dK3NxRZHlNCoT62ts8fjxcHI4WDR2Co
ikTbCtSMz+SrbeFZlu4J5HEcVjL1BleRC7rIjJAPDvYywAyc4U+JRQF9cIw8iRL7Qvv6FXvELhdc
OYY4eotRRnoC50N5KfRRQ9dmzb/zqoT2z2FpxwmIy2iFZIlzMBZTsTj0nf0mNF+/3Mg2Vhp3uMqm
8M2RN1Dgsp69Npmiy1RBp7AEBcbVGXAF9R9rlT77SAmmzV41V2wXiYHfnQQzYbuDLD/aBWegav93
sy8XV8MNCOlTHzWHFtAIq7xe1eJI3NslDGj7wJkgeGrsbNKhtMdLtYXcz5VfOLKElJaqBZP/fKxs
ZExbytrS/RUpFZTJaYEfH7gQxsnl4EPCs/pi0kM4faR9rrZLjyEsjuHRBY4YjIrW7MwlJYLntKAW
L/GB0Yd/Md+T5Vc9N5iQBOuxCTmUmUREcrrxW3Nfgb51MurlZ4PvYJlJ/qdAz26nSveeuRERD890
MmLpY7k8Drg0pC/iYxiTNz79OZNmz/arCv01DVbt0yZ0UnYrW5fKb+uo6lKDFLwQyK4ghcsSTo4L
k3FuTHBEygSkCq7CpGED4EirM48Kpd9sIrPRn1yBZV57E9MZhuQR70ikFmY86vhm1WbKkMI3vn7C
HEUsml1QzvQJXgzvKzkSp8UQnQkCwNOFheK8dlOicdrGE85RvVuYjHNk7zfFEy4RCvTWCKzQ4uZx
mNZyvpk1Mp7VjyenlSOj6FicOpvEsq2cu1mkJwGb1BVNbuiGUPImIdrIE5q/1ZcksxP7gXrhl9iv
3T5gSaDCarJyL+2K/GqXUV1RtwnoJNJh6zJwLslgSqnmtXvj1wZ08dgteR+SpbbkgkwTXDWF/goT
1uqNZ0+2kCEYh4ENWL8rPuuF/d1rWvp5HcTDlyQCvHvjv1/lKtfRoSVhJJVuAa7gGGKfTZe0KehW
geNrGJdtJc4Bocey79R/54GaoUUmjSIKdpA2Fm204T+PSzhROVJj7gYwF+Krt6F3BU/2s1bTcdGO
Fu6BMUwXSyJ3nxMcaSSGBw40MNlL243Ser7v3lHs2VSbC2iUSr6V/E6OaPEVxVxoGCXy/kXWVsAz
dgLTQszHKNJsTTxO+SlpRmsl+a0Jqh99UCQJfGMB48H4O8SDfwe8cWnMg8Tx353mv2C8vJdDx4O+
16cossDk0q4k0YxIODlmI8y90lMEasEAxojnaxB7H2zMgE0d1fpv7pft6OLk3FGg5Mci3jtNGtXv
N+Q5luWRzpTJQQ6ERaAGxjc0jIcV303xiHXpvYYbf7od4Wf2jJMnOsfpjJ/z8q6IqVhdwYtEva96
6MxKYIcEuuIQLftMlzPmTdxCIGSGGM0T88IoJIZPWQzhwfcMkZFNZuT5pGjG7gARb5nmuXT7njIN
fo2HWo+lLxFqScXR4sbmajyNMeWSPXU9/jHMUy+TT4+uKZ0k6OF+EyQlxBE/KyxmDrvZLb5XpoZy
9qHHMaruepfQWuoi35sr9tEClXLL3M1aNHrIaJj/atweIrGf8icK8BnujoLpnwhshh1F0l2IdANC
YLWPgN3S/20SMIExSWRhj3cwEp+E3fzqrJYata27KJ8PeEHOcRRpzqzFBQcpcIpCCUu0RqYwfsbp
8LvXb6qoE5aXPwH8tqmyckXREm3GBHauLT3d9bDLhjw1WnQEegPIgyO9bo/ujV+DWoCvadfEN8fQ
8VfhahhyIoPPsqjC7javapJIuMfoeK/rrepjmeBPY/tlgM/r+ZO03jxI6DqF2g8GSqn8bjwDec2M
65/vdOZsvS/qjhZZT0cu05qHte65LspYZlHH1PPPoX3WTCh1qpqixyjgB0ApCUZTsXkGjOiI/COt
B/7nTvn1+oI5AiJwR1kF7pOq3xwmm1KOafZ0Cvel2p1/qChvA4hmRM8zO5dXARdepy+stslPhkoI
sm/uWN2nwGnD+KaQm/xfdo5DByqtOWcLSA3f1bXdjzghn2eYQfNVuAqPtl6scYzDuys7DDd1dKON
DsN+fD0Pj4eN3Siag9l75xI/BNoLxWEFpXRDFuItZS0xUi0a7G/CZRsPAP53JAonJZL2D7QC55zD
Gc1vsEOJFAogeOTRRFqRV3ghBOSoJClEVRDmhImM7FlOkTsv/hRG04m+7NJ/KJMIhgI1OG1K2LYm
xwRlXxaBzF3OqhDAZgWtSDVBtjzpCfPJ+1OYtIiZ/cmGoW13Y3D/JBLLFVDGE9OYIpC0mDFHpDS3
xPI/zqySYjMShvg/IN3+FaVw8ovu6ccIquUBir3GSM8jl9C5/5ekyqqZnMro+cNmlMJ/t1Tig+Je
2dbdlrr0CoN3J5vlkXi95FvyfXWeCVAjIf6nTPGG0rs4sNlozacQP9y/gHjOn6ubn3HtTXGeohGK
knlGHA0c/haoMjObn2kui5F+ipx3PQ53aQWcuo94QgDhDDex/3GTnf4HOyN0r3bi5PZgd0p75p84
OfMLvkNInit7NqTkMlIgVbGUYqSOH0hA9JHIPhBsXZemsn1Y6a9LZzbyCd/15XisOFlB/ojKNHZU
p9DBXjo1ics0yYYmmmrPI3HB8d6m3gZEIcSu1iPydw6oOcdvTGjELVvJC2VME1Uk+MiUKttk95tV
9/9PUGV7KwrJXuvwyu9mLmfY/GUqRCInu/nyraeHvodAHhtk5kAR+hzmjl9U4BihKQplj+W8JeIp
2I8aL73gADzlwYl/ZKw8bUWfucc5S+xT+Z0SzH5LJ/CqVJMuNPOlQv/kV8Y5wfmiUcAPQmaPYu0p
J+f9b+0AeP29lqaTQw39hmkZeiH54r0BgALFV2lfMXhqz7Sh//ZTrynE93njk0FHlFI5P0fgC6KL
fodR/h4XSOn8z1dqlPRBd0aCH4Rtc1uzkQjPTrsbbTLxutAk7O5snS37OqsxhGXTjkQIMa2I9nmH
O0RhvVSr
`pragma protect end_protected
