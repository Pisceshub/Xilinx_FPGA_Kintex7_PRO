.GT_REFCLK0(gt_refclk0),
.altclk(q3_altclk_m),
.axisclk(q3_axisclk_m),
.apb3clk(q3_apb3clk_m),
.apb3presetn(q3_apb3presetn_m),
.apb3paddr(q3_apb3paddr_m),
.apb3penable(q3_apb3penable_m),
.apb3psel(q3_apb3psel_m),
.apb3pwdata(q3_apb3pwdata_m),
.apb3pwrite(q3_apb3pwrite_m),
.apb3prdata(q3_apb3prdata_m),
.apb3pready(q3_apb3pready_m),
.apb3pslverr(q3_apb3pslverr_m),
.bgbypassb(q3_bgbypassb_m),
.bgmonitorenb(q3_bgmonitorenb_m),
.bgpdb(q3_bgpdb_m),
.bgrcalovrdenb(q3_bgrcalovrdenb_m),
.bgrcalovrd(q3_bgrcalovrd_m),
.rcalenb(q3_rcalenb_m),
.trigackout0(q3_trigackout0_m),
.trigin0(q3_trigin0_m),
.ubenable(q3_ubenable_m),
.ubiolmbrst(q3_ubiolmbrst_m),
.ubmbrst(q3_ubmbrst_m),
.ctrlrsvdin1(q3_ctrlrsvdin1_m),
.ubintr(q3_ubintr_m),
.gpi(q3_gpi_m),
.ubrxuart(q3_ubrxuart_m),
.ctrlrsvdin0(q3_ctrlrsvdin0_m),
.correcterr(q3_correcterr_m),
.debugtracetvalid(q3_debugtracetvalid_m),
.refclk0_gtrefclkpd(q3_refclk0_gtrefclkpd_m),
.refclk0_clktestsig(q3_refclk0_clktestsig_m),
.refclk1_gtrefclkpd(q3_refclk1_gtrefclkpd_m),
.refclk1_clktestsig(q3_refclk1_clktestsig_m),
.trigackin0(q3_trigackin0_m),
.trigout0(q3_trigout0_m),
.ubinterrupt(q3_ubinterrupt_m),
.ubtxuart(q3_ubtxuart_m),
.uncorrecterr(q3_uncorrecterr_m),
.gpo(q3_gpo_m),
.debugtraceclk(q3_debugtraceclk_m),
.debugtracetdata(q3_debugtracetdata_m),
.ctrlrsvdout(q3_ctrlrsvdout_m),
.ch0_clkrsvd0(ch12_clkrsvd0_m),
.ch0_clkrsvd1(ch12_clkrsvd1_m),
.ch0_loopback(ch12_loopback_m),
.ch0_gtrsvd(ch12_gtrsvd_m),
.ch0_tstin(ch12_tstin_m),
.ch0_pcsrsvdout(ch12_pcsrsvdout_m),
.ch0_pinrsvdas(ch12_pinrsvdas_m),
.ch0_dmonfiforeset(ch12_dmonfiforeset_m),
.ch0_dmonitorclk(ch12_dmonitorclk_m),
.ch0_dmonitorout(ch12_dmonitorout_m),
.ch0_resetexception(ch12_resetexception_m),
.ch0_phyready(ch12_phyready_m),
.ch0_hsdppcsreset(ch12_hsdppcsreset_m),
.ch0_phyesmadaptsave(ch12_phyesmadaptsave_m),
.ch0_iloresetmask(ch12_iloresetmask_m),
.ch0_pcsrsvdin(ch12_pcsrsvdin_m),
.ch1_clkrsvd0(ch13_clkrsvd0_m),
.ch1_clkrsvd1(ch13_clkrsvd1_m),
.ch1_loopback(ch13_loopback_m),
.ch1_gtrsvd(ch13_gtrsvd_m),
.ch1_tstin(ch13_tstin_m),
.ch1_pcsrsvdout(ch13_pcsrsvdout_m),
.ch1_pinrsvdas(ch13_pinrsvdas_m),
.ch1_dmonfiforeset(ch13_dmonfiforeset_m),
.ch1_dmonitorclk(ch13_dmonitorclk_m),
.ch1_dmonitorout(ch13_dmonitorout_m),
.ch1_resetexception(ch13_resetexception_m),
.ch1_phyready(ch13_phyready_m),
.ch1_hsdppcsreset(ch13_hsdppcsreset_m),
.ch1_phyesmadaptsave(ch13_phyesmadaptsave_m),
.ch1_iloresetmask(ch13_iloresetmask_m),
.ch1_pcsrsvdin(ch13_pcsrsvdin_m),
.ch2_clkrsvd0(ch14_clkrsvd0_m),
.ch2_clkrsvd1(ch14_clkrsvd1_m),
.ch2_loopback(ch14_loopback_m),
.ch2_gtrsvd(ch14_gtrsvd_m),
.ch2_tstin(ch14_tstin_m),
.ch2_pcsrsvdout(ch14_pcsrsvdout_m),
.ch2_pinrsvdas(ch14_pinrsvdas_m),
.ch2_dmonfiforeset(ch14_dmonfiforeset_m),
.ch2_dmonitorclk(ch14_dmonitorclk_m),
.ch2_dmonitorout(ch14_dmonitorout_m),
.ch2_resetexception(ch14_resetexception_m),
.ch2_phyready(ch14_phyready_m),
.ch2_hsdppcsreset(ch14_hsdppcsreset_m),
.ch2_phyesmadaptsave(ch14_phyesmadaptsave_m),
.ch2_iloresetmask(ch14_iloresetmask_m),
.ch2_pcsrsvdin(ch14_pcsrsvdin_m),
.ch3_clkrsvd0(ch15_clkrsvd0_m),
.ch3_clkrsvd1(ch15_clkrsvd1_m),
.ch3_loopback(ch15_loopback_m),
.ch3_gtrsvd(ch15_gtrsvd_m),
.ch3_tstin(ch15_tstin_m),
.ch3_pcsrsvdout(ch15_pcsrsvdout_m),
.ch3_pinrsvdas(ch15_pinrsvdas_m),
.ch3_dmonfiforeset(ch15_dmonfiforeset_m),
.ch3_dmonitorclk(ch15_dmonitorclk_m),
.ch3_dmonitorout(ch15_dmonitorout_m),
.ch3_resetexception(ch15_resetexception_m),
.ch3_phyready(ch15_phyready_m),
.ch3_hsdppcsreset(ch15_hsdppcsreset_m),
.ch3_phyesmadaptsave(ch15_phyesmadaptsave_m),
.ch3_iloresetmask(ch15_iloresetmask_m),
.ch3_pcsrsvdin(ch15_pcsrsvdin_m),
.ch0_iloreset(ch12_iloreset_m),
.ch0_pcierstb(ch12_pcierstb_m),
.ch0_bufgtcemask(ch12_bufgtcemask_m),
.ch0_bufgtce(ch12_bufgtce_m),
.ch0_bufgtdiv(ch12_bufgtdiv_m),
.ch0_bufgtrstmask(ch12_bufgtrstmask_m),
.ch0_bufgtrst(ch12_bufgtrst_m),
.ch1_bufgtcemask(ch13_bufgtcemask_m),
.ch1_bufgtce(ch13_bufgtce_m),
.ch1_bufgtdiv(ch13_bufgtdiv_m),
.ch1_bufgtrstmask(ch13_bufgtrstmask_m),
.ch1_bufgtrst(ch13_bufgtrst_m),
.ch2_bufgtcemask(ch14_bufgtcemask_m),
.ch2_bufgtce(ch14_bufgtce_m),
.ch2_bufgtdiv(ch14_bufgtdiv_m),
.ch2_bufgtrstmask(ch14_bufgtrstmask_m),
.ch2_bufgtrst(ch14_bufgtrst_m),
.ch3_bufgtcemask(ch15_bufgtcemask_m),
.ch3_bufgtce(ch15_bufgtce_m),
.ch3_bufgtdiv(ch15_bufgtdiv_m),
.ch3_bufgtrstmask(ch15_bufgtrstmask_m),
.ch3_bufgtrst(ch15_bufgtrst_m),
.ch0_iloresetdone(ch12_iloresetdone_m),
.ch0_phystatus(ch12_phystatus_m),
.ch0_rxcdrhold(ch12_rxcdrhold_m),
.ch0_rxcdrovrden(ch12_rxcdrovrden_m),
.ch0_rxcdrreset(ch12_rxcdrreset_m),
.ch0_rxchbondi(ch12_rxchbondi_m),
.ch0_rxdapicodeovrden(ch12_rxdapicodeovrden_m),
.ch0_rxdapicodereset(ch12_rxdapicodereset_m),
.ch0_rxdlyalignreq(ch12_rxdlyalignreq_m),
.ch0_rxeqtraining(ch12_rxeqtraining_m),
.ch0_rxgearboxslip(ch12_rxgearboxslip_m),
.ch0_rxlatclk(ch12_rxlatclk_m),
.ch0_rxlpmen(ch12_rxlpmen_m),
.ch0_rxmldchaindone(ch12_rxmldchaindone_m),
.ch0_rxmldchainreq(ch12_rxmldchainreq_m),
.ch0_rxmlfinealignreq(ch12_rxmlfinealignreq_m),
.ch0_rxoobreset(ch12_rxoobreset_m),
.ch0_rxpcsresetmask(ch12_rxpcsresetmask_m),
.ch0_rxpd(ch12_rxpd_m),
.ch0_rxphalignreq(ch12_rxphalignreq_m),
.ch0_rxphalignresetmask(ch12_rxphalignresetmask_m),
.ch0_rxphdlypd(ch12_rxphdlypd_m),
.ch0_rxphdlyreset(ch12_rxphdlyreset_m),
.ch0_rxphsetinitreq(ch12_rxphsetinitreq_m),
.ch0_rxphshift180(ch12_rxphshift180_m),
.ch0_rxpmaresetmask(ch12_rxpmaresetmask_m),
.ch0_rxpolarity(ch12_rxpolarity_m),
.ch0_rxprbscntreset(ch12_rxprbscntreset_m),
.ch0_rxprbssel(ch12_rxprbssel_m),
.ch0_rxprogdivreset(ch12_rxprogdivreset_m),
.ch0_rxrate(ch12_rxrate_m),
.ch0_rxresetmode(ch12_rxresetmode_m),
.ch0_rxslide(ch12_rxslide_m),
.ch0_rxsyncallin(ch12_rxsyncallin_m),
.ch0_rxtermination(ch12_rxtermination_m),
.ch0_rxuserrdy(ch12_rxuserrdy_m),
.ch0_rxusrclk(ch12_rxusrclk_m),
.ch0_rx10gstat(ch12_rx10gstat_m),
.ch0_rxbufstatus(ch12_rxbufstatus_m),
.ch0_rxbyteisaligned(ch12_rxbyteisaligned_m),
.ch0_rxbyterealign(ch12_rxbyterealign_m),
.ch0_rxcdrlock(ch12_rxcdrlock_m),
.ch0_rxcdrphdone(ch12_rxcdrphdone_m),
.ch0_rxchanbondseq(ch12_rxchanbondseq_m),
.ch0_rxchanisaligned(ch12_rxchanisaligned_m),
.ch0_rxchanrealign(ch12_rxchanrealign_m),
.ch0_rxchbondo(ch12_rxchbondo_m),
.ch0_rxclkcorcnt(ch12_rxclkcorcnt_m),
.ch0_rxcominitdet(ch12_rxcominitdet_m),
.ch0_rxcommadet(ch12_rxcommadet_m),
.ch0_rxcomsasdet(ch12_rxcomsasdet_m),
.ch0_rxcomwakedet(ch12_rxcomwakedet_m),
.ch0_rxctrl0(ch12_rxctrl0_m),
.ch0_rxctrl1(ch12_rxctrl1_m),
.ch0_rxctrl2(ch12_rxctrl2_m),
.ch0_rxctrl3(ch12_rxctrl3_m),
.ch0_rxdataextendrsvd(ch12_rxdataextendrsvd_m),
.ch0_rxdatavalid(ch12_rxdatavalid_m),
.ch0_rxdata(ch12_rxdata_m),
.ch0_rxdccdone(ch12_rxdccdone_m),
.ch0_rxdlyalignerr(ch12_rxdlyalignerr_m),
.ch0_rxdlyalignprog(ch12_rxdlyalignprog_m),
.ch0_rxelecidle(ch12_rxelecidle_m),
.ch0_rxfinealigndone(ch12_rxfinealigndone_m),
.ch0_rxheadervalid(ch12_rxheadervalid_m),
.ch0_rxheader(ch12_rxheader_m),
.ch0_rxosintdone(ch12_rxosintdone_m),
.ch0_rxosintstarted(ch12_rxosintstarted_m),
.ch0_rxosintstrobedone(ch12_rxosintstrobedone_m),
.ch0_rxosintstrobestarted(ch12_rxosintstrobestarted_m),
.ch0_rxoutclk(),
.ch0_txoutclk(),
.ch0_rxphaligndone(ch12_rxphaligndone_m),
.ch0_rxphalignerr(ch12_rxphalignerr_m),
.ch0_rxphdlyresetdone(ch12_rxphdlyresetdone_m),
.ch0_rxphsetinitdone(ch12_rxphsetinitdone_m),
.ch0_rxphshift180done(ch12_rxphshift180done_m),
.ch0_rxpmaresetdone(ch12_rxpmaresetdone_m),
.ch0_rxprbserr(ch12_rxprbserr_m),
.ch0_rxprbslocked(ch12_rxprbslocked_m),
.ch0_rxresetdone(ch12_rxresetdone_m),
.ch0_rxsliderdy(ch12_rxsliderdy_m),
.ch0_rxstartofseq(ch12_rxstartofseq_m),
.ch0_rxstatus(ch12_rxstatus_m),
.ch0_rxsyncdone(ch12_rxsyncdone_m),
.ch0_rxvalid(ch12_rxvalid_m),
.ch0_txcomsas(ch12_txcomsas_m),
.ch0_txcomwake(ch12_txcomwake_m),
.ch0_txctrl0(ch12_txctrl0_m),
.ch0_txctrl1(ch12_txctrl1_m),
.ch0_txctrl2(ch12_txctrl2_m),
.ch0_txdapicodeovrden(ch12_txdapicodeovrden_m),
.ch0_txdapicodereset(ch12_txdapicodereset_m),
.ch0_txdataextendrsvd(ch12_txdataextendrsvd_m),
.ch0_txdata(ch12_txdata_m),
.ch0_txdeemph(ch12_txdeemph_m),
.ch0_txdetectrx(ch12_txdetectrx_m),
.ch0_txdiffctrl(ch12_txdiffctrl_m),
.ch0_txdlyalignreq(ch12_txdlyalignreq_m),
.ch0_txelecidle(ch12_txelecidle_m),
.ch0_txheader(ch12_txheader_m),
.ch0_txinhibit(ch12_txinhibit_m),
.ch0_txlatclk(ch12_txlatclk_m),
.ch0_txmaincursor(ch12_txmaincursor_m),
.ch0_txmargin(ch12_txmargin_m),
.ch0_txmldchaindone(ch12_txmldchaindone_m),
.ch0_txmldchainreq(ch12_txmldchainreq_m),
.ch0_txoneszeros(ch12_txoneszeros_m),
.ch0_txpausedelayalign(ch12_txpausedelayalign_m),
.ch0_txpcsresetmask(ch12_txpcsresetmask_m),
.ch0_txpd(ch12_txpd_m),
.ch0_txphalignreq(ch12_txphalignreq_m),
.ch0_txphalignresetmask(ch12_txphalignresetmask_m),
.ch0_txphdlypd(ch12_txphdlypd_m),
.ch0_txphdlyreset(ch12_txphdlyreset_m),
.ch0_txphdlytstclk(ch12_txphdlytstclk_m),
.ch0_txphsetinitreq(ch12_txphsetinitreq_m),
.ch0_txphshift180(ch12_txphshift180_m),
.ch0_txpicodeovrden(ch12_txpicodeovrden_m),
.ch0_txpicodereset(ch12_txpicodereset_m),
.ch0_txpippmen(ch12_txpippmen_m),
.ch0_txpippmstepsize(ch12_txpippmstepsize_m),
.ch0_txpisopd(ch12_txpisopd_m),
.ch0_txpmaresetmask(ch12_txpmaresetmask_m),
.ch0_txpolarity(ch12_txpolarity_m),
.ch0_txpostcursor(ch12_txpostcursor_m),
.ch0_txprbsforceerr(ch12_txprbsforceerr_m),
.ch0_txprbssel(ch12_txprbssel_m),
.ch0_txprecursor(ch12_txprecursor_m),
.ch0_txprogdivreset(ch12_txprogdivreset_m),
.ch0_txrate(ch12_txrate_m),
.ch0_txresetmode(ch12_txresetmode_m),
.ch0_txsequence(ch12_txsequence_m),
.ch0_txswing(ch12_txswing_m),
.ch0_txuserrdy(ch12_txuserrdy_m),
.ch0_txusrclk(ch12_txusrclk_m),
.ch0_tx10gstat(ch12_tx10gstat_m),
.ch0_txbufstatus(ch12_txbufstatus_m),
.ch0_txcomfinish(ch12_txcomfinish_m),
.ch0_txdccdone(ch12_txdccdone_m),
.ch0_txdlyalignerr(ch12_txdlyalignerr_m),
.ch0_txdlyalignprog(ch12_txdlyalignprog_m),
.ch0_txphaligndone(ch12_txphaligndone_m),
.ch0_txphalignerr(ch12_txphalignerr_m),
.ch0_txphalignoutrsvd(ch12_txphalignoutrsvd_m),
.ch0_txphdlyresetdone(ch12_txphdlyresetdone_m),
.ch0_txphshift180done(ch12_txphshift180done_m),
.ch0_txpmaresetdone(ch12_txpmaresetdone_m),
.ch0_txresetdone(ch12_txresetdone_m),
.ch0_txsyncdone(ch12_txsyncdone_m),
.ch0_gttxreset(ch12_gttxreset_m),
.ch0_txcominit(ch12_txcominit_m),
.ch0_txphsetinitdone(ch12_txphsetinitdone_m),
.ch0_txprogdivresetdone(ch12_txprogdivresetdone_m),
.ch0_txsyncallin(ch12_txsyncallin_m),
.ch1_iloreset(ch13_iloreset_m),
.ch1_pcierstb(ch13_pcierstb_m),
.ch1_iloresetdone(ch13_iloresetdone_m),
.ch1_phystatus(ch13_phystatus_m),
.ch1_rxcdrhold(ch13_rxcdrhold_m),
.ch1_rxcdrovrden(ch13_rxcdrovrden_m),
.ch1_rxcdrreset(ch13_rxcdrreset_m),
.ch1_rxchbondi(ch13_rxchbondi_m),
.ch1_rxdapicodeovrden(ch13_rxdapicodeovrden_m),
.ch1_rxdapicodereset(ch13_rxdapicodereset_m),
.ch1_rxdlyalignreq(ch13_rxdlyalignreq_m),
.ch1_rxeqtraining(ch13_rxeqtraining_m),
.ch1_rxgearboxslip(ch13_rxgearboxslip_m),
.ch1_rxlatclk(ch13_rxlatclk_m),
.ch1_rxlpmen(ch13_rxlpmen_m),
.ch1_rxmldchaindone(ch13_rxmldchaindone_m),
.ch1_rxmldchainreq(ch13_rxmldchainreq_m),
.ch1_rxmlfinealignreq(ch13_rxmlfinealignreq_m),
.ch1_rxoobreset(ch13_rxoobreset_m),
.ch1_rxpcsresetmask(ch13_rxpcsresetmask_m),
.ch1_rxpd(ch13_rxpd_m),
.ch1_rxphalignreq(ch13_rxphalignreq_m),
.ch1_rxphalignresetmask(ch13_rxphalignresetmask_m),
.ch1_rxphdlypd(ch13_rxphdlypd_m),
.ch1_rxphdlyreset(ch13_rxphdlyreset_m),
.ch1_rxphsetinitreq(ch13_rxphsetinitreq_m),
.ch1_rxphshift180(ch13_rxphshift180_m),
.ch1_rxpmaresetmask(ch13_rxpmaresetmask_m),
.ch1_rxpolarity(ch13_rxpolarity_m),
.ch1_rxprbscntreset(ch13_rxprbscntreset_m),
.ch1_rxprbssel(ch13_rxprbssel_m),
.ch1_rxprogdivreset(ch13_rxprogdivreset_m),
.ch1_rxrate(ch13_rxrate_m),
.ch1_rxresetmode(ch13_rxresetmode_m),
.ch1_rxslide(ch13_rxslide_m),
.ch1_rxsyncallin(ch13_rxsyncallin_m),
.ch1_rxtermination(ch13_rxtermination_m),
.ch1_rxuserrdy(ch13_rxuserrdy_m),
.ch1_rxusrclk(ch13_rxusrclk_m),
.ch1_rx10gstat(ch13_rx10gstat_m),
.ch1_rxbufstatus(ch13_rxbufstatus_m),
.ch1_rxbyteisaligned(ch13_rxbyteisaligned_m),
.ch1_rxbyterealign(ch13_rxbyterealign_m),
.ch1_rxcdrlock(ch13_rxcdrlock_m),
.ch1_rxcdrphdone(ch13_rxcdrphdone_m),
.ch1_rxchanbondseq(ch13_rxchanbondseq_m),
.ch1_rxchanisaligned(ch13_rxchanisaligned_m),
.ch1_rxchanrealign(ch13_rxchanrealign_m),
.ch1_rxchbondo(ch13_rxchbondo_m),
.ch1_rxclkcorcnt(ch13_rxclkcorcnt_m),
.ch1_rxcominitdet(ch13_rxcominitdet_m),
.ch1_rxcommadet(ch13_rxcommadet_m),
.ch1_rxcomsasdet(ch13_rxcomsasdet_m),
.ch1_rxcomwakedet(ch13_rxcomwakedet_m),
.ch1_rxctrl0(ch13_rxctrl0_m),
.ch1_rxctrl1(ch13_rxctrl1_m),
.ch1_rxctrl2(ch13_rxctrl2_m),
.ch1_rxctrl3(ch13_rxctrl3_m),
.ch1_rxdataextendrsvd(ch13_rxdataextendrsvd_m),
.ch1_rxdatavalid(ch13_rxdatavalid_m),
.ch1_rxdata(ch13_rxdata_m),
.ch1_rxdccdone(ch13_rxdccdone_m),
.ch1_rxdlyalignerr(ch13_rxdlyalignerr_m),
.ch1_rxdlyalignprog(ch13_rxdlyalignprog_m),
.ch1_rxelecidle(ch13_rxelecidle_m),
.ch1_rxfinealigndone(ch13_rxfinealigndone_m),
.ch1_rxheadervalid(ch13_rxheadervalid_m),
.ch1_rxheader(ch13_rxheader_m),
.ch1_rxosintdone(ch13_rxosintdone_m),
.ch1_rxosintstarted(ch13_rxosintstarted_m),
.ch1_rxosintstrobedone(ch13_rxosintstrobedone_m),
.ch1_rxosintstrobestarted(ch13_rxosintstrobestarted_m),
.ch1_rxphaligndone(ch13_rxphaligndone_m),
.ch1_rxphalignerr(ch13_rxphalignerr_m),
.ch1_rxphdlyresetdone(ch13_rxphdlyresetdone_m),
.ch1_rxphsetinitdone(ch13_rxphsetinitdone_m),
.ch1_rxphshift180done(ch13_rxphshift180done_m),
.ch1_rxpmaresetdone(ch13_rxpmaresetdone_m),
.ch1_rxprbserr(ch13_rxprbserr_m),
.ch1_rxprbslocked(ch13_rxprbslocked_m),
.ch1_rxresetdone(ch13_rxresetdone_m),
.ch1_rxsliderdy(ch13_rxsliderdy_m),
.ch1_rxstartofseq(ch13_rxstartofseq_m),
.ch1_rxstatus(ch13_rxstatus_m),
.ch1_rxsyncdone(ch13_rxsyncdone_m),
.ch1_rxvalid(ch13_rxvalid_m),
.ch1_txcomsas(ch13_txcomsas_m),
.ch1_txcomwake(ch13_txcomwake_m),
.ch1_txctrl0(ch13_txctrl0_m),
.ch1_txctrl1(ch13_txctrl1_m),
.ch1_txctrl2(ch13_txctrl2_m),
.ch1_txdapicodeovrden(ch13_txdapicodeovrden_m),
.ch1_txdapicodereset(ch13_txdapicodereset_m),
.ch1_txdataextendrsvd(ch13_txdataextendrsvd_m),
.ch1_txdata(ch13_txdata_m),
.ch1_txdeemph(ch13_txdeemph_m),
.ch1_txdetectrx(ch13_txdetectrx_m),
.ch1_txdiffctrl(ch13_txdiffctrl_m),
.ch1_txdlyalignreq(ch13_txdlyalignreq_m),
.ch1_txelecidle(ch13_txelecidle_m),
.ch1_txheader(ch13_txheader_m),
.ch1_txinhibit(ch13_txinhibit_m),
.ch1_txlatclk(ch13_txlatclk_m),
.ch1_txmaincursor(ch13_txmaincursor_m),
.ch1_txmargin(ch13_txmargin_m),
.ch1_txmldchaindone(ch13_txmldchaindone_m),
.ch1_txmldchainreq(ch13_txmldchainreq_m),
.ch1_txoneszeros(ch13_txoneszeros_m),
.ch1_txpausedelayalign(ch13_txpausedelayalign_m),
.ch1_txpcsresetmask(ch13_txpcsresetmask_m),
.ch1_txpd(ch13_txpd_m),
.ch1_txphalignreq(ch13_txphalignreq_m),
.ch1_txphalignresetmask(ch13_txphalignresetmask_m),
.ch1_txphdlypd(ch13_txphdlypd_m),
.ch1_txphdlyreset(ch13_txphdlyreset_m),
.ch1_txphdlytstclk(ch13_txphdlytstclk_m),
.ch1_txphsetinitreq(ch13_txphsetinitreq_m),
.ch1_txphshift180(ch13_txphshift180_m),
.ch1_txpicodeovrden(ch13_txpicodeovrden_m),
.ch1_txpicodereset(ch13_txpicodereset_m),
.ch1_txpippmen(ch13_txpippmen_m),
.ch1_txpippmstepsize(ch13_txpippmstepsize_m),
.ch1_txpisopd(ch13_txpisopd_m),
.ch1_txpmaresetmask(ch13_txpmaresetmask_m),
.ch1_txpolarity(ch13_txpolarity_m),
.ch1_txpostcursor(ch13_txpostcursor_m),
.ch1_txprbsforceerr(ch13_txprbsforceerr_m),
.ch1_txprbssel(ch13_txprbssel_m),
.ch1_txprecursor(ch13_txprecursor_m),
.ch1_txprogdivreset(ch13_txprogdivreset_m),
.ch1_txrate(ch13_txrate_m),
.ch1_txresetmode(ch13_txresetmode_m),
.ch1_txsequence(ch13_txsequence_m),
.ch1_txswing(ch13_txswing_m),
.ch1_txsyncallin(ch13_txsyncallin_m),
.ch1_txuserrdy(ch13_txuserrdy_m),
.ch1_txusrclk(ch13_txusrclk_m),
.ch1_tx10gstat(ch13_tx10gstat_m),
.ch1_txbufstatus(ch13_txbufstatus_m),
.ch1_txcomfinish(ch13_txcomfinish_m),
.ch1_txdccdone(ch13_txdccdone_m),
.ch1_txdlyalignerr(ch13_txdlyalignerr_m),
.ch1_txdlyalignprog(ch13_txdlyalignprog_m),
.ch1_txphaligndone(ch13_txphaligndone_m),
.ch1_txphalignerr(ch13_txphalignerr_m),
.ch1_txphalignoutrsvd(ch13_txphalignoutrsvd_m),
.ch1_txphdlyresetdone(ch13_txphdlyresetdone_m),
.ch1_txphshift180done(ch13_txphshift180done_m),
.ch1_txpmaresetdone(ch13_txpmaresetdone_m),
.ch1_txresetdone(ch13_txresetdone_m),
.ch1_txsyncdone(ch13_txsyncdone_m),
.ch1_gttxreset(ch13_gttxreset_m),
.ch1_txcominit(ch13_txcominit_m),
.ch1_txphsetinitdone(ch13_txphsetinitdone_m),
.ch1_txprogdivresetdone(ch13_txprogdivresetdone_m),
.ch2_iloreset(ch14_iloreset_m),
.ch2_pcierstb(ch14_pcierstb_m),
.ch2_iloresetdone(ch14_iloresetdone_m),
.ch2_phystatus(ch14_phystatus_m),
.ch2_rxcdrhold(ch14_rxcdrhold_m),
.ch2_rxcdrovrden(ch14_rxcdrovrden_m),
.ch2_rxcdrreset(ch14_rxcdrreset_m),
.ch2_rxchbondi(ch14_rxchbondi_m),
.ch2_rxdapicodeovrden(ch14_rxdapicodeovrden_m),
.ch2_rxdapicodereset(ch14_rxdapicodereset_m),
.ch2_rxdlyalignreq(ch14_rxdlyalignreq_m),
.ch2_rxeqtraining(ch14_rxeqtraining_m),
.ch2_rxgearboxslip(ch14_rxgearboxslip_m),
.ch2_rxlatclk(ch14_rxlatclk_m),
.ch2_rxlpmen(ch14_rxlpmen_m),
.ch2_rxmldchaindone(ch14_rxmldchaindone_m),
.ch2_rxmldchainreq(ch14_rxmldchainreq_m),
.ch2_rxmlfinealignreq(ch14_rxmlfinealignreq_m),
.ch2_rxoobreset(ch14_rxoobreset_m),
.ch2_rxpcsresetmask(ch14_rxpcsresetmask_m),
.ch2_rxpd(ch14_rxpd_m),
.ch2_rxphalignreq(ch14_rxphalignreq_m),
.ch2_rxphalignresetmask(ch14_rxphalignresetmask_m),
.ch2_rxphdlypd(ch14_rxphdlypd_m),
.ch2_rxphdlyreset(ch14_rxphdlyreset_m),
.ch2_rxphsetinitreq(ch14_rxphsetinitreq_m),
.ch2_rxphshift180(ch14_rxphshift180_m),
.ch2_rxpmaresetmask(ch14_rxpmaresetmask_m),
.ch2_rxpolarity(ch14_rxpolarity_m),
.ch2_rxprbscntreset(ch14_rxprbscntreset_m),
.ch2_rxprbssel(ch14_rxprbssel_m),
.ch2_rxprogdivreset(ch14_rxprogdivreset_m),
.ch2_rxrate(ch14_rxrate_m),
.ch2_rxresetmode(ch14_rxresetmode_m),
.ch2_rxslide(ch14_rxslide_m),
.ch2_rxsyncallin(ch14_rxsyncallin_m),
.ch2_rxtermination(ch14_rxtermination_m),
.ch2_rxuserrdy(ch14_rxuserrdy_m),
.ch2_rxusrclk(ch14_rxusrclk_m),
.ch2_rx10gstat(ch14_rx10gstat_m),
.ch2_rxbufstatus(ch14_rxbufstatus_m),
.ch2_rxbyteisaligned(ch14_rxbyteisaligned_m),
.ch2_rxbyterealign(ch14_rxbyterealign_m),
.ch2_rxcdrlock(ch14_rxcdrlock_m),
.ch2_rxcdrphdone(ch14_rxcdrphdone_m),
.ch2_rxchanbondseq(ch14_rxchanbondseq_m),
.ch2_rxchanisaligned(ch14_rxchanisaligned_m),
.ch2_rxchanrealign(ch14_rxchanrealign_m),
.ch2_rxchbondo(ch14_rxchbondo_m),
.ch2_rxclkcorcnt(ch14_rxclkcorcnt_m),
.ch2_rxcominitdet(ch14_rxcominitdet_m),
.ch2_rxcommadet(ch14_rxcommadet_m),
.ch2_rxcomsasdet(ch14_rxcomsasdet_m),
.ch2_rxcomwakedet(ch14_rxcomwakedet_m),
.ch2_rxctrl0(ch14_rxctrl0_m),
.ch2_rxctrl1(ch14_rxctrl1_m),
.ch2_rxctrl2(ch14_rxctrl2_m),
.ch2_rxctrl3(ch14_rxctrl3_m),
.ch2_rxdataextendrsvd(ch14_rxdataextendrsvd_m),
.ch2_rxdatavalid(ch14_rxdatavalid_m),
.ch2_rxdata(ch14_rxdata_m),
.ch2_rxdccdone(ch14_rxdccdone_m),
.ch2_rxdlyalignerr(ch14_rxdlyalignerr_m),
.ch2_rxdlyalignprog(ch14_rxdlyalignprog_m),
.ch2_rxelecidle(ch14_rxelecidle_m),
.ch2_rxfinealigndone(ch14_rxfinealigndone_m),
.ch2_rxheadervalid(ch14_rxheadervalid_m),
.ch2_rxheader(ch14_rxheader_m),
.ch2_rxosintdone(ch14_rxosintdone_m),
.ch2_rxosintstarted(ch14_rxosintstarted_m),
.ch2_rxosintstrobedone(ch14_rxosintstrobedone_m),
.ch2_rxosintstrobestarted(ch14_rxosintstrobestarted_m),
.ch2_rxphaligndone(ch14_rxphaligndone_m),
.ch2_rxphalignerr(ch14_rxphalignerr_m),
.ch2_rxphdlyresetdone(ch14_rxphdlyresetdone_m),
.ch2_rxphsetinitdone(ch14_rxphsetinitdone_m),
.ch2_rxphshift180done(ch14_rxphshift180done_m),
.ch2_rxpmaresetdone(ch14_rxpmaresetdone_m),
.ch2_rxprbserr(ch14_rxprbserr_m),
.ch2_rxprbslocked(ch14_rxprbslocked_m),
.ch2_rxresetdone(ch14_rxresetdone_m),
.ch2_rxsliderdy(ch14_rxsliderdy_m),
.ch2_rxstartofseq(ch14_rxstartofseq_m),
.ch2_rxstatus(ch14_rxstatus_m),
.ch2_rxsyncdone(ch14_rxsyncdone_m),
.ch2_rxvalid(ch14_rxvalid_m),
.ch2_txcomsas(ch14_txcomsas_m),
.ch2_txcomwake(ch14_txcomwake_m),
.ch2_txctrl0(ch14_txctrl0_m),
.ch2_txctrl1(ch14_txctrl1_m),
.ch2_txctrl2(ch14_txctrl2_m),
.ch2_txdapicodeovrden(ch14_txdapicodeovrden_m),
.ch2_txdapicodereset(ch14_txdapicodereset_m),
.ch2_txdataextendrsvd(ch14_txdataextendrsvd_m),
.ch2_txdata(ch14_txdata_m),
.ch2_txdeemph(ch14_txdeemph_m),
.ch2_txdetectrx(ch14_txdetectrx_m),
.ch2_txdiffctrl(ch14_txdiffctrl_m),
.ch2_txdlyalignreq(ch14_txdlyalignreq_m),
.ch2_txelecidle(ch14_txelecidle_m),
.ch2_txheader(ch14_txheader_m),
.ch2_txinhibit(ch14_txinhibit_m),
.ch2_txlatclk(ch14_txlatclk_m),
.ch2_txmaincursor(ch14_txmaincursor_m),
.ch2_txmargin(ch14_txmargin_m),
.ch2_txmldchaindone(ch14_txmldchaindone_m),
.ch2_txmldchainreq(ch14_txmldchainreq_m),
.ch2_txoneszeros(ch14_txoneszeros_m),
.ch2_txpausedelayalign(ch14_txpausedelayalign_m),
.ch2_txpcsresetmask(ch14_txpcsresetmask_m),
.ch2_txpd(ch14_txpd_m),
.ch2_txphalignreq(ch14_txphalignreq_m),
.ch2_txphalignresetmask(ch14_txphalignresetmask_m),
.ch2_txphdlypd(ch14_txphdlypd_m),
.ch2_txphdlyreset(ch14_txphdlyreset_m),
.ch2_txphdlytstclk(ch14_txphdlytstclk_m),
.ch2_txphsetinitreq(ch14_txphsetinitreq_m),
.ch2_txphshift180(ch14_txphshift180_m),
.ch2_txpicodeovrden(ch14_txpicodeovrden_m),
.ch2_txpicodereset(ch14_txpicodereset_m),
.ch2_txpippmen(ch14_txpippmen_m),
.ch2_txpippmstepsize(ch14_txpippmstepsize_m),
.ch2_txpisopd(ch14_txpisopd_m),
.ch2_txpmaresetmask(ch14_txpmaresetmask_m),
.ch2_txpolarity(ch14_txpolarity_m),
.ch2_txpostcursor(ch14_txpostcursor_m),
.ch2_txprbsforceerr(ch14_txprbsforceerr_m),
.ch2_txprbssel(ch14_txprbssel_m),
.ch2_txprecursor(ch14_txprecursor_m),
.ch2_txprogdivreset(ch14_txprogdivreset_m),
.ch2_txrate(ch14_txrate_m),
.ch2_txresetmode(ch14_txresetmode_m),
.ch2_txsequence(ch14_txsequence_m),
.ch2_txswing(ch14_txswing_m),
.ch2_txsyncallin(ch14_txsyncallin_m),
.ch2_txuserrdy(ch14_txuserrdy_m),
.ch2_txusrclk(ch14_txusrclk_m),
.ch2_tx10gstat(ch14_tx10gstat_m),
.ch2_txbufstatus(ch14_txbufstatus_m),
.ch2_txcomfinish(ch14_txcomfinish_m),
.ch2_txdccdone(ch14_txdccdone_m),
.ch2_txdlyalignerr(ch14_txdlyalignerr_m),
.ch2_txdlyalignprog(ch14_txdlyalignprog_m),
.ch2_txphaligndone(ch14_txphaligndone_m),
.ch2_txphalignerr(ch14_txphalignerr_m),
.ch2_txphalignoutrsvd(ch14_txphalignoutrsvd_m),
.ch2_txphdlyresetdone(ch14_txphdlyresetdone_m),
.ch2_txphshift180done(ch14_txphshift180done_m),
.ch2_txpmaresetdone(ch14_txpmaresetdone_m),
.ch2_txresetdone(ch14_txresetdone_m),
.ch2_txsyncdone(ch14_txsyncdone_m),
.ch2_gttxreset(ch14_gttxreset_m),
.ch2_txcominit(ch14_txcominit_m),
.ch2_txphsetinitdone(ch14_txphsetinitdone_m),
.ch2_txprogdivresetdone(ch14_txprogdivresetdone_m),
.ch3_iloreset(ch15_iloreset_m),
.ch3_pcierstb(ch15_pcierstb_m),
.ch3_iloresetdone(ch15_iloresetdone_m),
.ch3_phystatus(ch15_phystatus_m),
.ch3_rxcdrhold(ch15_rxcdrhold_m),
.ch3_rxcdrovrden(ch15_rxcdrovrden_m),
.ch3_rxcdrreset(ch15_rxcdrreset_m),
.ch3_rxchbondi(ch15_rxchbondi_m),
.ch3_rxdapicodeovrden(ch15_rxdapicodeovrden_m),
.ch3_rxdapicodereset(ch15_rxdapicodereset_m),
.ch3_rxdlyalignreq(ch15_rxdlyalignreq_m),
.ch3_rxeqtraining(ch15_rxeqtraining_m),
.ch3_rxgearboxslip(ch15_rxgearboxslip_m),
.ch3_rxlatclk(ch15_rxlatclk_m),
.ch3_rxlpmen(ch15_rxlpmen_m),
.ch3_rxmldchaindone(ch15_rxmldchaindone_m),
.ch3_rxmldchainreq(ch15_rxmldchainreq_m),
.ch3_rxmlfinealignreq(ch15_rxmlfinealignreq_m),
.ch3_rxoobreset(ch15_rxoobreset_m),
.ch3_rxpcsresetmask(ch15_rxpcsresetmask_m),
.ch3_rxpd(ch15_rxpd_m),
.ch3_rxphalignreq(ch15_rxphalignreq_m),
.ch3_rxphalignresetmask(ch15_rxphalignresetmask_m),
.ch3_rxphdlypd(ch15_rxphdlypd_m),
.ch3_rxphdlyreset(ch15_rxphdlyreset_m),
.ch3_rxphsetinitreq(ch15_rxphsetinitreq_m),
.ch3_rxphshift180(ch15_rxphshift180_m),
.ch3_rxpmaresetmask(ch15_rxpmaresetmask_m),
.ch3_rxpolarity(ch15_rxpolarity_m),
.ch3_rxprbscntreset(ch15_rxprbscntreset_m),
.ch3_rxprbssel(ch15_rxprbssel_m),
.ch3_rxprogdivreset(ch15_rxprogdivreset_m),
.ch3_rxrate(ch15_rxrate_m),
.ch3_rxresetmode(ch15_rxresetmode_m),
.ch3_rxslide(ch15_rxslide_m),
.ch3_rxsyncallin(ch15_rxsyncallin_m),
.ch3_rxtermination(ch15_rxtermination_m),
.ch3_rxuserrdy(ch15_rxuserrdy_m),
.ch3_rxusrclk(ch15_rxusrclk_m),
.ch3_rx10gstat(ch15_rx10gstat_m),
.ch3_rxbufstatus(ch15_rxbufstatus_m),
.ch3_rxbyteisaligned(ch15_rxbyteisaligned_m),
.ch3_rxbyterealign(ch15_rxbyterealign_m),
.ch3_rxcdrlock(ch15_rxcdrlock_m),
.ch3_rxcdrphdone(ch15_rxcdrphdone_m),
.ch3_rxchanbondseq(ch15_rxchanbondseq_m),
.ch3_rxchanisaligned(ch15_rxchanisaligned_m),
.ch3_rxchanrealign(ch15_rxchanrealign_m),
.ch3_rxchbondo(ch15_rxchbondo_m),
.ch3_rxclkcorcnt(ch15_rxclkcorcnt_m),
.ch3_rxcominitdet(ch15_rxcominitdet_m),
.ch3_rxcommadet(ch15_rxcommadet_m),
.ch3_rxcomsasdet(ch15_rxcomsasdet_m),
.ch3_rxcomwakedet(ch15_rxcomwakedet_m),
.ch3_rxctrl0(ch15_rxctrl0_m),
.ch3_rxctrl1(ch15_rxctrl1_m),
.ch3_rxctrl2(ch15_rxctrl2_m),
.ch3_rxctrl3(ch15_rxctrl3_m),
.ch3_rxdataextendrsvd(ch15_rxdataextendrsvd_m),
.ch3_rxdatavalid(ch15_rxdatavalid_m),
.ch3_rxdata(ch15_rxdata_m),
.ch3_rxdccdone(ch15_rxdccdone_m),
.ch3_rxdlyalignerr(ch15_rxdlyalignerr_m),
.ch3_rxdlyalignprog(ch15_rxdlyalignprog_m),
.ch3_rxelecidle(ch15_rxelecidle_m),
.ch3_rxfinealigndone(ch15_rxfinealigndone_m),
.ch3_rxheadervalid(ch15_rxheadervalid_m),
.ch3_rxheader(ch15_rxheader_m),
.ch3_rxosintdone(ch15_rxosintdone_m),
.ch3_rxosintstarted(ch15_rxosintstarted_m),
.ch3_rxosintstrobedone(ch15_rxosintstrobedone_m),
.ch3_rxosintstrobestarted(ch15_rxosintstrobestarted_m),
.ch3_rxphaligndone(ch15_rxphaligndone_m),
.ch3_rxphalignerr(ch15_rxphalignerr_m),
.ch3_rxphdlyresetdone(ch15_rxphdlyresetdone_m),
.ch3_rxphsetinitdone(ch15_rxphsetinitdone_m),
.ch3_rxphshift180done(ch15_rxphshift180done_m),
.ch3_rxpmaresetdone(ch15_rxpmaresetdone_m),
.ch3_rxprbserr(ch15_rxprbserr_m),
.ch3_rxprbslocked(ch15_rxprbslocked_m),
.ch3_rxresetdone(ch15_rxresetdone_m),
.ch3_rxsliderdy(ch15_rxsliderdy_m),
.ch3_rxstartofseq(ch15_rxstartofseq_m),
.ch3_rxstatus(ch15_rxstatus_m),
.ch3_rxsyncdone(ch15_rxsyncdone_m),
.ch3_rxvalid(ch15_rxvalid_m),
.ch3_txcomsas(ch15_txcomsas_m),
.ch3_txcomwake(ch15_txcomwake_m),
.ch3_txctrl0(ch15_txctrl0_m),
.ch3_txctrl1(ch15_txctrl1_m),
.ch3_txctrl2(ch15_txctrl2_m),
.ch3_txdapicodeovrden(ch15_txdapicodeovrden_m),
.ch3_txdapicodereset(ch15_txdapicodereset_m),
.ch3_txdataextendrsvd(ch15_txdataextendrsvd_m),
.ch3_txdata(ch15_txdata_m),
.ch3_txdeemph(ch15_txdeemph_m),
.ch3_txdetectrx(ch15_txdetectrx_m),
.ch3_txdiffctrl(ch15_txdiffctrl_m),
.ch3_txdlyalignreq(ch15_txdlyalignreq_m),
.ch3_txelecidle(ch15_txelecidle_m),
.ch3_txheader(ch15_txheader_m),
.ch3_txinhibit(ch15_txinhibit_m),
.ch3_txlatclk(ch15_txlatclk_m),
.ch3_txmaincursor(ch15_txmaincursor_m),
.ch3_txmargin(ch15_txmargin_m),
.ch3_txmldchaindone(ch15_txmldchaindone_m),
.ch3_txmldchainreq(ch15_txmldchainreq_m),
.ch3_txoneszeros(ch15_txoneszeros_m),
.ch3_txpausedelayalign(ch15_txpausedelayalign_m),
.ch3_txpcsresetmask(ch15_txpcsresetmask_m),
.ch3_txpd(ch15_txpd_m),
.ch3_txphalignreq(ch15_txphalignreq_m),
.ch3_txphalignresetmask(ch15_txphalignresetmask_m),
.ch3_txphdlypd(ch15_txphdlypd_m),
.ch3_txphdlyreset(ch15_txphdlyreset_m),
.ch3_txphdlytstclk(ch15_txphdlytstclk_m),
.ch3_txphsetinitreq(ch15_txphsetinitreq_m),
.ch3_txphshift180(ch15_txphshift180_m),
.ch3_txpicodeovrden(ch15_txpicodeovrden_m),
.ch3_txpicodereset(ch15_txpicodereset_m),
.ch3_txpippmen(ch15_txpippmen_m),
.ch3_txpippmstepsize(ch15_txpippmstepsize_m),
.ch3_txpisopd(ch15_txpisopd_m),
.ch3_txpmaresetmask(ch15_txpmaresetmask_m),
.ch3_txpolarity(ch15_txpolarity_m),
.ch3_txpostcursor(ch15_txpostcursor_m),
.ch3_txprbsforceerr(ch15_txprbsforceerr_m),
.ch3_txprbssel(ch15_txprbssel_m),
.ch3_txprecursor(ch15_txprecursor_m),
.ch3_txprogdivreset(ch15_txprogdivreset_m),
.ch3_txrate(ch15_txrate_m),
.ch3_txresetmode(ch15_txresetmode_m),
.ch3_txsequence(ch15_txsequence_m),
.ch3_txswing(ch15_txswing_m),
.ch3_txsyncallin(ch15_txsyncallin_m),
.ch3_txuserrdy(ch15_txuserrdy_m),
.ch3_txusrclk(ch15_txusrclk_m),
.ch3_tx10gstat(ch15_tx10gstat_m),
.ch3_txbufstatus(ch15_txbufstatus_m),
.ch3_txcomfinish(ch15_txcomfinish_m),
.ch3_txdccdone(ch15_txdccdone_m),
.ch3_txdlyalignerr(ch15_txdlyalignerr_m),
.ch3_txdlyalignprog(ch15_txdlyalignprog_m),
.ch3_txphaligndone(ch15_txphaligndone_m),
.ch3_txphalignerr(ch15_txphalignerr_m),
.ch3_txphalignoutrsvd(ch15_txphalignoutrsvd_m),
.ch3_txphdlyresetdone(ch15_txphdlyresetdone_m),
.ch3_txphshift180done(ch15_txphshift180done_m),
.ch3_txpmaresetdone(ch15_txpmaresetdone_m),
.ch3_txresetdone(ch15_txresetdone_m),
.ch3_txsyncdone(ch15_txsyncdone_m),
.ch3_gttxreset(ch15_gttxreset_m),
.ch3_txcominit(ch15_txcominit_m),
.ch3_txphsetinitdone(ch15_txphsetinitdone_m),
.ch3_txprogdivresetdone(ch15_txprogdivresetdone_m),
.hsclk0_lcpllclkrsvd0(q3_hsclk0_lcpllclkrsvd0_m),
.hsclk0_lcpllclkrsvd1(q3_hsclk0_lcpllclkrsvd1_m),
.hsclk0_lcpllfbdiv(q3_hsclk0_lcpllfbdiv_m),
.hsclk0_lcpllpd(q3_hsclk0_lcpllpd_m),
.hsclk0_lcpllrefclksel(q3_hsclk0_lcpllrefclksel_m),
.hsclk0_lcpllresetbypassmode(q3_hsclk0_lcpllresetbypassmode_m),
.hsclk0_lcpllresetmask(q3_hsclk0_lcpllresetmask_m),
.hsclk0_lcpllreset(q3_hsclk0_lcpllreset_m),
.hsclk0_lcpllrsvd0(q3_hsclk0_lcpllrsvd0_m),
.hsclk0_lcpllrsvd1(q3_hsclk0_lcpllrsvd1_m),
.hsclk0_lcpllsdmdata(q3_hsclk0_lcpllsdmdata_m),
.hsclk0_lcpllsdmtoggle(q3_hsclk0_lcpllsdmtoggle_m),
.hsclk0_rpllclkrsvd0(q3_hsclk0_rpllclkrsvd0_m),
.hsclk0_rpllclkrsvd1(q3_hsclk0_rpllclkrsvd1_m),
.hsclk0_rpllfbdiv(q3_hsclk0_rpllfbdiv_m),
.hsclk0_rpllpd(q3_hsclk0_rpllpd_m),
.hsclk0_rpllrefclksel(q3_hsclk0_rpllrefclksel_m),
.hsclk0_rpllresetbypassmode(q3_hsclk0_rpllresetbypassmode_m),
.hsclk0_rpllresetmask(q3_hsclk0_rpllresetmask_m),
.hsclk0_rpllreset(q3_hsclk0_rpllreset_m),
.hsclk0_rpllrsvd0(q3_hsclk0_rpllrsvd0_m),
.hsclk0_rpllrsvd1(q3_hsclk0_rpllrsvd1_m),
.hsclk0_rpllsdmdata(q3_hsclk0_rpllsdmdata_m),
.hsclk0_rpllsdmtoggle(q3_hsclk0_rpllsdmtoggle_m),
.hsclk0_lcpllfbclklost(q3_hsclk0_lcpllfbclklost_m),
.hsclk0_lcpllrefclklost(q3_hsclk0_lcpllrefclklost_m),
.hsclk0_rpllfbclklost(q3_hsclk0_rpllfbclklost_m),
.hsclk0_rpllrefclklost(q3_hsclk0_rpllrefclklost_m),
.hsclk0_lcpllrefclkmonitor(q3_hsclk0_lcpllrefclkmonitor_m),
.hsclk0_rpllrefclkmonitor(q3_hsclk0_rpllrefclkmonitor_m),
.hsclk0_lcpllrsvdout(q3_hsclk0_lcpllrsvdout_m),
.hsclk0_rpllrsvdout(q3_hsclk0_rpllrsvdout_m),
.hsclk1_lcpllclkrsvd0(q3_hsclk1_lcpllclkrsvd0_m),
.hsclk1_lcpllclkrsvd1(q3_hsclk1_lcpllclkrsvd1_m),
.hsclk1_lcpllfbdiv(q3_hsclk1_lcpllfbdiv_m),
.hsclk1_lcpllpd(q3_hsclk1_lcpllpd_m),
.hsclk1_lcpllrefclksel(q3_hsclk1_lcpllrefclksel_m),
.hsclk1_lcpllresetbypassmode(q3_hsclk1_lcpllresetbypassmode_m),
.hsclk1_lcpllresetmask(q3_hsclk1_lcpllresetmask_m),
.hsclk1_lcpllreset(q3_hsclk1_lcpllreset_m),
.hsclk1_lcpllrsvd0(q3_hsclk1_lcpllrsvd0_m),
.hsclk1_lcpllrsvd1(q3_hsclk1_lcpllrsvd1_m),
.hsclk1_lcpllsdmdata(q3_hsclk1_lcpllsdmdata_m),
.hsclk1_lcpllsdmtoggle(q3_hsclk1_lcpllsdmtoggle_m),
.hsclk1_rpllclkrsvd0(q3_hsclk1_rpllclkrsvd0_m),
.hsclk1_rpllclkrsvd1(q3_hsclk1_rpllclkrsvd1_m),
.hsclk1_rpllfbdiv(q3_hsclk1_rpllfbdiv_m),
.hsclk1_rpllpd(q3_hsclk1_rpllpd_m),
.hsclk1_rpllrefclksel(q3_hsclk1_rpllrefclksel_m),
.hsclk1_rpllresetbypassmode(q3_hsclk1_rpllresetbypassmode_m),
.hsclk1_rpllresetmask(q3_hsclk1_rpllresetmask_m),
.hsclk1_rpllreset(q3_hsclk1_rpllreset_m),
.hsclk1_rpllrsvd0(q3_hsclk1_rpllrsvd0_m),
.hsclk1_rpllrsvd1(q3_hsclk1_rpllrsvd1_m),
.hsclk1_rpllsdmdata(q3_hsclk1_rpllsdmdata_m),
.hsclk1_rpllsdmtoggle(q3_hsclk1_rpllsdmtoggle_m),
.hsclk1_lcpllfbclklost(q3_hsclk1_lcpllfbclklost_m),
.hsclk1_lcpllrefclklost(q3_hsclk1_lcpllrefclklost_m),
.hsclk1_rpllfbclklost(q3_hsclk1_rpllfbclklost_m),
.hsclk1_rpllrefclklost(q3_hsclk1_rpllrefclklost_m),
.hsclk1_lcpllrefclkmonitor(q3_hsclk1_lcpllrefclkmonitor_m),
.hsclk1_rpllrefclkmonitor(q3_hsclk1_rpllrefclkmonitor_m),
.hsclk1_lcpllrsvdout(q3_hsclk1_lcpllrsvdout_m),
.hsclk1_rpllrsvdout(q3_hsclk1_rpllrsvdout_m),
.s0_axis_tready(m9_axis_tready_m),
.s0_axis_tdata(m9_axis_tdata_m),
.s0_axis_tlast(m9_axis_tlast_m),
.s0_axis_tvalid(m9_axis_tvalid_m),
.s1_axis_tready(m10_axis_tready_m),
.s1_axis_tdata(m10_axis_tdata_m),
.s1_axis_tlast(m10_axis_tlast_m),
.s1_axis_tvalid(m10_axis_tvalid_m),
.s2_axis_tready(m11_axis_tready_m),
.s2_axis_tdata(m11_axis_tdata_m),
.s2_axis_tlast(m11_axis_tlast_m),
.s2_axis_tvalid(m11_axis_tvalid_m),
.pcielinkreachtarget(q3_pcielinkreachtarget_m),
.pcieltssm(q3_pcieltssm_m),
.rxmarginclk(q3_rxmarginclk_m),
.rxmarginreqcmd(q3_rxmarginreqcmd_m),
.rxmarginreqlanenum(q3_rxmarginreqlanenum_m),
.rxmarginreqpayld(q3_rxmarginreqpayld_m),
.rxmarginreqreq(q3_rxmarginreqreq_m),
.rxmarginresack(q3_rxmarginresack_m),
.rxmarginresreq(q3_rxmarginresreq_m),
.rxmarginreqack(q3_rxmarginreqack_m),
.rxmarginrescmd(q3_rxmarginrescmd_m),
.rxmarginreslanenum(q3_rxmarginreslanenum_m),
.rxmarginrespayld(q3_rxmarginrespayld_m),
.m0_axis_tready(s9_axis_tready_m),
.m0_axis_tdata(s9_axis_tdata_m),
.m0_axis_tlast(s9_axis_tlast_m),
.m0_axis_tvalid(s9_axis_tvalid_m),
.m1_axis_tready(s10_axis_tready_m),
.m1_axis_tdata(s10_axis_tdata_m),
.m1_axis_tlast(s10_axis_tlast_m),
.m1_axis_tvalid(s10_axis_tvalid_m),
.m2_axis_tready(s11_axis_tready_m),
.m2_axis_tdata(s11_axis_tdata_m),
.m2_axis_tlast(s11_axis_tlast_m),
.m2_axis_tvalid(s11_axis_tvalid_m),
.gtpowergood(q3_gtpowergood_m),
.ch0_rxprogdivresetdone(ch12_rxprogdivresetdone_m),
.ch0_gtrxreset(ch12_gtrxreset_m),
.ch0_cdrbmcdrreq(ch12_cdrbmcdrreq_m),
.ch0_cdrfreqos(ch12_cdrfreqos_m),
.ch0_cdrincpctrl(ch12_cdrincpctrl_m),
.ch0_cdrstepdir(ch12_cdrstepdir_m),
.ch0_cdrstepsq(ch12_cdrstepsq_m),
.ch0_cdrstepsx(ch12_cdrstepsx_m),
.ch0_cfokovrdfinish(ch12_cfokovrdfinish_m),
.ch0_cfokovrdpulse(ch12_cfokovrdpulse_m),
.ch0_cfokovrdstart(ch12_cfokovrdstart_m),
.ch0_eyescanreset(ch12_eyescanreset_m),
.ch0_eyescantrigger(ch12_eyescantrigger_m),
.ch0_eyescandataerror(ch12_eyescandataerror_m),
.ch0_cfokovrdrdy0(ch12_cfokovrdrdy0_m),
.ch0_cfokovrdrdy1(ch12_cfokovrdrdy1_m),
.ch1_rxprogdivresetdone(ch13_rxprogdivresetdone_m),
.ch1_gtrxreset(ch13_gtrxreset_m),
.ch1_cdrbmcdrreq(ch13_cdrbmcdrreq_m),
.ch1_cdrfreqos(ch13_cdrfreqos_m),
.ch1_cdrincpctrl(ch13_cdrincpctrl_m),
.ch1_cdrstepdir(ch13_cdrstepdir_m),
.ch1_cdrstepsq(ch13_cdrstepsq_m),
.ch1_cdrstepsx(ch13_cdrstepsx_m),
.ch1_cfokovrdfinish(ch13_cfokovrdfinish_m),
.ch1_cfokovrdpulse(ch13_cfokovrdpulse_m),
.ch1_cfokovrdstart(ch13_cfokovrdstart_m),
.ch1_eyescanreset(ch13_eyescanreset_m),
.ch1_eyescantrigger(ch13_eyescantrigger_m),
.ch1_eyescandataerror(ch13_eyescandataerror_m),
.ch1_cfokovrdrdy0(ch13_cfokovrdrdy0_m),
.ch1_cfokovrdrdy1(ch13_cfokovrdrdy1_m),
.ch2_rxprogdivresetdone(ch14_rxprogdivresetdone_m),
.ch2_gtrxreset(ch14_gtrxreset_m),
.ch2_cdrbmcdrreq(ch14_cdrbmcdrreq_m),
.ch2_cdrfreqos(ch14_cdrfreqos_m),
.ch2_cdrincpctrl(ch14_cdrincpctrl_m),
.ch2_cdrstepdir(ch14_cdrstepdir_m),
.ch2_cdrstepsq(ch14_cdrstepsq_m),
.ch2_cdrstepsx(ch14_cdrstepsx_m),
.ch2_cfokovrdfinish(ch14_cfokovrdfinish_m),
.ch2_cfokovrdpulse(ch14_cfokovrdpulse_m),
.ch2_cfokovrdstart(ch14_cfokovrdstart_m),
.ch2_eyescanreset(ch14_eyescanreset_m),
.ch2_eyescantrigger(ch14_eyescantrigger_m),
.ch2_eyescandataerror(ch14_eyescandataerror_m),
.ch2_cfokovrdrdy0(ch14_cfokovrdrdy0_m),
.ch2_cfokovrdrdy1(ch14_cfokovrdrdy1_m),
.ch3_rxprogdivresetdone(ch15_rxprogdivresetdone_m),
.ch3_gtrxreset(ch15_gtrxreset_m),
.ch3_cdrbmcdrreq(ch15_cdrbmcdrreq_m),
.ch3_cdrfreqos(ch15_cdrfreqos_m),
.ch3_cdrincpctrl(ch15_cdrincpctrl_m),
.ch3_cdrstepdir(ch15_cdrstepdir_m),
.ch3_cdrstepsq(ch15_cdrstepsq_m),
.ch3_cdrstepsx(ch15_cdrstepsx_m),
.ch3_cfokovrdfinish(ch15_cfokovrdfinish_m),
.ch3_cfokovrdpulse(ch15_cfokovrdpulse_m),
.ch3_cfokovrdstart(ch15_cfokovrdstart_m),
.ch3_eyescanreset(ch15_eyescanreset_m),
.ch3_eyescantrigger(ch15_eyescantrigger_m),
.ch3_eyescandataerror(ch15_eyescandataerror_m),
.ch3_cfokovrdrdy0(ch15_cfokovrdrdy0_m),
.ch3_cfokovrdrdy1(ch15_cfokovrdrdy1_m),
.hsclk0_lcplllock(q3_hsclk0_lcplllock_m),
.hsclk0_rplllock(q3_hsclk0_rplllock_m),
.hsclk1_lcplllock(q3_hsclk1_lcplllock_m),
.hsclk1_rplllock(q3_hsclk1_rplllock_m),
.debugtraceready(q3_debugtracetready_m),
.ch0_txmstreset     (ch12_msttxreset_m),
.ch0_txmstresetdone (ch12_msttxresetdone_m),
.ch1_txmstreset     (ch13_msttxreset_m),
.ch1_txmstresetdone (ch13_msttxresetdone_m),
.ch2_txmstreset     (ch14_msttxreset_m),
.ch2_txmstresetdone (ch14_msttxresetdone_m),
.ch3_txmstreset     (ch15_msttxreset_m),
.ch3_txmstresetdone (ch15_msttxresetdone_m),
.ch0_rxmstreset      ( ch12_mstrxreset_m ),
.ch0_rxmstresetdone  ( ch12_mstrxresetdone_m),
.ch1_rxmstreset      ( ch13_mstrxreset_m),
.ch1_rxmstresetdone  ( ch13_mstrxresetdone_m),
.ch2_rxmstreset      ( ch14_mstrxreset_m),
.ch2_rxmstresetdone  ( ch14_mstrxresetdone_m),
.ch3_rxmstreset      ( ch15_mstrxreset_m),
.ch3_rxmstresetdone  ( ch15_mstrxresetdone_m),
.rxn(q3_gt_quad_base_serial_rxn),
.rxp(q3_gt_quad_base_serial_rxp),
.txn(q3_gt_quad_base_serial_txn),
.txp(q3_gt_quad_base_serial_txp),
.refclk0_gtrefclkpdint(q3_refclk0_gtrefclkpdint),
.pipenorthin(pipenorthoutq2_to_pipenorthinq3),
.resetdone_northin(resetdone_northout_q2_to_resetdone_northin_q3), 
.rxpinorthin(rxpinorthout_q2_to_rxpinorthin_q3), 
.txpinorthin(txpinorthout_q2_to_txpinorthin_q3), 
.pipesouthout( pipesouthin_q2_to_pipesouthout_q3),  
.resetdone_southout(resetdone_southin_q2_to_resetdone_southout_q3), 
.rxpisouthout(rxpisouthin_q2_to_rxpsouthout_q3), 
.txpisouthout(txpisouthin_q2_to_txpsouthout_q3)
