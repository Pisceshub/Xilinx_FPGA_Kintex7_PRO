`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37344)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9JQaMgpupSUIgDmsbAQQ3DL5vC3Qu8u6xK0RRu4TKgP3/eH23+g56iUo
jPZoY4COC+nKJ3OZ7Sb9z1Kyz4UaOr66gyKURpFvQScknKtIVqiSQm8PeE9TBY0wRBLH/W6f9WPN
OACuVEw/1VIkd7am6hZuE2tsIZedoeflOAA94+0pd+gieXWG1iIRamWXUnuKb0lDHzgot5Bio6xk
89TDsmu6OlxuFc56qqfOAhr0mhDR3N/d4vu2E4YBQmVZkzcYdxUPItGcRxnIaXPFYew30QoTWUw3
pYZH6VDEnLX9VYwkZs+qjybDauc7qpBN0HHkjJ0tSrDORpuWEY+HeEnvRmwna6LSOVIy1/H8BNVx
3KjJtiEey1WokqBni8xXnoUV2XkhZJiZiv4AmrHwW2Wv/gI/Zxbp+sSZKJFbL2ARGBOHglN7tJrs
gIgolGK3LFtYg2VkOpdIR4/FCQ4hVGh4oSbw5i7loxlsd8VtUne1MfLxGgjlhAa3oaYX48swYJdt
8h2VkfWzYs3WspXX9HEp4jbmjapK67oMtK8pfTgHEKCvwL1YPF5YH0IFfYEuP7PVZq3VcRLsFZ63
LSLQxgXYprO/ROjsKTjGlkYhGZh2J+/O2EFEt76YnVywyqo7SvPbWVcvfkapFBOgqqgOeO6zTxGK
dZASnlxY+sHUXDsObWLp13hZacOn+E6GCFeaXa15QU/qcriMQEZ6plU8cWqrN8u23OCGnjfXDRN2
+XYECSeUNU0oVee6EAyyMZIRIa7CBqYEIrZ3AmVIkqv1XUKuTNZHYBaT52AXoRL6UlEK4U+yzFbi
fUM5Y1B14+BHDKzznXTCf6opYS3oDAJxWruqibjaxPTqWY3cSMtGWVlBsOMoKfwbfwRWsP8T1EuA
JSuwyU47/SFjd1iKKUnb2e/dHFclRzfHY2sKymZuhJYg/mMFNSLmoEEb62+U/ePCXiZ+QF8S1FGO
5fA7FFbLyWfM8TFoPeZoZ7RehS3kGL+b8Dnr0uPpvx1FWY4xVf6OBKteMJFIsMPFWThb/oWIZLIk
TZiAP4RufrlRgCzhU3Ap2i/7CJpOedCiZOEso4J2BOY9n7RNp8Xf34GUKPljaskCUuiUjf9XWQUf
6T+eeIPFwZtygFDrfRKauqXAtIDm8ZubggOtsTY9LjbyYaqHCzgZNzdMH2PFw0UsWU1k39nne7Ie
b86CEjR1zmzu5R74XwMjDxeSlD38JHyp+UO5omHLhFy3zB8qFMoQYehV71YMjFSjq8V2wuji8cCg
sTNjR8aEtJVZy3cUiNpeXkbGuEHSfDLklUTVI3iN9ZtXtyGhvLs5Iah7emQAMGuLk4zyqr0gNUl2
ogWa37FiQ3KFiibuJO7hV96uj2d2xduIJ44UFXimWsiO8MejCPLETRW2dPLMYGMan9pte9PJhiXx
w7Zb5DwOgXNnzGZvS+gfjdfOqhqOqG3xfBTW5PzJTuSBwc8J2OZjuF5+942ft8o0wCN4BerAPRaH
/iMOtFRAJOoSfO48NAyQdip5uI34bK/Gm94AVrsocbLl3GoB30olVsYzZ1BlA1snQRLOIPu9/dRM
VG1zrqPqWVir18o7STRBZBlkSOL8E21HXbwkSgzcMBjrVWja+zQkJtCGt6Mu0girWIJh2VYcvvC7
eIoltZoF7QACXNbU3dJycsrvV4q4wL7svEshhTlyD+GWMrGbQDyEf6s2uVO0lOeJwrRkvnlXP1A2
66OUEFEBpljH5hgadWyWMePz+J5E/kTN8vlJBn7pi82wVZ3N4UYzGBb51ucnc1Z3gPmEh0CHR1/6
9n1vNhvBPtUDuz2esxCfjt3Bc3+Tpf5/1+8gpht6sanSl8VFDr/sW1fxToLmoUWfodkBClDMDooV
v60i5Jt3RlTHxMLQWAyrInn8YIT+S2IGTawsoK1POz/g6Yt9aIEbVlsXAxVWYd/rkkjQ5TuEasCO
FMSueRJW0KUrBWi5ZvKBUCM1HPjQ4Xy9wQhWGzaRAjaFiwJ6KERwL7pjS4jqa0E0uwEqLyupwIPs
lEPwkCdqBMb2y1ncMU6d1jP0riBAUZ76864wvvmAzLCRUmmBuiYiE9K0csc9cR232a8QcjBMkK3R
LjxzkdNqDeXgy5zenLbdaJ5L1j1vIHLA9k58MBIrQaVh/YL1MHE3d3Cl3SeUrjlAy3POGbrjcNh5
ozdjctaJ6VI4wDiyqBeBA4Xk9uwGtvKXUCqPs91nR6+OKed+PCWmsaaU9f2nZIgR3IgJSEBLd5W3
H37MGu2rd8185WW4NKk5dfeUEqe1R2ZmRufr0UyC/BjsYMDWquyUhEhFS/9d9wlcLMvpWa69v/my
HT1iKP4i52RQbtp6Pp6cqjK2OOb3kpwpGESdblLu/ek5wW3E6UzA3qXzvTxo25HhVh7e5xF6cvNe
bS3zq4e9TJWP6Ms+zcQVhKNa6+N1XCCzoJAIylPg4FwLG/FQSZKaj/54qJpQaMp9rjdc6Ix9RCHR
DBT3D3cCgwpTnVET++inYLpfCyY2vY0G8k6ORbRNm7XLdfwAYTejNRh5pS/1pAf02X436yS0oyby
O0Cf3uO9oGiZv4enlBjCkuc/s0t94W6bPY22G4W/s6+3W40HJR28qskfM5haS/xw7RnyhjYF4eY5
ixiwWnH3w7C4PGjr+MvxCBE+o2+F70ktpkN9u0PcrWyv2gjGJTyGCs0Aa0SCi4qTcd7w1T0ACyGt
ujvXbNDR2ey3FD5hjV9bf2AMq2gQzm5IbkZwtPPgU0ApDXSIfFxcWr0KWBqLUdWaLrSKmADb+WoD
7fHiqNFsRo6Tbr1hfrocCjpZ8dskr50trps8QXo2UjLOipvvXfnYzfpRIDMsIL2PamrywxvyCWF2
TYXoO2cEFU3WfiX66l9Zkco0aL+iG2AV5/XW3S/OJgno+vAgAk/jsRAhfQ4RIEdgCFXRWBcHaLS/
PB/I+rDC3XGaVlRYsqiZmxdCJwmM5SEnxNmo1QT45Ib/gA8f5o7h/3WmFPqw/viZIX6Io2uHYQLj
4iXM3R00cRjsG8m2S8wPZ9CN54yFP2x4Eq2VUyqKmWBU0rT0shAOEp0LQX/EMi6MeG5Eo+zylleN
8uTax+BEwyejUq+yRN9YtW9MyLdvtGLj7LpnWp6bsZWfTuDASQFjQ+qc006qhi8nH2Q7rbrDEv3e
LtBtgHSQ0xvH0D18MY3a7LSPyCxg9jX4P/EyKhjxFb9DtnogbiOcZ1xDAzVTlh0BnMybPsFSXXSq
RhdglRXLiu5RaZXZJmscy1HfOAmSFtalQao7XXZBidGGpuSldhyuTdP/YLgCsNNyY7dqj/bFwILz
NZIQ10cmiC5CxGGD8wCJB6B20isRKTOl31MByAnuzHKyaa1oZ4+dT4OIMOjJackgXeEp1t+5GVRN
r1BaejNDih0LjYhmIA9gSeQLw0qWU/wM6yiyFK4s76qUyxlH0KLXmzwZA1WnF+0vWrULOADXn8Fs
1q4238lAnp2vrqP65t87zorbPbxILLOf97d21s69zMRl2ng9++iR0JSRz3QEomqstfdjzpwg+wkK
ART5N2czt75dr1cfjuatT+KQagQEMYFTgLcevhrozFuYTYFk0UO6/90uBTqMfverAzah+Q+JPQKx
Et5HUSEwM9waCG5VdhVYCN6+FTb4arp8I5IiyQdnkYT065AFlcpiY/flSFJ0GX1+fa6TehYEXV6Y
8O0u6QtPAZjiy1Wq5z6FQ0YwMke4KicIzFC0Ca6P7iZtyzNkefaBKOiiDPsGSrSCz0DRriPSrkwH
2YSv7Is9AExf+ZX1AVAq9rtfHaM0BGfdZ/XLLHo2Q7bbhTA84Z0b6qiKBFpwkKuVn05o9tK0BKyk
JD/DjE100WQOoMnRCNale5QwVLo9Lozly7bnuVGbqrJiSqph5PgmEA5O9qTtrdjHqJwIntL+PxvC
kmhbLB0nKa4N+IzsJxN/0ztbHsk+JvlpHUYF9qjAnBKePGxUP5OJlgUD8eH+Zu1ufIym2Ua2EOP9
Ide8p01jU8zpohKQIGQznCzdFq/PwcVny5g3vsOXykwan0T9tS+Dc9IoQiTNKotlyWFLGGwEx7uu
awqY+/5fJctji5G+FJKJBfKS34cMEfU3BJrHmaP1lUEwx9Hqa0tg6ej8zAJboLBCsM7qvOsMoQRB
djKn/piHkkiGISY3bQuMFEJyxoUrCKqqYhXyXlo/1SpQENfzsJK4+NyPYvodnS8Awlna+H045+iT
UK+XgsHJoGR+xWT+rm/Rg6lyO5H1FPQO/eR7xQfFe5V8PsIpTTKhnfAJeFHsHarGTYaaMGCJRIBv
k0fo1UFBTNzC34TtbuSswYrZkVyy+2vsqzyaryFSXG1G+af616ItV4NtLMX+cPBmcZrA9mwCj6BH
mcqRNgwMVAuYUjm/t4UnT95fYefbYT99ZaiLWBPLRdiMB+dEOUCzQvxV9kkDptoaTCEG/1DtGNTs
YYb7tm292Z97xOg/1AovbKu8NmlNkENZxagX5PcnjPtR7zOofPC5uWgJxLxsKNJOc33VyO18rJbe
SNA9pn6RAJyWTTR5dHuE4SUCTX6u3dk4x5uLBEKteHxKZFj97XH1oGJm929Xk4dgO7wnaSX7rrQN
YAmfsUUfQPqHn+Hr8iZn5shYfnvG86mjsrD+AyBSjd18F7pnA+4Y7xDzKHSqHeaepngu+xcWHnL2
8sbmf5vHsJPEHQy3pOS6EuO8qTgjOjEC40bve7XadHsCzTAfx8pnzDq6wGitoVONw0nfW1oR/iC/
gnYh3P/Q8O5NgwIRKnoLntgRKacMGlDsrRDn4t6ctw8nogWwEiRHoJT4jsMiyO2LZ5HH3QOv8DZc
RvkHyXJhFs/IrK8OeVwfhBVnA3StRiK8hQ5HQe1UZndJSDcC1SGHbmkjMb8G6u99CnaUb2KzmTOq
B0n6KK/6JDp9gHEHo7zVVlmIGyCjWXqZpyrXzjLBBd/AybEDMF+5ULC70Vh1eThULI/s26XlUYFC
jHW2bf+y5HW4GeNnpi1QcX7kYKlZhI3BoGNBVWatD+ZDcmA1Yr3n8As0H416C/sJqeYFQmcSJ5oV
uuAXno9MBhR9HKJax3gKdCY4FKvFGk5s3lZpoEQDr5Q3CYcws26rd2pcF+V/VLUH/6fDIy1nMbGD
OCwoEd3Lqx/xJdm8aInGmmxozvlu4dyVHbGiuyUKavsC2bEq+AxlbdBgfw+f3GugUXY3Vqsh74ty
sQOMU4LOsue9pHcL/UUoM08SLmBBKlnY3qQIxyr4Jzmn2i3H0WphhcOOJkQItY+hGrMOSzjoYWr3
ejDyOk8Bkg6UpYWa1RmpnzIq/6vdiMA2ClQYCybwkMdcsAZmRpn0RkIDhjVIUdLEa9wuIIYmt9ji
CNbifQqbGNf85Zes2A/+9Bou7UMAZP1nkfyyFtiX41YqghZZEfhAYVqen+xHvz80uD1nUPhVUz7z
ffwNq1U9CyDuZgGx/M4SbN+yf1DUzDOeyuaKnMjGZiYbrf0sxbFmTeLsMM1sHSBxVwC1P0qemuvY
qFlItHhkoBEu3r2AAge2wlvS9QRQeJes+MAaoWcjMA5CFdJ8hX5QoYzH7gX/Y8TQ3tR1RNg/czv8
LO8Co2S60DxWmKfWLcFwztRu+EJTqH/8wAb9PUa0fkb8cx0LCbgcbLOztwMhEa613TDmfZnk82sJ
CDXW7xEHK0uryHHIBqWAzz9/tdA3arlGFTPCPJWU+tUaiTGP/Ir+cQ1H5If5OqaG5rAjevOBiyt8
MgM8hravL+w0KA1pIsoP2iA4/Tt/2BDSibvaE4N/SC3YwdglBQ4qQN6qn8uNT62n8FyIbx0bVGrk
hBYcX7SkMiWZYbeQSAIzTx2LiikzzNWM6HeG13pMZXrMWJdwO2QfDRxCaUsA/ENEoqcTV0hpn6CB
Q5a8it7x4+4jnjg5ojdkxG0F0i2aHmzENZLtENd3OatqSAFo9ZJ/DlKwuDqlZ3L+ImPa1Oj2hr9w
QYeI6W0vgn4WU4qWSTxninzzPnbQFG2WwRXRj7tNRml/Iz0L1qx1Qv0/HWrw9ui3G/GdsP2YdZgL
6t4JFCaQ8zU2UfYNRpgl/bm7Lhec1frbi/phIPGX4sETJQHgINsyVJK+W8CvVrf5mEPLx5erv9Fu
H7byL6fuY6w3RCtk7TCxr7UPI8i7OxBhZG8CAoHAjDTAOtB86k7J6lafYB5UoWHo/ac4+ecepJhU
+fU6o9FLr1VQjc/xc3rSLSeFiUOpGClkRYyCK/ANY96z5I3cxhC5TFkzgvPsaP3OhxkCpiFW8SVh
/RCnf/91tBas8847B8XMbTb+FhRXzd7xIypE2ENYDkt+TWp+Zn6vWUSQgZ7iAK5NupY2b1uNGbgm
DeiIXI01H+ErN6p62+7wlCltFwU3f4B8TYPeTF5CX/inNV70VlbOzLItXTKjZX3PLq2E1gm6i0Hy
eZPEanFqznrZCLD3LchTmQURBOdK+hZ/IhhNxFi3zXxnJe06d14cMiU66PztUUhWdpn0h+xIvUDq
7nhuPKTscgG9RZG/XzmHHIlUifxS0AsfgckUkg73MF5To1ls7HfwapfGKDBdNQl66+r0Z0ggtwbD
H/sEhHbkllaw6eNi/6PE4F3uEiZSBhm45TEXJxb+xYzCVhg6k9vXf/AJUfLRLIfFcEynYI3EPKfG
sa9+X87GlnG/KDt17deDNPHWe08nzoRlf2p2eiOWE7hy07hN0mN+kSC2Jt9Vg4Zr5FfWIX73MHUu
7pm+Bw/xNTYUTyFLcV9S5hZ6+Pp1aajxJEQUYWGkFMP8AyFE3iZj30N0dEB5/7dvapAAbUQfacp4
4+EPanEc7jPhmgKnMxfPc45OMYgB+QmuBOIzHjpVe7RxdEk3vNhV1UHP0wwGbaVUD6IUsJhjTrkK
8JfiwSnnmpDYnD4xTWqK1KDShsjJp1A3eT9NQJALYWk64JBfsvE7CZjwBazIhO221iggcY7b0a7p
BDeI5XDN4bFV/NsBE5ulq7ODz80VbUG53Q9azXfxSxK1bXfbxgossvot3Pu5IoStAoUuKQXWgteh
AjFmq4I7H4XXyEK62Cj8jP8xLujyqF7dQ+12Hpn3iDeK7D1taCSCC4AzLdw3gqFSEY4jUNNU1ZiG
Aiem+ROPrkyWxJM9j9vOwZP23WQVAaHdNY91q82XSVyZujAnXqkbGyRtftCPmGqYGgbKB8qgOsW9
QGAJQUdqZ1e7RY5bnLbrf2Hjoin6wiAfiFlk/BhJqrBXLxI+qwXPwwVfOVjRYJ/aZ3hlDpt+tzWq
J0yjR/rQnsJln9a7njUWR3YIqpo1EmsBw0LUiv19b/8j22ZNQUkkxmMjMVuECHr29KS2kwMPmAXT
j76v5FspcNKnGiChU12TOL0QuPTtQZ0l15yPiGS6xwvgqz37Kv0MLkbKR+07cmY0CU2Q1NGijIZB
fy3PYgqFVsadARhrSyFpx9J3FuNfxotKcluAa8MLZ0y8wWRcli51YjiPkDSWoeDW7dv0JEj2EA7x
f6+3kcd6I5YThtGESxq9+JmJlcKTQFmTC3Odyb/sn+s1GNw9hEQ4vpsV49JF7O5W7XizgvKFA+rw
RK23hX/dWxmI+hJtri+UdMf0QzgJRti3/yZweMQkiK50HyQAFQW/JGSpDjuOMeyTkl15fOMYEzNN
psx0FtSZXiTnqKxkSEVhAYD1jQRuviSFFY6qdz+YskhCiIHSHYul1wyRn0kbPRk8FCr6zmCxU56k
90Z0mRi/MaupOFd370QaxNnZQ4/YTXHM0yrURzWpz9rO1K1r4YKkkLhrDwhhQZwVaaMLGcy0VE2c
hn7opyZOmkrGt8iqzLLwXd0ot/5DFW8uF3QdW9w3tnHeJyLFfjGzC0DJ47985dZwOd3pjd/ica0R
vHePWTwp3mCZ5FCq3t8yc6qP5/8I9r/F2R3OY5MHHJV5JF+7fHP5CgbrWPyFk8xh4x+4VaI0AaWX
Bo3aYW8bXc1UsEQEYptXjAJpgM7BhMTckSYVmUmFGyW2+abvOFcIbhvHhbqoA19rCuhhn2M5fwr5
QBWCSJ+tf1UuXpsSV62bjgH/kOMnz0QnS+6Jz7bEddikioiwzlHT1eqDz8PbI6/RhGM9frPmtVvi
BqgB5PGbVHDCvjNqHepcrUIomXWaQtyD+lGx1SiG0vwiBpeJLjTbq4cB3BScXfY5SA4/DTKpgH3Z
DRalrsy7XE3xfzg4JVfC9oEVXZzRJlvgPEOMl2XZlaB6yd8qJfICNDtfjkg0Q7RZ7X9FZk12vOIC
gJmJsCJ+6hn0A+gQF1YEBwEuY6hgLk/8wlPsNxfVeDL7uiZnmbH/VGFOxrgtyQaMte/6nDL5Tb2A
ToJ40MkIgKUAQGVyYTrViBUM1fIOGpledKBb+WG9OfjXrMuOb1jt/CQ9iNzN7sjseGOnUb5JuERl
TYZYtxyf1Z++fYvHXn/9pg+iM8XVuQHiDRG5J25LRw/jndtCCtDRWrJ+o9RJHpc4RF5/zDrr8LE4
C+iAyuDB/MQqyhRtklGSlGBi5rtm2jfL1kRblfg5uwGW0tZDwy6aaNgP7lxLlnxH6v8oc74Z54OR
hs66sSX49hJpBKCMlAHlJbnfpzyjT6VHfv9+haWnfJ9MYKDqJEdnh3Bzz9Mbsoj1tsApcIcoAcoV
G8jNOApanTIJ4YsmPcCcQnslLVpvRgtnhNJ0SSB4J+s8TizeXaTd2uzu2/QnX7cEACOj1rx6vg2f
wY1IMt4Hm4Eyb3Lx3+FEDKh0304fOBIQEC0mfLRw0P0Xy8BdCoTdTTwhssOkG9OxFfBwYNWhEgTu
lgRXTRsGd9rEv/5S3dyUzwrdkEfrz9ZWA3wUeE0TUCHhBzQTuly5g2K8GO9oGtvBnJkOOzU4qZ4S
xywcx/ot2t0BfTUeFWRvGVMe6S3HNO/gcEsNDOraO87NIHWNklPWK7vHsxfin/4ih9rte/ILtXsE
8K+sKX92IjVKq5tKnlTtfDBQhhN9zdprOWAtqHQO5+uzLlNUCtHC2zCLleJWYTE1UTUUGpwi4tL5
G+KwRMnT+lmUrbJVXpcbG6r9rMrojfCPgXkIKdvaXzAGRmgkDT5VEjuNJwAoJbOCty1pnlf8fKqj
5GZIa81x6Zy8jLeaJFs63NCVYp/tUrAR/mqy0opHNXHQOEvEFJ9wDOa4wj5IcURZ3TB1dF4SOP9d
2Wh6zel2NAc7YdqnmD1z0IRTRAJriCON9Db+AbJIU3r/KqosieWsiEjxCBkhhhYBRZm12gHCndQC
ihVa0EqIlfuBhdfqIiEFGLMZ3gRwTMkIgn370H8Ysr4TSR3ORhQY5EU2AsbZ3kkejbrBtV6/p4rQ
P2pO8tn+k9u+i9nbP2bP4Flw9+TKbeJZNSGmm3jk5V36iGRS8PrdQRAeRie+zs05XEXVHjEhQlPh
qBKvm/NeFkpXrgqHVcnmSctOPuFSPSMKT0Ums+Oh1ecvdznptk84Ilr9xB7Pkj4UBUn8if9Xmbqo
YAcrkk6APT2YHXHU6juV8tR4zeV63rRoj3VWJ5kKl0nlgYXO13Vo3MJ4bbtG995Ub5lhCBK9IMP8
9a3nGLAbKlI+3j1jDOGu99ttQlclbLUex+tNvPN/+D7P7n+FPbQ/x8dvreIY+7cfxI+W1n+bE07a
Qy+oLHFOffIBuwgkwNWbfkwVsr61XtaDZvWOmcu9mTVFY9x0vSHgkRVbMQHNE3vm5/1u4AI05F1a
ZRIV7685n5worekNpHVc8xPEidWGx+8WiVNcXYT/fzMacv+2dj0h0jK6g4tbdggfuU9j+jfbhO3y
pOnS9oFkHzScw44ZCcZFioeAVXkLTn0hbQLEqZ7UUZw/04nihRV1Y4289OsiQnbrCDpXeKCEogQV
d7lJttW3jPQq9nQc6nsfJT/iul9PdS9HP66J19KwXcvkqhwz5sHzd5tLwfDcFmW+D+dOXFL1ReX9
qLEaUdIt+UPduF6u0L/gejdIpojSJnqzJw8qyW7ZIl1GA7IEkwFdBcDweSM8BkhQWaEk+VFU1nUW
RE7V7hyC+TXU0/uDMY530SgglpBC5mbXNuu2Ch0qpRxBCsgI7lmL5jJFm3z7n7ud+1gW32NEPIg4
fvu5mFym1tMTFEsNLkmylikZicDQh83qNGV8jsbQt8U/nJb3frF6ioETCBUqs9W1cdLw/mbNU4xE
BwASTDKLYwV1jX24fa+6Q+hNtQSvkmAFonC3rDLU7GRwQLTZZ6rVcVIGtdW6B3gIoMol8QZade+C
PxjUjqrNSZY5vX7OPJgHn4xcsUgNT4UNiyLWDkGcXTT861li50kazBJKHyLkXzuACqfF09FxfWx6
iFJLSM4l6/a6f/JTbsPWkRNYsbD5DkTAO4k6aCU9G3nK+qUwTQ7OQFUgbG7eW7V4/cfjl9gb2sZk
eaFOBQ3/x1Kh2fzTIZPzAEt2sRQASwQJmEetA3dwzRUiZmBNKVSWVkvumBgNZ7skv4Uh4iRBKgGf
+fl8kdCb3eobvqv7TseqX8bOYs1pBFzTNHmWcGgAXZOEaG9y3234j4jlLTle+1LCXW8EZioVAmSe
Pr503hHcQC80+b7ZkeUC3h8qtDjdTuuiRV4dl6w91D/v3T53T1jL2kFvtnxI/dLYtgBPwKf0juzW
Kdqp3wfnQBSJtEAN627Ww8DDXKWIYiKf34Y3nJXfqe8WhouaRyrqkpf7fIJWWbsImIRepT7TdBAa
Hhf+YHNGwmPQ+Bli2qKL76us8z7IG1e80o1TWUf6o7dfDqM6Zv9L5Y1HbrCI/qw70H/G0STAH8DG
kHuOKiCj4ogqgBw7Y6jpzDcdO424Ig9Tg5RHJLVwCypZieQsCo5efUa7OCkIdJKH34tTZWjCdr/A
9O8ktAAmJHzr0BDANSqeWl2yQH1NPgKM+9eAROw0qXUTxHx84XESkESY/fXsBZZ7TqnVmk68NHdn
aGUL/lkY0cu4eti6dmQweDjeJdmBmyuuRZTyN/7qYWKMUiXM3/N1hV33P8b8E2QE1Z0yGajN9PWQ
PuAasTqntinpWvBWhHS8kux+fXQFs65xn/p5zPppJRAskd7j3EFneG66o9fEZwHsEcWTPS/h+4Vu
X9sbg5ScP0FEum29RB5zWt8ZV1TERne+FM8obAhxlQU2BhHE1kpmC3P4v9Kdq3g0lDBHkU1iLim0
1KLtGvjtRF5ETJZ2fKEtNZXr7H1AlmveIBTy6HecOYOE5Dazt67vEWWWUhg26u/GGZIGGiIQ3Ure
+t6YcWHJQXlciPYKpnJl1Tu3+ty9u+uN5FBpIMZrhSHH87BKjnWa+e3IyuebyTiFzQqEOzfNMxnc
lyhlGEOLfPn76F5wTjziVuZsfx3VEKrogVU9HGBLMw+Yow21pTJxhOloDkaZExNgFMmZFXQIQzQf
T0xxHYorBiIa8yuU1YrAka1CZ35wGJBymi99sZ4sDZXa/T1HpSa7lX+VP0M2HdO9n3uCXwkvjSvz
t5VwdiCIPsLqE9c/COSgssoz6bcIaDTFjWke3b/cMoOqHJLf2MdgakodvbHG1zq5bwMEWbjdOf4O
oprxPxd0WZo62ajNhRvaqJQnv6i2suwIAVAWqIj1GHOEQqx3aZVjzyD4fi9F+dq1DQqNNDx9jUjG
5oyy/3FJ+vpxjQviOaWFokv++uHlBVCtYEviOFSt9B2JmZAt/604vBrRpQsWXEid+aAf8g4dxnXu
3PeDfY8OI3qbF/KtwYO8PwW4Pf2YrtO46teLz2LkqAFs7AEwSZqP6K89hRqyX44QbQe3xvhSbKPX
4wioU91v+QIyaFjGLJcmO1YIQWv0GoKFzcB+VHaupTb9ZlknO8oiW0MgUaZiORKs30DH/s6ZMuGt
Yum1GrJqrfbH8gQMoGQx++el9WZxidtdVBy0rom1OGY1gDOuQ6bLRy7vtteDRUwn3N7NZjbHUiMN
BBOa4YmORLwroovkCMqM3Aq8S6aRGSNOqTeJf92TEkpyWC4ag8sL3V1shCeYUOzakJk2gthbyXzB
VE0osh1UbOfX2+CO6FYif+NrmBrackijmSR3uBp/BBt2YAmt1hM/jb4tm2js84jcImZ9APReZ3S9
5JjKmk2MubeEct/CumZ359Sg6Hf8UImd4FHdBo937LyzTSyZMkwLeLqPEaCMERXGo/SLwKQrLVWd
kmvZ7FBDKilNEn2s1lEgVqaf40xsh5iWDxdrCbk944BePlsSif7bhRivwy+4+0Nbogon7whmWdng
K4hR4GtHeO49ZQFAh8zxxLMT8RkWtN6DluwEc1zVDjFjF3ztP8GYCuV+VXslkJLEA9dUj5g5ONEC
0UM6xpQz95xdO3wDiLCDUhHViPm9ElKqm5xOvP6MHB2dBGVxOupu+nTgPBgGrCmW19f8Pa9wATxB
y8nJNkJdd8g34vM7T/VCSHb9w5om49f3VEjU9UApV0k4flbAWqQ89S9ImUE1EdmcRdsTOkTTaaXh
NG8KSezk6fDVMBAByU9g01VSDTUkhKHLxc1DoMsEBC1NKKUGyhZsqKnkBXOz4RdInjBYmvTqqUN4
TkI3AU3OpMj9Eg9844GLLmUMt5oYCJba8qLkjgBoYTDxFMtC5uwNxFkCNvmzxu6/HnGmB73QMCBH
MD9yafWOzbsrAEwCRWvdKauzWbXkpRfNv8G8jmU2mbf7Fm+2pGoBdXDHnFL39Y5j4LjqIQq+h3PN
kdIebrlqkevSeCazoTk0FNNWAYK4ehEkKllsptf//7Wn4/Z7Q1+Jl9uW4hOgSx4WNRboDbctYzze
2CSVg70zI0YPdbmPT56y6VO3uNKQY7gq8irH4Hm4cPRgcGNzSq6ftkoW3mYVDzapBEAuLa6cfOuL
UVSt4lM7WuljYJsn2flfT1gQW/2+iZLdeITjGrAbq8KTiuNA0S/7U3+a13n5NMWJTqRI31yZ7uxL
uHWiet9AorKbv1a0zKgesvqHcLKNrFrnOf5XNF7p1CZgOD22sYyvQZ9ARAhcT3MZQAooxgpj3YnD
yhmlrU8ZCPWBkHo0MNauK2ioeqTWR/1bOIThVEEMGaK9qZOOCtOWbO4ZntCXNec+jB4mye7LycWV
7j+0tyGnHZ22oIl6SscK45ffMxdnbwjarxBzhHntd0dpmRARRAg6oIIALGJ6ncn41aP2avXiNaxy
C9/WHFqrj/gVqQ6dug3EQg9svrklaBl4uX2gU3x748v2+AdCnnIZl89SQJF7CW+iFBpf2hOWBQbi
fblV7YgR5TPX+g8leWip2cI1uWk2Ss5prPW5D0Y4MULsnAFFv6a1jnTRpPgTYwIncd31TnCW7/IT
GdBYILLtlQLwVyvd263er+Q3dxz5IwqECk4F1T5xUHwP4nOAJmZzVeEfhbLYsGx9I3Y7z1VfzIm9
73RznKuypC/cnHuRpVQ/dkSxBf2Py600ZmdNFKk3bXoBHlZm+MCXGhhmACIDm+sL2CgZ/hmS3GjG
HfLtCKbe3vZYY9WE6A1la9J79GKP41Di96E7VEeiExquKJpshyTM81P6lG8ptDnP/Lqn7wLPmAnt
l+ymSGizfrB2PPF2W1x4J5uUz8Fkr+e/+DRkUiry2efAugA5dZrXqBqk+2NunWyQU6Bw1n/Zc/q7
Qoc0QuPG39uEMOYBCmw2xEgnwfunZumRh+q8xxrwKUNrmuGkwbTmdL/y0hue5nTiIVecn1TA6NO9
i4qQhofPKRFSgZBgfrTCD65DubHA8Ny96oN0MS0rcoFZmf1Ngl8T0oM30p2jtwW+5AIyKjk3R2sV
sEImNcu7jnisSWfRbAX8n5nFG+Ed+GW1dUvuDsOIbN13UYvN5kNx3C9evUbZhnr4jutyHX7jKeSv
ZU9qA62yYsv9NbAc57xkOOW1WsdghsCkPTJoCLPh+ulB4UJkJ1Q269+XLP2RdDVHQxDOu1Zz+nBP
ujJtUE8TILywYuoA2UbFPAOd3VZaIwZml+vmefwjRZ/cq5xM+tr9GGimeE7tW/jyrZileAS+k0j+
Nre/4DQ6wR0we3/28hggvCainGEjm+1JDr606O22kGd4lTXPA7IS/1U6eVHbAI0k+55hr9Z2ukoJ
3Fn2uflYopcIARomYxEl19XvvRozpwUPkdWqVxBKJT9S6woKIjQW67bs0gBX0SJ9PIftJJewNCOd
rE/Z5q7n8e8s54Pbzunrip8QCmFNFCPadfUM6fHgt7QzHvBWYr+zm3m7PIug9h6BQOVBPKEI4yBn
gPKA+eP+ZVokz/lnx1CBaZnAI483IiSk7h74tV0tYgPz8Ynl6bBFGJCAcgsdf3mHggZLvXurVIfE
aaqLcMcmH3oleX2ypwT+UMGcg4I1SPSoA9eNB7XjhWhmWKymO2HimkU1h0r0AkrIhMBE/8IRpQa6
sMcXvS6XVurWN1krVPTgPqaETCPFJZTDtu3HcCFblB+M3KyzSDwb8p7cO4s8DEGd1g5cXWAKcEId
4xuwLecUTchJOCpRQuGizm2N1HrQJfSlh3XTwVRveAjTSwVUgUDYE9AiX4ZAU16R302MkA1eOqyT
jGPzjX8tjByEUiEh9WsQIR79Elpn8bW0v5l1WQIXU476rroStZCiPkwQgdU+eSrH8am586bWmcXy
VBZ4gRwti5OTekwUD5aKpAP/l3CNp2/LypVp88q+Yvjp4KNR9bZxMEDIGqOI1xpnragbsLJtmUFG
6GI0yWv6GBVIfULducQ5BL9X1OpP+MU/j8GFvpIFAgNc0pS4teCvZ9wxjWHQRpCqKG7OWCd/faBV
OMkZdnnE13m/QJ3F2eVRplAmQ+rNhDV6tHal5EQWKd45/xbgxJeSIBlGGKzHobrqgKzxBM4oz7o5
xQn+bO/6oDpChoBDDj5230t+3KBodTyy0BDl/onrZmF5aEs8P4mAWERmwZCAP4673DKVWQRxA7AP
QlOSeRNErbnzkqA1vcJ9hcvjd1N0FlfR1M8yxSS+Su4Mzc4oKfyc95AwlanQJbHOqS49BaXDto/f
pFvPHWFUiDfKUB0aKyLDyn8IbF1upBqqrh2wnpgT7OINte6GZd7iQICgSdMUoiyU1w0yTh8PAdU3
aN1aGys4bfqg7O6soE5jobu6omS748FsDHe7zJRyx/avrCxTwaDc0l5f7k9OnNY3eQXRegLeCsOB
VjpunUAHNTB0wjm54sS/eiN4qlkvSCCPH33FOGEW0JSU+2X1XSdJ9jVUhPd2Rh1cUlN2c5CIp+EA
sm2Q/Hloxu95/IfL7uUF1KyDMQ+fX7UZYAKtSjcokiK3IZ1xGEDTXWUKo/9wKhG0vYSVlE/Hp6a7
g6JoPvr3OGKqIuDW3usDVv0Pg1io9puskuAdNbgSfp8Hd/qn1jahqiLkmT8FSe1Lkf5KAYLYTQlT
0VpbC8NYb7LIMXGh0CL1bcin3pQOf6Kvfl/ouHHQe32wI32FIHjhyBOtNkqY5HiERGiuDNBT20xu
80LaVLM00KJDtF2Xq/BPgApwOxtj3Lh44klqeDUdiXreSDZWlRc9GpmKRDA1oBIFNh0MC587RpWR
fCg1rleSHiNTXyA8q5mTDoi/CyUcEHGD7qlFL0hhO6rKGFuYDikg+ezZ6gaS+FEcSY+7VRKaGEKe
DBFA6XaAh4bUIcW0IyyIEq5eY4M3U8JL2RWzv0eJfMaLg6JEGAX3Cl9KtojqsNi0rVE6Xq8GXCjh
cTwjEXaPyCIrAtXFrayxgBcrrRg1g86inkOm8XazecUcL/hFdmZDwzLMnXPSnaOk8/7aFRdg5UBT
nxVvUNl4UUY1vMnlCLgJ69p3KixsD8AKuoa1X+vyS0PuVkeKCZk5S2j0NypBRgyd9cRSlOBPh0f+
1XlbPx7pYV0hm+cxB06SfVBW3R+diT2Mhb1I1bOaR5Ua7lVILCQpIawTFSXb8deDeSXiehBpcV7Q
gC3c2HxlV9WrnMjy5Tt8CzQyUc6cjgqMiLrPc/3LU7taofza2y89J64uGY89/qi5PvAd5rt3sjSV
fpz0DpYnU3rPYTguQgPAE3Z2v+V01SmH+roAXvSwcjIMvrb1l7y3xY09Oen1FcZb041YbasUKiQt
N8mOmO0ROg1wZ7h8fy67ILy+gtEQujM8GZr3V7C7P8w1ASE3WIAahguzv/9NZ9zvnYSHOp0nxl29
apyNw3szCHfrfc6rqAxzlW7hSgl5QRqT2spHRCJUExdP8Ruc2JT/hyHgRrHps+W36ymHT9tLhSKn
r/vgjiLfUAYZzsqVwsvmh+r61WBkb9uhnZjI2GIcD47lzFYGVJNCHRY6ySq2KidiLGRQ1m61edWP
qiYuwQfsH3qXQl2AkADulcm9SZDLmfmQoOlr60Lkmwgf2XX+cRNmQXsPXy4iJLNTp7sVBfq9EzxQ
ISul+e5IUyj5RhTxyIA3encGJS5Cq1xjnZVTPi/pCCa9MGmExzCEIGa7dm70C5mF0jT7NHVMHvBC
q2DDRTJ2VYkHG9a7TS/K9GLbGh3vgI8r157fytiDAyyFHU4Z/pRJE8cctNPYy9BwSPpeY6DZbMuD
5MMo8xhzOE4tmEkxgEL/Ic3QFLwRtvm8FhQId5HkoA6DxPyAbFLQYfgCaSPcGujXx+UNPcS/wEAN
tMJUntdr936DJdm7yiCr4lf6BeevSd5vrYU/E+z4iBiC197WvMl120aHJebozEnbdZeQntQ+3nEA
P5Y3w6I/6Bnn4S6YTNKIzIaJwV+LVYvNbyhOmgsESi0AAQJbTAA3Tozi7LyVydAbmhcWaoL8ujFQ
8JTSbU4ba0roLzGbfUPscR3UFRboF7ZM34NnA35z+r40z7yXE05pWCVMP6bFtqO2zO8KOCjtusR3
+tWtKOzrQnt3Zzqr2ANN4nkzdUCAb+0ec+yim+5q8ZhDalj0RL3EDVkitn1U8j7YC8mfX/pQo1e4
mjmmOGJp3xFrDGHv4r5/5fY7Ao7BJasVVhZVn9iPxuYXtELwgDyf99ezhGSXU4WR5L5MXAdGE3GL
bqbCLC9ws2PAY7Pgxqm5hBq1DPrgVFZJ9V/pwWlREiZ4PsIj8QexkaFCeI95G04hJREhaj0lZV66
tC6CKujKH14FwjgPdgyp/n2LAdnNvTedyYHd4TnAVJ9iIh5FGvQ8vzf4FF3s3uxcc1vZqhjjlfe3
Xfah8Di9fG/YGI/6ToPe7GkrRzVyCH4nq+45VNvLYS9tXLxW8yq7LCp0e5z1e91dayIUe97SkS+q
r31LOzNSwQWkzyARe+gXAG5W6ytIgH3XxOuXtsah2QjIBJsSY/8dUqyZW0BppUCjngUHXm+zEW0t
iUAh5zO9D43L1xSlBmWsh2a6mmrTlzdP2FmjbYDyNDHrwuHAv9xG0jMAamTPwoJORDaThD/PzncJ
Tl3j+PIMIvhSxmvv4Wrze6qdHHsXM5trhj1Q/XLWAP46JY/zMBuoqcehHRbMf7dqjJAIUF48qLOw
rDKFltwnlN2yXjIIDIX32JBB13c4SCNEg6wu6kN/lCG94PYXd+METzSxOBTexi3MjOyzgq+b9kBc
3cGxC1AmTSo50NZL1K4njvY/Tnj9jPGKjCk/Fg0EmaWtkQ7QyQO42kYevUPWfh19j1XAMykAVh0Q
2DKKo0+MyOg7qRVi6ApSugFbyVVnpij4KMEuVLOGSx2ko8jiaxipVAaHocDhxb/wY+GgHTuAyWrq
6voEdSzfnEN5tyKBs+doJp/GPDOiOiapHuWQ6+Nk+gP+PRcyGpuAXzguKs/UiqB/rGE7e3MS1w/v
10mzee2cP+mgekCPrY2JjfRsGYY6TQ3B3wz1BZWM+6eJWKAlDV18JKKgub24ATKfvqCB1G7bw0V4
0wNEgyx36wzkO6zZzSAYQu3zwvTRAorq+tduFxndvM8un/xFZi64Ya9ToiDNx7n8XQsadS+IGcQN
VohnQpZWhDNuChG7ESxIYqdOf6g+vVxEOcXNaoXaued4mEKut5rkbkRXiNwhPMuyZ6P+Sx7ILG1v
0rQMqBGi7yStRFyMeL/15CkxCCIf+QxNziABlMleFEjIxI596vA0FQBqlr/yPx2Jr4UUp3T2dVYQ
HvKybPDd/nQQrkNzDWHn4bxObcW9TgfhkG4oKHiNOM9ZxjNlen1B5V7AnDf1XbIu/i/xv5Gj8cRK
UtYJBDfzgt7HMfWpQroOeleS1MdQ0DNc8m+kJWNcngd7QSekFv2IQWn1lU3s3Ss18nsdew94KXb+
8BnIju9cQ84ZqEyQGOaHnntOvUZitws9HrT8WEr2mOv5H9+hktm9idjndb9O4B8LuMUG3bsQZGkw
K+v0fCO4hZZ0hUfbdnlH+19SchY/oMAfXAee+CKXW3BfHCqEkZGxPe9btubW7r6IDenoNaBrZVnx
EliPdktx6MlnnyxkVOT4NI8CAGDYMGvDI6DT7s3h7rKswvwcliawvNmRvCHZ05IIqVALp7IsDlno
+i0U3ROWiCQ8u1meICMRMCP/DUgLceuY1M/cxKvyx/GQMqCUvqgZHYyr0iZZzhgTA5RDOOQxqfFM
xH/RYDh/CAsB7gm4dhE2gX4K3tuFWyDzyfjF+eHsh7C6swAoHeWEu8uiyEEkmI3OgfZFsPxBNBTl
xXt/EfjVYMtDJ+c+Nq001z4RsIRvgBnWQvL2VJq3P9KpHsq0hA3VD/r8CnkIljfRnO4OCXbWoIdD
0ZybWrMaxjbDV78ICF2wxBzhg+eMXysLXsuS0pLDnwx0zKe/Ou1SdPHUoAXywtjQiqewuEW4jp0u
MMOC3rZisbcKpt7OAjbNtB4e0f/GmHikCxL1BoAWfzCILyoUeG6qNJ9hEidh3b9RSiSNy6mPa/+Z
cQXc0rzRMs6ifaEnZuiHDPUImlTtOsV/biDB9aU2QEsrCLW05grN/Af3m75A7eBYc4dwypL8WKi2
edOWCetZgyg0t9XWlcUrQDP4oZqnTEnQK8WW5a2Eekt/G5H8FyYRYYnNd1Xr5Ub5VCG3QFwsN6Qk
4besZPxQgA4A2+c9uI1R9T3BY/2XhoYTFSQvvlre14Q/K+6qWQPrhzvProh7W+Ve6rOzH7lFmcqS
eF6w1ZkGF47we1Wpled91yEJ9U58hOXfqvF1qz3xXsOT8nPQp5/jL853iYTQfBA0Ru4Y6Kf3hu33
PueAoJlkah/6dJHvxvd7mlfSeQqzXS0EBPpu4tWscld4zW12RohDbrfP1E0JoC980bYexPoaE7GB
XpKAKHweHM6Edm5zM+JU/Lu2gM71Xu2iKXgLHV6ku/BMp+yiDcb6TAXhnhSqWzaisV/d3hkjiJQp
X1LL2i6VONbounuzztBHGKreefh9LWX1p1RdEMayHKuY0+yOjEer80poHel4kdj8m+iem3QojOaO
z+TCJS+bqTFKiXMS/9NjtH9NKmHTT/6rVYW6s17OsUhFz4cUBmFeI8nRBeOMGW40rwXYDQO2xX0V
Bqg5tXWVe4+sO5Gj0LK4KqtbJyaYf6JBBeMh0Tt8CUpstgfxmzcQH+ruabCuwsWs2sQID2IcZQGZ
pjNH7Y3fCj35XUwhY0iw29q9ayxjMsqiLgBnY/EeZj+R1RimtR/PhgkfOxW/68hN+ZRKobEdFj0d
Xi0v/RDiFJwkpXDlBxyA0lNdf2iWvuwDiCoHM5j8g1juWDDbqQ6+blNaRCu+OrFDlvoVegYyM3+k
/ztmP1OPfk1jezTPTdAmoU+zFTdvzdhFDkPGklQLBk8j+YLSFX040FgY7MZU6nCubZwnsdFW2uys
8rMbTYDXXK604+P/M16c4SoI3AQ60ApdHK6RJJSzBAUR5o/fmoZ+CEfkx5n8I4EBY5hEyuJdjKdI
e/2aOddWgU+/TCxRG5RVVFoOnyNNrsV75V9PfZT47LoRZj4ZrivkkDWjtqHpTQtzLqwXj3zyFJBs
GCEvi9tRXpk0O0HqLaUlr4kNEPaXgTxDLWBgkNfStodAGsOC7RPlTC1E75Xw6+RfGJBdPGN7yb7H
g7q6tpEMCwNw20Nh27Vj9ddQl1OPSULEy7NPFt13AMo9Dxe7PSTaRslS5hWm8sU/bTtHL1YH7U8P
XuXsr9vXS9WoF8tJ/XxyryCKggS37ex6Oe8Ng7X00/hWQTzJjLNubg+TWIWSsFiY82aBktsRCnR8
f59lbVdRmd363fHuQojix5u8p6FHwR0QtosOEktCcibk75rhTUs9zLq1+82+RXrZOERE4/4aTPPJ
eBc9Es89VoNj/xzrdR34ItQIraQjykru9qV0+hU0T1yINqvOczqjdYIZinUQ+j4FFv5JCfQMZ7ps
+tdGaZmifFhbxq81Fv3CQRmFyYD8IWPM1nwflS+L8cSodGv6aG+EmeCxkdARRXMr5NKmgAwLtwUX
yFDw7UhF2fje70N2ZM1771sfs4xm0sKqDruDynKzHnLy7kR7vTjLxJgDGj2n1/qlobyZ8mcsSRZ6
Nf3YQ/8sR22vAP05FQmAwPK1S1FZcO1OTvuWy+vyOBRsccDSF4TmF0fwiOLVkO6TgHsRX/ZRjRd8
aBLBAbX4wBVVoWxfbHSXJmSUoH4+YQyT/Uw4JkplYUmmrfsch83sIv8tRqUWVW9fGf31vCtmdj8H
zEY0dsLV6FAKezIInCdm2M3K6EC/6scBQNsEr/p5uM4+xGkcEfJnTdf2lTHzNDU1YH7X87hM0D4l
yhdBlusJzkoU+XLO/EdY6ilQ3SlDzDwMYhGizoIWeNkrlKuOOl7CaesSel5Nxs0NJIQk3awh/hM6
no+irvYEr7RCvqrpOPu3HGvtt8mJ6KmF6fSLFanS+K1iXVVirfGt5d9Ttrx9yv0aBrpVgI+EdDtT
cDz1/gTaDp1LhcRotwH0+m8dzh7XI/uxNBTHZRY4XTI/oFMJBegIEj/Njq9j3FBoLNyghG2/Dx0T
BR8BSVzNMPXXZjfuaOHj0r00R8PwoweoLzvt6MzJGeiM9VpJJFH25CGT1hk57l+3XOupC1AkiXM/
//mpvGdKDgFULnxJpsL8exJNcU4Ow/iiB5BsIGw2+ou8pcuihY+tgWfcA282DkFlS6iSkMIBLrto
ZQDNKMHHAaTbx0IDofrh3PmqED8OT7+hXrmBKg30FP3q4kL+9bpjlnAMf+GUfiWNtFAZK1a0iT8x
8YOlRWXo67hfaFtyvh4/6ker50EOpnwBbhwgE3bEUKdUBVnduoq8TlfUcUmQoAYGXOeTWyg6vrxh
7NolB6nlQ7M5VMsA6BvpAdsixI6QehsshDCQKbiXYtYyYvJRzOf/l5Au4NzxEjwbR1sKXkWuSmxk
WwXGOQ5TLtcQwdh1ozKmAGVsuIXq2r4p0echLd/sliojKn+7aX68arIhfff8g0MGCBvWnM7NtMDi
+PhArDlTvRMT5ZM0u0QT8a8GvrETxJhq0E1cVvnObcRGxsEja5rp1Xa7/zr4bDvan5OYPPs4LMak
fSiTDrnKcD+2iQVWc03fiXrjKlSzvgnH7WkNlv0QujX1TKj59oxsTDSnFOQXV6xV9t0opi3NP+0R
ic16i2LqKQZi97UMXlYjHHZ0LvTMCeh0WiFgtHDo+5n1IpLXz8xlqTR8lCMQsJgUBlJqQPPu3Y5N
Zf7rAh07muyKUJ8mwD7pzVFxmqG/xcpFiM7++QROQa9WYXL8REwFNZkZYRjcjsTcOTY+E1wanyAj
cMgZ6+OsJLc3Qc8JUoWbkF91FyAPLH6s/DKhWbL6e6nB7kQFvNyC+uk7883eumef+ULCBqbD3txg
1dYERfdzW9cPQBsZDBFF1uiXagYCuh2cH/BqF3jua11dUf4bl1jNwuSHcq77a346J7xJKJ0GnK1K
9+ZdGv1hZCD87JX7qwDu/rq21PvbgNEjIMttiE5J2LIJtTT3QzSiSeJuvDwqjzFzxe7/xYHvIc8A
wPn208cWiCzgJObdgnu1xbTlE577mDZbzdmFJtnLLb6hpdDezBnKaNqE3fcJuzMKjBvsDHfqTSyE
AWDqZffgQvmgcK2O6molkTeoTAqswie/Bgs7mq/Se5jliSXzYMhC3+EQaDPC/SH1WizGlJ/aj9mA
VvcatlM743NHhOy6kXD080HRUJGSf9lkm/yiWW+AcOD5pTdy7N8o4wzw+2Z+1nj4yfPlADOM209/
XMy5Mgc8srCr54XM7dNK1hUaLwVj8+QorN+JluyY7MN1Bgv5tmWeKFEp1HYiILliXw9q3o6DLbEt
KExANRO3hqC4GLhydkApX4lXLfErXYO66kPkH4aBMjpRlq3/uoz09PEYKV4MG94XC4R3SzcLjnz7
SR8AWc3FR5qg+o3+igmMsR3Abtkf2mNMOzq3EpElVDsJvIICN9jAE/qI9knI9by0F0LTktnNcAM8
hmZxY3SdO2HKq3wMPTy/vvWABLSBPRuZyPrDUL74Ym/fPNPmzE/xJLFKuQYUC01YJVD6oRW5TyrJ
OsiJnQaBk0jAZW2bmrfATrG3m52G+31avWxvgkFdaQW+huP+jlrqvAJXLQ7VwQRQpgHBOiUtjT5h
fapejVgsLEH3Go4ATdcyIqwdYdAznrsBiyrbIbBL3Ci6p1PVW+TM/3WOGEwPJCPAdg1cTD2lL+UR
ZWg6s3dt8+B5MH/c5X9w9vjpXs+fNR6uUO5GcJKklHs5ZzDurFRYtNM1ztwtYrywdhmYDD7sAs8x
lh0IqHQWxNh2QK5hxvUk5iFRtpb4f8xhJiduydArHCEw3w/N/PvefdRfOey07//99I39Ms65L3eU
kOp7S/6/Tfb161+Pc9oOhm25zb7ZxQjP29A9BKMAlLJVcwJ4qHbYiTzYBdfyBGlaNJHQ+f67GiBa
IlCMoOKz6uoTxUPcPwcL3z/Y3j4IsHFDl9qOs5Se5TSQeWd+FCsHtRDicvsLZ+bnXKnSPhkS+POs
nkVGdoC8FUoTAuY6WaLsjn56VrizFxsf8eOzWz0vIYvcKhK1aSCaJhNwvdBcLWh+ZaZH7o6T9o+Z
xfkJaQ8E3aWClfcCl581YbJzJGa10kYaunDJxFPOHSgbwNNIJp0qsH3Cd9SUnOy460l8oYBoSsp4
Ig7GuFbFSYVnIAksPHkrUFjyDEpllXIgHqipecr8tZgKOuYE8JAUe5j8qhHFuiYLy68A9Ai1aUgt
XdMgQ5fPI1Y4z+5KpIgSbf12/lO/voFNVbB6ZJvbHaxrQ1KUnuOMFDrwxnaoMeuNSRkH//s8GTvI
1bUVd6CmAZD1fg3jl5626v4Ix5ffYVuOBAj2csP9i3n7nv4xVnZWPR6pHIEP9ofeazF80pEkk9CT
upQEah9Fe1vWyAMJ6O7ZTUSy3zSv5pntnNGykVhEYObpUO4FYbBKsWYjf8P2OjUDep0r9+QlANsO
6A1D55DmvYQhhHjO2DAU0wyAORFyZkZXpxN52SUaddms8Yl9VEcmCbTHT3T9EgXiMvmYCkIJRQVe
bW35JUNAhu8K3CB9JZ5VM0QvlEj5PG1H6leysVMww2CgGHntM8yp32xEQ7Z7TtjDeF+Hde1A5YB0
HByG6SFawe1iw55YofSsA7Tm75wEyoD6N4X18/q6id9PWHlvE++G3TMVFNcjdhcB9UUGxcg6E56e
YIJBpbEAHEztqRkPglgF4ZgZBKzFenYQL/YoQL3DZ3np03zXW2dIm01Jqd4jU7kjGodNQoTebTqr
9L8qVwuTHV3/7lL6+xto2VWUjInw51lliABSgHkMKXKp1VJ3xb4bvxqBK8r0wU+JQoav+wqAAejz
Z1SnbaePVfvwVWP82khFCZY/OaVcIwOxdWS/svJ51UbH/hWEOW5Cs54VgMbBQxLMaQbseXhtxpbe
dvPok5t73LbP4FBs8MgviUc+QZUxobepOsVDOnSECH9eCDO1iueqgCKnyGxfgWRqq9mrlgTZW/Vp
ym20D1lcftyrO2JRMkTSDpgO1aO7dS/0OEp9QQ5EH29+G+vV0Fs8AHK5ZDsU5nsYkhwDm8vPOPbF
C6c7fOLVqanCYOhjDFANe1h/R+vmkrasyEvOLlZ4NavtHHS7m8VFfeEgRnHCbG5s+DFiboX6pPYy
BQ2Aalt8mydwjCeuJj8sGTnNlsit26VwPuSVeGMOWLT5e8KeOScc//qyONe50vMNAhnnxKQtM8va
GLQoRBFcYrErfHZPWl4uHwuIXAMhfFVvxP86uGtfHoYAM5D1QZcEoAqtapw6gLgaG8nIF9vKXs/2
H8NZiRt69CvKlizPylohnsAgJ1qwX9Mwz0XZknrmpkmacqJ18Aqnb/rx8XmKMoepw5dyl848McMh
qq5U6Z36ihM8Gj0btaR1EEW/jZ5tq0MCsYXlTjDlqaG+xmrHPIHcxk/i9Nwy2R5Y3MSWlP84muD2
IZQHpnJUj3S2jSNEYSzxSJ5C9A+BpdM5Qw2+IujjfzrkgdCKaUyI3bnyBo131gkiiIsxABauB/qI
hPfyHyQ+fmL+b8nUOuLxLsX/kPlkXOKKLuUzr4Sd7LbdgzMTHNgtBps1Lbqb7mNsi+mXeXNLbshW
YX1+Ln2/T7fr+t2ws0KdM6KdZWRiryDQdxNfez2QVA5hQxaLLtgyOoXTSH/r3oq2ropxLsmZr6s7
5YaoT5GOZy81jnNpr7j+4JuJzvuoTUA48LmQ31jc+Idf+hQJhYiTLGOrgyhHpC1mJCXF01pt7Gkp
mNVwsE4XfRPurFfWHJjmIiJsEOVwIIny89zSomP3oQmm2k8BkdR1isPaKiYRtlh1PqF2Wa59of+D
nYlarJXFFegtMkyHgqqM/Dhc8m6Rv3jDFBRzoI0kA19++9/vEi38kFl8AWH/Et2KVFobIkFsnS5n
Gz0T+BaAFQLYUczZ+PUlA6f528MbQjJCWZXvR3EfC1P6v9VSTFpGZAqwKD1f4H7mf7dQjifhYObs
bbd3UB/BqFE2w5Em+3DI9h2VQz63/Kgb1tf2If6IisOSbIGXfvKhVXKBTuVGis6q2uIE75LrEZXD
VW/PBPKgsISaxQoa13FoegUCPrfedhy1rwDLYZQbB8sPZEVWXEXYUDBOVdQQ6HqJqnoqDvV5+BPl
b/vNfTgKdV2GXS2UhxMnbnQbaFFC/Ecda1FEDXiD2E8yMs9ruv1C+XLPU1FpcDGK+WkG96P1jTDn
rZwmmaEkg29qXY30dOTEa5TWWkWckqM2FuQi0Bp9sqnhxGZ7bV98ijHBPyarlkdVk+g1Z8NOsgNw
6oz3X1sdytraZm8tqFMdzASTw2JcSlipBi2difHqpW6nk1zR70XjUI9x/OqbzA0huNZRAvWfQxer
9S/ER5ls1HxBgERcgwxoPhzlLjcEGVAc2flKLza1rOVoTYsbWDfgw7ktTyJwLbu3M+Vhbln2sTLS
Q3gQP0XO2AJQ1NVi8bJx/AEde9ue+bRVJiu655RLciQZAfR1ec+27K8XyQaCSJ1l9EKA7ZSm94j3
XeCBJ++RyAicRAx45h0gW5x2se1kgALEifIpHuSasuTs17Gm6S87SsZh14RYluPXluPkAkA1OFh6
gtOa27z865XRaHJZk/nn1d3oHLBgdDBESEipeKqIrY+M1z/qMB4PE68158EWrZkVhk8/hG9ic/JC
gvRVpCpm6yEKtXUGmlvcsltH9koGcf0QVKYkgySAK280Trt8Kp+WAOnAuxDca7MN588JZINlN87U
J8LFSFflyKq8VfgNXM7NSxe3wl9f6hFdFRPpRTqnXZOPN1HJx+OiNcxgJm0S5aWR42+Ca3Lm71Ca
OH/7sNVJ3906HuKmjxDfz2o0rQxnteakg/MuZnaMdp1phbw2GNAHOZAzjkykMPiCaveGVYEHoO1R
bS1GXSLRDIW7yCDkum+kt9PW7HRiyJN0w2fsRkZgBD1nsOw1JcPe500EwMW11QAqhONGHFjoMvoj
Bac+dfuIfalipSnLHJFp1qo9UIKcHFIX/1Tz241Lf1vZ4j1SKX2CX8rMloiHXIj0UP8UacyQcG2o
lifUjxxXSN/CWqZrRGs4Q1xBC1EEevXIeLhXceL/+C+8P2CLgUFhm6BjuhUI43tmydw7Q+H1SZkg
cxWz/WxHhxpuTnayEdAsmU8pSwyfrvWZs9mQkGlnCec+E9EQmtX5uy/2arIQG/FCOVUV+oQ+onz/
qOmy9gILSrs9zb2b41NK1UIsecmQJztGLaLNK+KSHkeQcsGORUUvGAzZWWn4+g0HRHWOGu3BmLqG
1Zb205QbiT3QT0Dwkkd7BC5S1cjP+y9cnBXJ+UqboY8Ytp/JoigYy2ewcKgX8Gp8PD3KkEnKY06j
GxiZuFb721Hs5Mxn1sXbqx8WWflDM6SRBnB8mLY1HC20NtzHQ5Aobp6grfyHNFMQn1qxP7E8+oQC
+ejWje1UzKug3GBN65z26JgoLZ87d69feTSRSH9XelwzmLIvev4MsbWrcB73nsKU5G8Afx5XwrS7
8RdtKZFuYXzAUjNHf9AXr9gdh1sVi0pJ9MnFa1UdbwEuqElbhSnPDb7YS58z61ClksB3Rmn7b6J5
wdOiiPif2lCCnZLecniau/xxt7NP27gTzaScLM3gzqL/nE2NqdBJjLc4Xm26F4G0bkmRjqYXctaY
yT2MGciIQr2TOIITwnuFJiLcdaoXGs8lU46nD9dSVrBVeUKLbJCKaqpcBBODvnRDb3qWBE/hr9xh
8k2ORFiJj3JgLUd2zpsvcMSHKhzn57h4MQdtd4m+r+B4J0EMkCrFaYv4Ja294HUw7CqoB8mQ1yP7
PjbQHTNQvU9mCzxvaXrS1ewnZZzP04DOvjOkPlvWHfd6Kco3WQ+K7K19M+lVZcsETVYee3eMsBjW
kyaqZ92Xaig2TgqBGqKs8etPoj/m4lDKDmM3pXFLvqvG/uyz1LQQ6kn06fMg7lOLQMBuU1ve0mwQ
dU94fzEPmRaS2dhQAEroD2npLCzwIOLJdngzaUDX+kdqFnNF1A6vwmh4iJmF6VSdPZtoXokCXwH0
qA55MOJHk4gEX8e+WGpT3JYkuSko016QplhrfxVggVjLMQDE8bno3rCSusuyEKyVTHcG8HprkX8g
YSKYH/UnzakotpKKJsULsDTJhF7pCAPq5dXvQjVaNgv6Fo+iBG7ikxBVJzFcEcKEoau2+Y+UDn1B
GyGJJLuvV+JuhfJf9UF8LcUmBeTuFH6VMVnuZhYfm4qqG8eC7vCnB7e3VZAuzpsahBoa6z/YsUUA
4Chcm7+Muiq/+Dakeqt4+WTYIr43e5ZCRE1zU/52SvpNAwa25PyBrqFCRb0DTHAgYsgGpzStfOqE
kNLYRlJ0TM9WPBKY3qXsJpMwnRws7s1z41X88mwrFi7hAm869sJE5Lt8MDQUsXDrrjq30J0CbDt/
DDnwONRi5Tvdj/4cDS+MY/pecRU6u/66EaBMUabEpKsUkjdRIaNJcChxl0CtZDtivKmSfCxfd1TU
CYvYO52n1a0H1zmDZXYU/n4KRfdZtwd5UyQ0XdYK3w/waNU7q8tVrbnCDqOR9+iZq8+fXD9lPjmR
7PyyHaLfRy+TZjEm0GWbjKV/fmJMKP9o2ujmCVsLB6AoddRUTPYjZOE8OsigIORJozvDt+Ko4Ibl
/ug4LSKMPTFMlb4NuTH5uyBb3UFJ4QQQH+5OdgtRLVpyd6rexlAp2d3CzZrl2vizbmhSKuSlMzU0
dO1nuTLIWMYnPv3ktz7ou387Ed7JhuSKdKI170WnNzBA3klEX4EGLsvwIOYcN1HunMY4Riz0N7l1
u8Lomnt2xuocrVDmM/jr4SIFaJETJkG6wJvGiiJjZzARzehTQL3GOWG7sVfr4YlNWlQVaDI75AvZ
INojWIJmpGTeN1Kr25gFeEViPKzLfAEN3agEQe3/Uh3nqtlGuZGifYoosjsjV1ID8taQYJY8RCW5
Fm9LKcwevjR0gqrRNmjyDabEOg3PeKq4lo7jGFsRyU/dlx3bD+l4BK3JK0AKLDuKxXCh2mo+HUB0
168FUICLUZj4axd0NgfOzRQRHjP4Erp5yPfSpyQHuK0mYkahFKSAi78YxN6yqlmYqSGWbnosbEtS
0Bwj1/VdPCK/PNxSf3ThQs83JzKaOEnQe1V8Y06vQLYR4QjaqX/gQYiBQjBBuGuZVDYV10ccIsOD
DR4vjLifK9hYof1LxEdtQpkuHPtF9x8aZP2QJE9fDi0L0lBmTz1T9niu2h//a3/qbL6yGvzB4dKr
MvFfSzIP7OsDz+cVDLUyCygXOnoFdOCfINelDz517QamfeWDzYWbPVcdJP+ckHUX3Q0pYX+hYYvq
7uokUrIZPe38/I44siLIBAcy8xTuDjjOA9sdK4K45AzOzwQbUDF/cY/4B2FCbDyx2fU8nEA3M3fF
0mpeV91T9zckYjOAnmWUo1P4dIV/NoVrkjhZKQDtBCjFve0scx7CJe/BCwBieXdUDroeefEGAG5c
DcpFInSqnUR59LtyJKh+S7Z9uG2U8hzPcqZuvELPuF3jtGq2jLAfBes9/cNl5245VO74NuPYDvvd
aPIDoa5tmK78KAk4G7OT20PkTbOc2e+kfBXFNLFiA9xTLB+xdf+TuRwrvVKvJC5eiFGrbfG10TeS
GuR2MjK5O/ZA/I9JE01VjJ/jo2hER3HiB7AUN1G9TzjMNChXTHi6DfQ6azGhHockXcqFW6Lg7cEe
X9XhsIn/qf7bZ06N3qzuEL52GBC1p4x0f+l75aFPYMI1ThTr7/Vo9CLPhVihp30foPf/4bB0TonJ
XrT1pTDQrPx1Bkg8QI0O2pPQ4xMLXivKvkvPzmjIeIZoKkFYOST4M+kXNOuwoqQGxo3FhvjrQJIX
3l6hNkQ3dG6wYE8Qmb4q7fwRPJm3q5ewH2Q8m4AYTicCme9vGTGu5sdJmvg3WkffiWTk/94aTDcW
cc7a/BTSCVe4TLVwkcv8/Xub1OtDefnpp+Rj4gZW/6JXDKJGtPLGWCRfteQLAHXcForBh6inuixf
sgIMoRsRMtsSsPiN4iNj7VjP7K/bcxD3dGoBuahWP2GUCNuKDcsQjlc9DgH+BXPQtDpn6wDh8+IP
U7O6hUZYYqfIrWAcWmJuQLNV8xZsmsUBiYzUo/1nx7w2AjUaQ4Rvr3mfBKgnh1aUuB2/bqizYY0v
lQn40vBXxGXFJU/QaKdZrhC99T8z0AmWl3AF05enm31gYTRjJ5MB2eyHArlYDeDeiwj/yCPxgHZL
oZNYFZW9oDEie8B5m0MZAhtuKCeYVmtu2MWj6a8D4juvDNDuic5D3rHc2L/M131ndVE6XTJGTYAw
wmIahTQWgdqN3+MehxtxbEyHII6W/K7VaKjKnlPp8wqvXCO9+Flv/KqHGrEUjztMU5QLX0QiSVBd
0ycVUdRqRoITBy2d/tsjw55AD2dZ59VD8mIrro8gI0jpXXRf11V5YPXxlRMPgANLcFSDpNWXZYu7
d5wwvQ4+5gtmkv5XjPkfdQkuTDhxeny+wwiB1CCc8kbCtxp8TZOx7/jgBrL5xktmy6WuYNFtyY4S
pXgVz5TyN1Uzlwzt/qoXp7GbBTy9c9ESIUPyKQFskcUMsDz8asbe17CqEs+C6vESzDB8B2fB5tTO
GkY9dQhC8pw0yxPWEC9o0wLzs1hTW97YT/5crgxWsvKoTw+wd3MrARjeYYdu4jXlBh/uR11WAlo0
dzvTYroaL0TOfxAgeFKhlRFteIMH4ZsXB4+OtD7hWV8mKw3xuS+tuAvKjXaXvzkeNxh4QTUpjAFS
QhWQVBTtEZazyXctKqSSr0BMlKhzLg7jiiN3JW95Qw42Kh24VSukaNBVukDFBFnSaadD2rnBZ63s
7JJmwF8osm9tLV7hSHdSTRaG7S2gE3En0OkISDeyNiUFaCN/8mivQ1/FmNWZskrC1tHv5sy21ewX
eKx8Axb9iPOvu0Ex49C2C2//z9B2G9etdx5zhEMVHjq1LQacCzesblXs83OyPw23G9OgtLdXOfHM
7MIpHDd0LtK0u6XdITYQhRRR9fXt/wh80+Y04DYesOm94mxG1tfhtnrXlDCVPknbRPRhUE8AdAxs
qn1IZrvVmzfZC6tdoZt8inD69yaeucwEeJemhoEsZASWK6w/pOH7XwN2NPxZdG07pMmKG2Qb2ljM
ePJovoxBxBmPEErqZAYRoGmv57/etwGVYr5yY1fm+VEMmK79gjLc+beF/GtRKw05lABVJkekGNXD
JBjCrrCmZ9O/Gc6o6bZIhI1v97kyE/6iAPtFRoSkOtYY4l7tp3zgF8ayT8/rXikMdbieT6/xITYe
1J4vbfpRJdITw0u5EtoPlnElFoDivLbx6eq7hauh5c4FqHFb4by4dTqEPwgWXzxjA9IHShbnGq41
VoMLtruJiU3U7DVpDX7GrdRX347NajbdyuHpi+mG8DeG703gnkiLgkw9CAoxIxlIa0bQxl0Kz+Fn
yzPVj8kkfqA/BcjmyU3wfcmB9UP1rxmAVlXZ8bsyDxVhylGWeRcmxXtPWlfZtvMywjy2OrhrlTdc
Z/yku1cHb5t9aobzSPDfKCTm9VSRP3jf+BSMfJxaqbDjbb2IzzLfDqKwA//Rp52Fzpq9RTLODR1l
I1HrmnYsOHvkm5mYL46kUqrCjwXdwG7D4knJx1edZrq0fC6pW46ERBaKyzPuSTny+nBZSe5sAH2y
XZK9LxFDzQZjqzbxDQGpBFi7FMi400np4FxkcsZ1E9pSliq1GVVUf3mi4LYNMZp337TAaDgKmWNd
4iFC3tB8bGpPEN8bq6JOY/QVtqAfy2rW2i4sYmqpq8IXdK3SBhxkT9vB7Rawq69WVE/hieyntu5S
VrLvEkAd55XL2LLmqd9BXFIAN/ggM51cSC6H3a3baTOLfX6cixoLv9yc1+8DzCuw5bOK1JreMrHl
HIwjcitWa8K/Jz3WcKFhY/FQdX/N3zp1E/rEzWcB5D+V1rwG3u9xYIFOqDar4V+cobOPW8EKJi2Z
YMha2swzLWO4s9UhbIf+aljiXHobEtA7cRY4FoY702VFO/T3EF1GMbpSX9DzOSuBdvQnJi8VXoVe
dCpf55fvl/PqkphRqsrH3zYErZgNfkVoJhHQOC3Hh581JoMG0GrumSS6OJ4Y4r8760ndoeTP8hBq
YkbuFMc75uruR2P58IRTeY6I6reLFT/W40lr1nbUNaqtBPjrJLD6atPOvemriC8OelaGPdplnUsu
aBu8RdGN5xGl0cEZPJu52oNTU/T1OyEFURH2pL0gtmyolE2MSiG37fJBi+MaFE5qYOH8k4dacxWO
qqU+HHCM1S+8tuqqCdh3rw+iHGellTQqVA9wJ8Jeti0hUGbLE0QeQOAjWQxE5sT0ZiQNqAYG37le
xyhDr0HbLsvMIYBRdZJR/kbbmITKyUpuXKvORbWoBRaRuXiCHndql6re6p9t7hzKEVc1PadGbGM8
rIdESOI9W+iYf6VWFfnJ4dEJx3l7uMkG+LESjFxd4A3EZPDGyn464nfBUKHh0WMV9pmyDO5BCblQ
vzUyDhKwFoW9tXYqmzeSSoH14gASzfgy69c3/Z47yVe3IPocOIdQAyl7CdIuS+BvMIbumLanF3tP
2Unp692Q7u9SzZFN0sE8QJqZ8F884oYf6xQEwXWFc4IWKiHRv5Nh9mI6wO3x5ZQNKWjR/y2Uhseo
HgcNhWpHYEGJ9KFP9bvy1rWuMd7fh5uQGzunvOF/nfQbcwMXoC6sCrmYP6pK19GC46skY12PoOCc
T2NMZ/S99r1HnqrB397D/i5GWN0AvJBJnqsxszREz1O2XlyRpnDswqnILtSRgL+4P5QOKd0pHmnA
Vy1Tcud4RyWhrW834ysM3XkljyXxT0e0F4ysqEcfrhOxNmA4tHy/XTdik2Duc/ZDUQQaQqcVsXZp
5SlFEGhSqzWPibV722WttwvNtgk9+D+OtpXse7YkD3NzqbFy9BG0mwlx2Bh5DTp+QZ1p+rqU3VJi
0gkMOzrUeNTZuyzjrXQoyq+P7/a5SguLcM5Oih4OeyEuyFo9BheVKZtKGq4pnJ9ETg0eXmwe5gzE
mPy7RMF9BlTbFPvLWC10fcO8Slyy+gdmXVnBWvBpgvvVDrD2iB+RKAA+BQNMnfZQqg5at8PHdEzE
h1WwQe6Uc+P+lxEbGMvICNB5V/t7+cnN2Wn7MTapFV3HgIGkN0cD9B3FP+uT1AIXBCLaA/Dcfsyh
iJfGXPZlGRi/fiD/bKFyOlGjgiqf69sf3J/j6m7xU8qfZepxuU58Kb0mTD2PHK2iklf/fXpTNv2I
nhA9bVWYDqym07qT0HpkZzC92MYIUtzGch3faA2l3Np5LoB2kO8LLyevdh6GFJ1qrkPDDFRGfY7a
axMhiyvdmEkDoSVnXIALXME0vr/R/9mwB/F3wDhucj+2St9OO+BHtQbpQtsnh9mRLpXyCdJR91ih
pLZL1B2SYWJqbC4vzRpW+gm40k8Gfjq39Oj+ux3tp0qlJzoKBgsshiIkWXYkYfEOiGaeJolDeco/
N5+ybFcwSILZvYPWjbwlCheOSwrti8ZLa2eoyPUZ7q+VxK2Wzix9WmdzPbY6V2+j9Mw838qONU1C
qvuA7bcC3WV07jS8+cOWZlgaMTIf9GhQYOy5Pyg+lye4ZfnKrzuT0NBSW4dpvqwc1/et+R8Csxco
GNnqx7ru8Qnvt+sCI1oMJcAl6XjAza0svD24ufjX9A9ymwD5pzZVGSucctORSeO/dVRrGWTWfVhD
2LzJ/jjFOiGj/lEmIraGeePWk+suoM0fh4xuRfrDAhFPZn1cHNYfUcIom9zxj+ljAeunjQYnmriS
I+i6ir0a6toNlG3YjY74nuSRkLSEPAmX8LoQYa9I2hs+5AoZOGFuaVpFQQxwuxuL6laQ54nSte5H
52Fuo5yW9RzjXxNTS65ZEjywHIKs8nhtev4i9In+vCHBYx30XvT79snhnw1SdSLs214Suu0xGRlk
5UWdMwVYYiIlaFL4GJglLO2rkk68W47YrLyd//wagYGQr0I4pDZlhNQ/A1eoS9O3WmLsiG6YW7TX
16l9DW9dquEkM121ZnwT5UmUdXJKMtU8WaKwxoOz9hnndXK2Mqa+6tCNP01qYN0jiz0I4lyLn5Uy
Uh/jPNkwS93pcqr5npAt2liie3+6+o2I7a/N0An8k+5HsejkEwb9YsFrKySyGzs9C28d230PpNxf
J4hmiCCQapU7IJklwOdacOAR9nJeAOR9MggT568MR+8DsAaMyvOJQXaLfUSPuSHS9nsTUYZ0HOvT
5mGp6CSNxvI04V2Ef5Zo41/mOgew26Q2yAIiUcmGivz1H2NH6GfhxshdShx6ypRucsSfE7NoTuyj
7p6ImBdHo+Bhizr7fKSWdQjD2CiI3sSiLsTr5WL+1zkSGcwfSnpCFjyVoSzNTAKJiq8EyWuUch/j
MPkvK5x9HC9zqTIK8267P4GvDXjF+n8mZklDaC3C2bsEZ7+h0DJnHIOwdUc+T13gXcuWyj9Xpquj
X7n967FAqCf+niYXpQSD+/yabn3J7Za5sWGYXmj/CxQuOjGcHBA3ZK++EKl7cj0SlFP/+3BF6j75
MOQHmRWyKQ6nQiEm9n38QRAndANwez37Sx1HHNgLwEtHQDo3plpfaUHa10s2s73Cv1FR9l7LISj+
sl8y/vo6p9K9Xnpj7Tq8/ozIMkSb+bxjzKoOXmdQka8BwVi9x3U6z6JvkNXXgRb0B6uzGOzG2IAb
dP89Snl22H2DTWBpw1hdU0QM3scOdzm8pqRAO6o4qmRVTnYSBHVQwSyMAtA8mlZDay0yLXc5gfop
c9MJLYsOJmVtLUS/hxaFJQaKKsq23CcrYeJiGwetn/Nc6tKUPDNYMvJW3UiBHY3E6eBItNDyEVIQ
vdATlpfg/lefAjxcxp6pnzYuxKrQUNqctWmwoHbBIA78pb8jU8jHl3BFi16xTel2h/HHtUCpEYLb
VVxV3GLaf99rCZHlr3UuXYq7ODp4ezIFZzzQmVqv0cnnxqQA3wmZW7y+hXrQ1R4h71AJ0YYIzawm
NAD0ZR4qnYJSGdAPll1yqseRw7rycecIPYjEq/s6oBpSuuX6bGC2hcH9IrN+52qCC7yrQeZCFSdX
xPZp4Ewl+pZ6mxQ47d7N6cSFalKZf00egJUU/RWPhf2lg2SoerEv7en3KRxK19n9+HTPjyTGm1WD
+M241mdBhnu5HaGMOk94UnLZMAAMZGOWi7BNUUW5cbb7JxB6qxqEvnAaqI3A22lOqbpUWUhpUJN4
UZBZ0oH7fYokJj6uXiMkVUxxDCd2DvrihmjH3KzhT7vy7VXjr1yUcxcdmeY3WJRebcKmvhucjL0x
JZGl/bCb0KyZovbOilBKHiEHJOBhnDVluTQBEiuQMoZqkcW+Po0+yJFh0xSlsSowN7izyZ59bpax
BTSvWyoo6JEr3MBggtMRRJ7/e32SrYHSgW98LK8EMGatxMXVJHzB5iT9pruMzibu5p4JtzIvurMh
o0hxLA/rB8EN3ruxbDH7dwhRhFRP3otZvBoDsd/yoX0fUHa/56V8XDbL+b4pocODTCj9womiK4Dt
9vXOW3tqAIrZpMMuPJexgikTDYbAeKc7DYKgjILsiXK+DrslKMTMt5cat265p5ltzGrO7CPREyr4
EJWulzYye/sRNY+HnqXSOwCjmXDyMBZLzaVa+6nIY6ryl2kEnnuJ65eMzGJQ6ePiG+rvOiyX5dgO
OZwtmz3evqe6XPcMwNVsMjo5BMYDG/6fCXfnrT3PR+XIVqUFL09EB0IqgtZmJ8GZAAWpbHmpWx2E
XESrrpPZU5WbKNwSRkAPTd7ujx4ABYPVAVJTS8MkidbFu5k2ecohYB2esSHA3/JWNlAqsB5kiqmJ
euRcwyjsItPuFu01dbOoCrwj+5i/KQCC89icgE9jX/Ze3VIYzo2K19sZgjF9xPP1Tb0rFh4N49pr
5ECZAunS41LyUy9SZPlaKKzCEy8apm4VAndrQrStE3JAO1epQxeu1tqV39iv/9Mod91YFvW4W45r
HW5WLCvfdy2eXKkJp/Hoez8ER+kQSnoiXvafRs1VYxvrwQ7HYMOS2mzCYwJl5MvD7yfJCKVcHkL5
BErUGaOTXPU3ULyPV6ePRxRTDoXSBQf09idKrLEOXsz+8wg+TWcfvWZpP1Lpcd7RBIXs+V/QQ+lt
M/iUf8XZRD5V4xOK+o7VJ/GPrfGXr2JvW3SZYO/hHErgr39lWpxoyWi7Z8dRWDWRawT/dsVStGVd
sbz4jVPIWcsTpBEtSmjmVIx1t2yZXZOFxAWDwrTaa08vkjShGGa6YAJ5/rgTSaLUr++CPhbx98Zv
9KAdpnAUAZv1j3yuwSzpqT6vc/NQB+yuFWfqOUfUexkGOt0Xr4ymvWeAuGtJ7Bg5D4MEmHYHGh4r
yhwJdmMK3b0CFMB+wC8/9dgC/CO9pe/KNMeJa0dMo91aPBNbdcS3Zmqu5aAmoC+7dO7nawfg6hI3
wJ9OFBN3ci+itwLpS/D2R+IGe4LcM+GVUEfbQFdoCtX8+KsBWle7DJzoPAEvz7D64bk1nxL59fZM
hmduP+Ecag3HSJpO8uVra1LKRvayIE/c8Ujm9xJXLfn+rCTgZSq3GTHVVabVsN/4XInVnptznaF1
GxaKjX8AqXlNp4G2yOtKdIQmFQGv09oJD9XJutAHlraxaBJ9sRa2iSGX+tVa452FwtZtaI+XEmhz
JVSUgf7ENPYn1JLXPyuW64Sl0d8rh+YZVWYSrp0WX/wrL1XP33HVIQwePc+rv3Uhs36X4os/CEvp
vTzDm1vv3G+2EFWAn1o+IyPsJ9jybyYwz3C5+vWkEiPS/QSOTprm/7DAYVND2qm+aTa4gL/T66p7
ws8UGu9kn+EgNyz3EwEoL4M7Bs7kFn/VvqyMVprVzpg7tIMqWB2okwJBZJ20vQ+S+G0+rqLYgLod
vDu6aaQ9a6LVsvJOo+SAqg5JEI8Yoq3XkvS90ltd7/wGmYfsF7hUyz3YidBQMCFslOFEN3uA0eDr
UScuUAucFJZulbURA/0Owt32WMdvyh+rNG76GTFfkGYDZN2Ss6gEeCYyJQziBj2DuE1ipHZeZWxo
Ow1hWwZgMiNFdWeUm/1SUKJ2+GRMtbpsfrqj5l6dlhiqncHEAzzUX05a9e4Fh78IJbFCQNVYVSRa
AZ0k8j11+IFgoAvWddowH6E2oElU0dmgGEpUqkj6c6vWHoQOCh2b45EJ/IR+urdsrvmmrFvzvDWO
WH3lSucwPneRzYpi+XHcrVPkrGV1WQX0omZFPZ2YseLfWQ4whR3YU+GRmTVWqpcGTnYiJJuJHGB3
mJ1PP77jqpUtpUg5Uu47qUJtJdBKyBV66RTWwlAa+tYj6mx3d6X3Ka5LClzu2iPpCaEa/n8li9hS
U0AvhrtquRjDFtQ7zVujGKyjVoVo9Ls3VeuKNwlWeaYhLhG7cWM16BFnWUTxOw6bOaQQa6/VMlra
upgQO/RKxPf0pTFSQYiamCFOfIDNyVFl8XsJ551+qtSmy6W1fKuZv0iJDqYpt8gFeVCkFolKQV9W
zXukC9dBNQwUsmV7hDvBXPYykrwIe2kbIRZwK5T5CTCVMdJnrXgwsiKkn6oK1KoU9e+FBCx2tQg6
X+kfxSab/T1TWP9+QH7Gj4METpJsUG4wyIHlJ6UtwKJ5yB1t0bS9rs6/edcD6xLMc37uuGl6kSYg
XyjeV2CmWNC3QLGa/gti8rTBFQ08PY/EcopP4sSjVar6GfrrbZenpE9LDgxiFHwTBzq5HSZuRsoE
IYsP4hifKQcQaHaDyxf0hQW8747Zd6RIMjXOGNbCQfqWTBrZNfWfX33jqWToRKN8bAxTO/FDY3xm
UcVnchFqkbBsLAqfCnI6byDqzKLWxtFjdH78X1X8u+heu3WCUYm4Zlq6VrEtyUOXLOazZSv9/Fiw
07fG0E33GW8PaONcY/ayhLkmLMGTQJN1ovNZn0W+WYqMG0xm/JFjCoCFvodFCrSxgDl0AiBvo5eg
Bi4TokQhngPeXqChDko6KdVmkbw6MW5Yn8G+tASAKwXUkYV94IvAmcF4vSw+ZaovfZKtbbIn4I6j
RaLQtWkgul118Wrt3Ky6N7J08xUdpsMd4zpMrXVRButX4OkpNs9leEFhGxBB2wcMa+iZwTzqJzc4
VohwZOnGfzfzwrTJzQMHPNEpdSgAn2SMyQSz+1pUAph/zpgXfeJwzouDOz7EgC+Roi2oJUP6aHrD
JCXRQeLhM0fAEGuOyuaSIT63DjllRmDIYrMgtdGPLO2cMss4YSoJYxXkucKYPv9cnrZbBaBwKhTX
96/0r9AOVOOwvXSOv7m1QzuW6+OZYSsfvXEyXyFnav2obPXkkNBSNW/sOFbMT8+n/+7UgiNtiMkM
LZvE2U4TyE339NlkJgck2M3NpLE0CxMdq69d5uyahib4zE+AkPfd8fEZ0fVCwhwIhoTElMOfjKPW
Pha40BMinGnni3HPCxin1QG31hipA66vHtzKL+jRAuV8dDuSe9q3ir/kkKLrdF2tUHuBqZt9DD7W
4rG/GJvja+7p8g1oSne7gWhgYpnxnWNJCHIV0KM7yiAvY0PqUZv5+rap2kFNgEOncOssq3Ioj+4b
VgdXjc1uzjqvD/wfYDV7KeCAVqVk+rF4+LStoVaUdw+9p5gEu5kjWLIzXeQJxmwGlE/w/CZgCawn
s9VVVhWws4CQzKKFIcl2dnr7R04Wn0lYyX1JxlntYWe+KZnmuYNo2UcCgehUuPlHA3/DIzj19hfY
wmpyLnvU/CZCZzJZu7ddWcrT37UXQqoM0xs6/pmP2dBbmW5/pvO/HKodxf/yK0N7mGASvqlqJGVN
Oo1xWVxeb5hvv3BjP9Lg0DHOc/GvD5MS4TQdtvrnDyWpJgHlNad47eqDOu3P5eLFYdiJ5/G60RtD
/ZPk/CFs3L8FO+rROCJVRYVJ48F75wUOmmgokxEPunp9m5aRXleEanlfYqs9w6KNf5VuVu34JOiD
yKjzep6I2A3/lUGJYRPdnuewb1slFKWDq6cmpFUbwRlCWilOQa7frEBUznzJH6yecoKvcwfz06oc
381U6ktJK8hPoBnYo3GByE929pEzvt5iN6opHRW3fsIzydmk6Migt+vidQ6jSKrYDiOyA5v/YiE5
UmDXDhrm179srXOvKOhsMN0I9kSVtFM9o/h20htT5NrjFfUBkdNl8Tv6p/QSQqFAZMkgrureCocJ
XuuRAKBjveuSvAvMFQ6dywY2tUox9W7bp1WTdXo3Lact33maZwA94pZKKXf4g/jN/6bWLn/Sy/qp
W2/N5U5NXtmo0Cxch8iDrmJwLh6cEX4g9MvRcMNjMAoQag4CHcj29UGASo5RGZu0GILpOZNBK6PY
Rb/uq9i6IQgZRR+zdU5FYaFB99N6q9rU2lUNJQg1wSl5I5IIfSLLHqNXvnDGz5+jNrNrwgbztwJT
Y0VeCU+LLuSZY+e3IgXtT7JaJLhe9RmMjWr5wXq1zUIqHKxUlWh6bWuWISHW5t3QiZY0duaKfAtn
yuzRPnIiRQhYnYAxJ2XS+4jJDOpPvBBHKUxBisbAg5t8Qefi5P5Kx63tuo1g7RP+V/UJwNIyIz7S
alUE6yrtPzJy63Re7Ii4O3GVGRGE/Awea1nMwgaS8BcSpVAUg426ze6tvgalz97Gg2ZHLHGUnk0I
pRYdrGKo6B0i8RoK9heybXxg8oP0LSf4XWxq5pKHhkCO3V5AMHIDxAlbWnoCg3ccBBp/dwYhjiUx
St9Wl5cjrDb/zKzN2quaRuBB78MZ0z+/s7m5I0W6sTRB6ilGP992wJJbE5p1BqVgAUOqoE56JxOb
aVDjTwBrMH6Qfairk4qpgCl8tFUsXhn1olVBUdtCf0rxtCReotRJ4vFSochfIPCEwdg3HIMvHH1D
ZYWnEid51U0YToqgX/qBgp8Pwhf6JdXWXai4bmhUzKHUtAnGs1+I8Wv40svfqLXZb9Qv+u06Iu8Q
g4pEc596vkhQO/VP/eCXJHGczcZMpZaUs8WqM61huhMBhz2nV8DDR52nUgUq05XxflVeDb/KamXC
Kjn1DeqHo1rqh2PteMeOkZQiA0CxaQB/blsjyRmM1gdohUlODEo/weA5esw2h7ue0R6jqe6PYDID
x+zkFHj1JrJMDtDuyJ22ZgtJn4Ek35SozgHlYCUsdVpMj5hPyap7q0TeMqyLyHhe0yuHJ9AItvTw
wJdKBgJTA41UQHRCStXtJ+GR14H+rK62SjwmgyZQWNNkKs8UnhUdxXlGI3z0NUsUZ5JDdkErFVFm
Tz35P6OUiWlLDFtcRsvW7dklRS62Q8oBdZME6jrSyca+tW8b5YGs1kF074qoBDAJis9PxCGMCdCf
Nut5jf6ByrQSU4M+hcKXQjBvcerQ3yoaRthdW/Zmq2PDzNWxPcCLQfwPYtZ6ssQzkY4NlVA+SHV3
ykbYOWmDsmoxces0oJA/JI4aBt4MwLTFQnZFnms5NM/RNWbaSh1r+tiwQ789mp4wpKxZ+NlMS2Fw
sexg18fvxWBXZT5BmFFsjuw6UfQNlNxs17RfTTPDQuxz3hbR70ca31pACy5U7rcaPkQN8wecKDrF
KpkQJgMwoJbxWwkNbWcHsGP5evvbmIs+j1uZDRETu8V38REcQBdbxipqaBcZN0xW/5SOOErPBynP
NIt1mhajqj5sREsywd1Bz24obnMfEK9nQm8II//w0/3NScc/d150pfLnjaQOb4njrdjQ969pMDFZ
0ydqx1oUoXyMZNXWD7rUduy0bAigj4YLqp3XfDc7nGTBn/g1mZ2HfF6J1kLCxHqnDowYOmTpNvuq
mRQG0k2B4hJ8DqJtYhyt51CcWzz4lndW+vq6gTFCfKD/x4RVZdasVZRpm9vGmKAlJRMCCfuxbRA7
SUtvP+bboRDVEJW9s9//Yrop+dOTvl3e3FKde5oaOc/YokkmNpG1LEfSQ+m92Zp1dxDCcyYsyeyj
0+kmsEjsy6G2XT608qxA34FCmN221IJRCAMhZ7pc+IHJ6NLIfEVfQ0xsy4X4f+gmgEFGcubavjrc
AWPkaZzZ0HwVOaA2nNyXR3oji3IQuvFZ2HkAfjExaxNG5/QCU2i0QZaJdS8jcllPIgl6/6JCqLj2
nqWP+UdQeZhCXDjs+rXNJ+aM1Vit3A9pHgTSVnhlIa5Uoe4B5nB3RWtK4htku+hqBNq3HDjF8Unq
LUNdYTGpDdQbcMMUnnLZXXgB4qQXbSKzWQJ0cszlcYVtHRLZMCGnpgcFAdMmx63udKuvTfA35aYl
aKvSqXNjCF/pXJaEwUM4b6P4mwoiOmCCTUntr/l+lq+HxBLQzjOc+kR4oSsCFNTBDQHZ2887c8kV
OOQmlJIaHlacZVs/5uyAwamKAckI8bKiFVWLLAUtWYaRsFglpB8jO/7suvjhxqWAuToSoHWAqS5o
5YXOMctIF4X36lGVi2r7jPKUZqmpSUXFDyRggqJG6nuA45GSUcKZ2ydNx8rKxJlL+xGqxsA6vy4d
38u18cb+NcXekGuNli04jerXpuCwHvIe1nzL9Y29GzMDq0YpSxv+pSgIYv5Q2ozcKO+nmJNTYVKd
+WXdc0fIEt48oOtcnzA5nsvc/Ea6cMftca9DcQMzuh73t0PV7JxUtocQvmjTcXD1SaH7VIcJBW5c
GLqlmd24awSm4yf6jcuPTQgTe+ozM6puQFU9+bQjuKr+xDIolmLC1h0z00DNuglmt78+i0HybUgU
iPwiJuYBPLkaJYUf4lT+XDt2ord85nawE7J7xy6gbJq8MMx5RkPiW0S9N7G8UZuIdv7K5RfeQKJ/
BQs7hQcFD9omGm6IvZ3jqOo89ZCCIWG5FUdDkWut9PGVJ91oqY3Y3IDIjUdW6MwNw+hBamnHETDl
nFgtQqPyUhVhkQ7CdwnnKdrT3/89FrPqUnHsPFzo2N/m9zK0GWSp+m/1IeDPFSQ6wXnTE4vWZknr
1kbA0wxZkDgz2TpngOfyOxp7tAU4sQgbXXpyfxX9sMrLQwPL2vn4BCEoFWt/3vpqYkKvCPfkq76a
fSPeafhnCZQwrdf7N/pODwKgxyxNi1XbBr6yjr9UStRujLlmiBrgh2k8SDL6nvt5arfBmlRQwJWi
Zy5/wSk9FjWbDYcTemkjcRrmaa8hVGPKSlya5mh79hkrW0TYJp6wVmKeWxmVqjO4LhNW3GrcgDKC
pQR6qaWhLq55/MpzYcPznlMikc0JoX8Ib0yEWczZ1SORSJhCdXLQRdXgtWWep5gNQAxWybSuCQ6L
eqWpFFuT2o+F+PPzofm0NNo/hfbxLsLx15FQHIAQJfVzmHQRtYDvBlVR+2XARamrk1H/YFU8KZrC
2ABQtbH5lPHbt0kdtKHfZ8fqnVR4x8G4C0wNqdwkB/0BPo+J/lD6lZM3YiUvJ0SNCOZRZ9AR07J1
Pw3XhzbkgKH3OXm+8wYsFKxbC4tWVGRfc4qwXmvvf7iD3ZMLTeKxTQ8vsSBavZU/l43KlbUbnCPz
KuJHBELnOZkzKNM43QVCFvNPfoMGzdIXGisn6RkTUlX9SqLoGU8xKGl79SFujzZswQqDcF2ySFOh
vBEqpKyuszodQXLd7Mapx0qSaTajiGwDtiZoafsc/Ei3Darfk+Zg9bTf5MzkjvNneMEbz6ZYl0iH
Wc09k3irXTAaXDxk/E1f5rQKUGvitTXMZ3P/3gGrjfxeFB7gy29pIN0XC87tHxaHEaKgX3Lus/0v
sr4Bfa1Wthwiq/t03o4F3x7wfKo5ntUBkOK0QoYtFFZIuU3qtBHjystETeIYRfH6rZf0ygMj9Tt2
g8QiYlfRE09eDh5QkCkXY40FvdH6v9gJpfpoWRRWCLd3qat135utnclRsSymFcv/q9iqAjjiBbVn
WdsQkHxLEbvmwYxhp3eLceYnG59a+SRy7cV5858CRTAX7Lch37PLNfODZUVyRwe/DB+NtrSKVktl
1JT4wkH515eknEuor9irWz5y2LQB4OOjBdH9jQyr+xBxAXUiQb3FeHeyI9qvhe29OKMJhKWj8JlG
fnq6BfQPHnlZ7J9LlUVggTuctbkxM4LenBTneJLzIpb6IzCkcbojSQUyIyIr2ATpfezK+crtvp6/
e2KuLiO7f+z+ZIMjy8hoKWdskqJ/tFGCHcf/1XzdYn5HbICt3or04LvpcdwyMvRtkvUjTw9X5eRj
zgNLPL8Fx+DRSxAFFbx+bKdd2fFYV4tS5NAidNgHQJTuNC5ltxQVk7/DFR9TxdPKscBtzsXb1tnp
5lGBtN9VXSFsozpWRu8U2G6i3j7/gktxVxoASJRvQATI5sQmNhvAmaEVwVZ33B/A9O2Fv2206+qD
mHle3B0ipKNZ/5cyDFqOKHkg0rGWTLHGnN/Dou6LmZO9knUjyNDmDYz6bumH56uqwXW6bm8FwyRv
j1HO2kPlmdAkp4XnONh/J5flPh/dqNXz1rq/rEOS67LWON5JLm6StP/Pqa8z+32OL5O4OubTYNfn
ApZ0dNWiOzlVZkkEZLjxXYE3H4FMdfgw80UYVFFprkt+K9Mp/RkUAQfUwwqrFVz/ZQOYUG4Lu0xI
m0IUuGEXxB20X/i43gkRTLRYWNwqM00aWjqP8tGrU8pO6Jx2MtCI918oaWWgzAJaefWe9k6uvCIm
lGvKyMBfNEh3EHF6H/w5GdsmR+Je9skspbfOUFtdpxNU9NXg22SweGGk09rJCE2K6pcd+mzWKsqj
EYSD7l1qKNgNUlBSUEGLQmzPkwPIJGIElL7pznZOwGcCefVS2d1RYFCtpJpd0f4C1pD10yRXt4um
FO+pnVg69n+7u5S2BfgKAElqiuiNaiGj0zPPc1jEdjbvnOWleGCa+yxIibrSMgk3vpfpXvmWaSlS
Vj+gjorLXC44k2YC0/rmRK6TG9EbSwcoWQz9qO/VNbrzSSK/ApUmIJJHtKDOnF58D6iW2Fs2AFrt
pq0CcgXX/2T/E5UyoEGpjwCwA6oAFEucwQu3dh3oiP4jDcTaPHvYW7MyIoNDjZLILN0VcWUekaGM
UQFlIM34klKTvJhX7fE6lwXe18qt/KUdwLS/ezvbSmw0dlwYEauChTzDLbevtbcFc4w4xSxtYm3v
2DsHONCIx0uHaaz+azP7/Fp6Eugsd5Mx6siQwLdWB5ZL1tTpy06kmtigHgbP87KALs59Ve5pzaIn
Nin7ooqrH3NkbiCXnbrht+TszDl8MM8V5NqHKLQvFkpS69Pi01jxE0xwIGci4si6OhtFwq3lXK8K
M5RFsCXICYDWMgt+UR3bXB3HCMZCI1BVAHtLxchFjGhVKytTFrdAmdV/xypR2cPcsjyeHOteEcY+
neOo69zqdDN4euszqIqhonWcsPIIufr8PUKdqL5Rqrr0KipvU4+DQHovD24xO6GJm1E40PDBJFou
q/988SPXHbEiEmqQ8ebbFiz6SR78WsNRFXzE5GbECnrTfpifkenhj6h9ZHuExWdoqS4EahSaq4Zs
KCEfsa+7S3gIZWq+V7/HYWiaPj52LkPJOD2xG4ORL6JqUEtXdvPo+c/z3BjghVnCgarXTQ26WWCc
WM7PHLWt/a140ZGB09aWmB5TjqFxZ7xuI1etjXjaRDl4ZFuU7BuIRA7auSTQoONd07di/i0PfWOa
baFOvKdz9h2ws1fW8RQYL0DtYr5dYsZlmusClQQrkZBF6Sm2EPdl8xM2oT4GwVjWAdeB7jlBn64r
NnZroiyGdNhQ1Eolnqjo3yzLWgltcF4sUClLJmlN7AixEqMsnOCsXhtn0FeoLWeawHhBDVg10+bk
i55vMwvT/KyWLkl6oYLfmhoj84js/L8QH/EqdkYrYku7tcltJPnxWiFmlSVP5R/xdXmQagazH9R6
hACh2HIOdIIRt3J66W9ApexJFp6kl+yfW2kwb/NtEPo5ZaY2BlXpjStFJmGs2Tm/alCma8zuea1d
bPGbgPhxrS3iT0yktIshymZrYe5+Y0KnO4xueJ77onZov3axmPC/c/nnXS1ic9qjCpwPJ3slKzMe
wqoAxIHKjR5jpTnHRp9pGluGOFjA+ipSH+8/AOea1CybMLnQ+i27kdnHmAFj4vQhZMceWJNHSCWt
9jCfhaYBtl929VWIpyaP6eJhkenAs/BvupLac4KrOCVYXTuQ0GUlSSgg/LCV1nUc5nCvyieYwxdC
pmYEI6qX+ZV2vSEIfGrofhIHUA4YHs3nE634FlkU5CLj0m79rPxABsrf8E19QvV/A6K2twfhXVUG
AoyGFVSN4Tfbb1YLdn38kNFnVctcEaTwq+pOqedWjasyZ96Nt/3acO8Sfa0iFWwPALFoykCJkeOu
NsrC6ZgfxhrSbdglOL2I8gWGciOXUB5igGJ/wWo1s5egvYEghRSLHzRz09Mk/csJFNWlspkUcXIw
uJEEvnRlRI84MdztUpBlMQ2wlhVCkBdiyycaHMp0TZ6qPNsQJe7zp7gAL3bmi1ac/fNWgBE0Xlsy
HgvWtRK2n6R054RvFLhf+hhjRqABmBjNX7OND5jZ3EqjF6tXnPd+IlsaJuXDY2FQyMbWY4OGuyv7
ndKDNLLCHoPFgUDA/XUupKLn4mNGrkl/1LKe1XYnAaMkRjhgG0gfq+B/21J37/Pz6S0T9svsNJy8
+h7TboTMzOJJvy7ZMf+eEGQMebKMbtE0m/iucbk0w5Y2IjxPsNT3NVTA2WNdgXquQTwcuCFFOIay
c5PLfdpylDkNBKqco9HSI8hUIWiXB09AsuULDzB2WwQdixfd7c3/fwU7Y5IUxSznAHylsV4iJS08
U8+ZEbc7LKSL+gBAVlaUQ5XnPm3WqwMw/nz5H4eG/AqAiri2Pa4/C1CX8G/tCc7gz5jpZJOzBCHu
Mwy1j9qk4jJfCu1CGYyxHwFmVZkSUhjOF+bLxlHEIe0O0u22RK0YHTgkRNIkXCf/hWR/7pSub84i
j8AxXzCOfruY2fmTadg1PBmWrvZYrRnkd978Q+T92gvf6+jfXNv6sKujbewvVPpLxYjiuKGD2dZK
jWu+bLrT49lz07OvtduzZek/S82yOw5KQ85RS0vuaT9iQaku4Wb6t5LgC9oIWcfAYFS4uXjZV/nW
4L80/wD30qUZqKhimfN+5ARCztucXRgoCv3XYLRk0Etamr3JEp2DIvuBfKJZfg9d6b9/wVsvfp09
ahb8c8TgfSgMXvJmVj0eLTIVGZZOL34SU57/ncKfT2cy2PH+QWkTSUrmAxsnxEHOscJwOPZFD8xU
njmSxav8eBYFvjvBoTi7g4JtzWnQFkwU4atW9QMNxKbnVRJYF9n1PptC8m/IY8gDkd+JL0zF2QMV
5Ubvt7t/4MF1yAOZK+VQ2Eo+0uKhsfFenpmeh6iIf0HFyzwStzYaCu3PaVG2PnHi5gi6QBwkWye0
GInwjqB/bVyX3CoA438fcvqg5dEzvZ9CJrt3K7dL6fDxBOEzIydWR8KAxhWVrEx7s09g41Jte+i8
MmOwqQmPL/8QqriIaJkU8SMb6ucqGuxkO2geL7NZi/0WoOjZ6noT1/RcyP80OFyWmMagw0PDayTr
DinUCNvGT9MNeouk6xQF76qBR2EQFttWhDTMBLyRgWr7OBjkfkrbYXsg7I88FMwgULCl0GwiHVyB
lXMKVwuJLqMNlPyWFB8YMuoMa+ofNdAudKKvoBDMNFAx9EW5VJe77ri2MB0HErmIRLvR2zhf+y8l
kJgDqWarZcCCVCvOzvgwtHs15Z6ofYYEI8XkspuC9rqtjpYxHhKkOMHEdvQhkv1BePypXUtDCoP8
DcZhulD50Et2essurMl3lL1cFDbpH2Qvs9qIbYkz6LUpp/gRRs4xBN45E3V95UXLiDzzbbbpw/yC
I1lMb/fzUmYHB5JsHuTgKIE1jGyXoYTjYItJxrJRd8TKbFwBJcHLSxjz4lolp5uleBmUtEIQVAwT
uFBwMRaDmh8nWX2z2wIZqTzJvjQRnlsdau5hBdIgqJYYJfOuPeNhTWhDru6rB1JifR4hsJgRA0U5
7ZX1T18AHCEXZhq87A5Apmpy3xaK4ysFUHvIkRbGXeAcsyzcVJFS3dEhhE4jkEi132nfthGyTJVk
oP0KqkfEVdeekr+QI5P+Ee5Jpf0DKSzKCF2mr1wScdNKBkttmkWvDfLIl2GO7LyQoZ89fiIK/qV1
LQuyJdIXTyDHdg8+rehLWvWSK+QKOa+BcKbyQrFV2OrLHyW73ZAKhjHZRUAdHow/Z94FsgVsC7i4
sDlWjUPab92v0DYlWz25MOXcYS7piPtG7IOJ1j0p6AO2147gv31N1hZBEoSjEyOcpj4ZWmL8KG4p
gFKS6Ihn1BFVnyUJquZnr6aws4YJggd5ZOuCUbABzICaN2xgwBhC38Ju8D/slVwatb2F7kYct1dR
ZSyzNfcpL+8BFBq7ucQ9RQFIK/2X3V0w/8dwpkSarhI3r7ltfNvX0Z0RAAGlK4VzwB6QF0sadq8W
vsILaIDLSh7Gts1raSXoCR4jCgSf0z0QMdcRMWeH9rFuBJOFSASQ65gbGfjNicAQoqbO7dcUdXls
tuajv5kU72s6ILk+WCw8mWXkSWhH8apQpE3BNuw7ZkTakpzUZSufH+ay9uboPPfZNkn/W4UzzXAv
KfEBiftikFJc3mmzV0FW89yYM8EBRqdJgTctA9nWRmahB+Z4vTloXXrusSId8VQ+dzYhF7XvbK+V
uQemtlzd1lt0ICNsVc3Iw9oe3xPooJyHGinwHNbvZZ6PTdMxJrutAVWmt5BmHCVLub6p/yDnKc2p
w6LvXhBIRFph8TYIa+tE6u/ArZ+Y9I48oU4zbiIrYHmgx4cTpYGLEiib3rSEkafXeqNbvIMejcfv
7vppeloUpaB/6kLvS2wsZGFUOjaAIeq8d46uvhOWAtxhiQzX1JXHCiYIZC8Rom/aVmh0yObYPSG7
xtJ41o16CldJNSa3g25VhSnhaY9qP37i56WAoEQmCgbZ29EHZ5bOipjyQT50YnpSL9oQDbNgfbAw
ITLYHAdJTwbJYHIUzF6/8M0RURxz2s1UL9umLYuhSDhNhURkN0rMhZGP366HOsSZLnc5n5/ynjjy
i5ssyICj+EZVfyB2pYglJikT379DQcf1JSZrTo8qtwWu+al90fHugufCKP+rJiMlG37KpXoiRcHN
ae+mmEOGeFzP//PBcZhrbUS48jC6EGwOMqg0keDDXDa5Jq6drIuLo7UevT5n84C5v4P8jf0Hxdtz
s5cMauCX+089WmoFL7CRv/YgIHugwM95ZUxHMvglUjL3FFbp2aLAypSCG/LWI+oB81j54R80L4KQ
Y6RfSuwIyuVEZualm1MdEtCFCHLDzf2s9mK6gZ74csfO0zI/vwPnIJorFKFf0J8YoCeBPibm08eu
HSWFkFmbMbIuONsLjAtheTM+5uzh/9XX+y8r0TmgJACVCkTcLTky62IMQVA+vRO61COktjtKBBcH
q/S/8QG+B58nYyTuCAuZR9HAiKmu7lyACnsRZfmE5LTnAuNazLjAYLU7YTYmaOzMxh25QtMVAsNh
riAIrjbPZZHpxfdwRySSIDWdO7JYkPmtBWXQ575Tn10x0M4TpqqyQOWeNT5zdPQrlY5Z2/05fNOt
NESh5JDIJIqLtIhRgTjq/lIM3IersLF9SjDlsb1ykQt8SDuwjiOWalzyeDhyIHHUTaBkLh2f7xMu
hLF9hVD3XjWjsjARs7RzWrZGIVNiX1R5pYovy6DRo4UAybu0ubRzW2vbIYPFL9CYKT4FyuhG6dUE
umHPSR1IhDBXCGnTbE9MIbDcqozNyukJy8DrR+57KG7Q+lydvcLeUTHRg1MKHKcTXMF9pxpFYCpu
9cMeW7DBYqYkesqLcfQS88IZdX7Xh4+/vuv3jKR02w35AVtEiYWm2ShTNnQKIhj8zzbIR3ktm3MG
U19z7TDl0Axo7FcqmfHEHyo2U+aIrD1VaKyz4C5elrxxFxs23NH8L8QllqjVei7YgtxNLyxvi4IT
YT4VuWY1D5wbR+FF3LnyDairCedVMUnjXU/0GOFZK4QFK5VvBKhJfmvrLAijgNGVzIJOqh5FC0ek
p5uZ4SN4RQRurwtKlp2XkmRQQn8CfeEQ/ke6j6IDGnepO4x9nJuP2zT/jDBYbS2wq+YuIySkuODE
HulOxcjaojEHgV7mU5MqqMmTW3hQQBDfkqpyU7cV/laLMndYqerQhmVlBetl7K60GuiawNTZ9DLX
l1EmQ3BypLlOA9C/dtgoZKKhO6d71zq72m1qWYWCanrFq29k/xz9u9TXQINwTDFIQtkOWWzrhGrf
rdDXgB6x8ePde6JM3UXBOaeXQrERM1JaGaDtOQPSK6q6NYHw9/ZDeenyl7Urumi1Iwe2pj265u0U
Uk31TX3MMzrTGmnR0XSYC5CQIcJUSISNeE6VFk6ZAC0PxXoGL1XysyTcY6WqC6wbPycpQ7UolPL+
Mo4GnrKnFHBEhbLgwjb3iJD/LE1cfAWVfxZE56ZyoYui4I2eb0FUtSm5q5DwzEeLkgUlr/ySSfHQ
OApliDRMzPrt/nq1Qw20e7zT4GKOT7dNx2c/d/SWIjAzAVbXB5YkKfXBehza7JL0mhcfFw9k3lqZ
UUhwqJgx+BvsEso4+lDoKvVAm2V9nVstGznZRtWVbUwUU0E7hcCAAdqB9E/CiQBNLUuJrAvtqN7g
QKhc7WmpcD3iKOnjv8tOMeDFCuLfbWlgADwxE/4BpsopskYQ4GVJJD4XunRW1iIDNf574CbIGV6F
bVDz5G3MSRGHiXyqJmJPQvKeKnUQEXv+AfXqi6lHtqaZkrxGF6ZsU694EQ1i5TRYrbwDSyAMGewl
TQlI4UwIN1lrYSxVq0f36gxPZ3t0FfZUhsxwVHWyg4Q4N5haJp93MqScPq+EUY18ihm+MLCJ/j4K
bROTXwZWlfJat70GZiVWdXYNHa6wGmCiYDhd7VSCp316WGTkOe01nyAk2g6MBnXDFumJY4AZXVNb
3znRYF5OWTpAHY0W59dPU4jxxC8Z86bQA6VwNKqSMkDZnP2uyMS8nh/GaT4GjU09sZHIeSaO453k
zDPjpdt1ZinRIJ8UFLwS8wuqzuntv/ONSdZ5vB3QBmy166flCXsbvVAYoOsJpIDjfkN4mmUaDCKg
m/82YXviD+PIVOUOyOAnRKsHUupPSyvxwFu+vHFmYqdI7EJdXlzuOBRzLb2YM7Gqgcuxl54D3TPr
ZMNjiNCJRScqLz/pIVkC4dlTGhrLcCNY0d6aIuKBKvHgkcCk0ilSmoNl7EzGiKCZCSNlvSbyLOda
97/eRXFFFIB2nWFMRn6gRvhOJym+vB/ZKeqWuSUDm7fARMkPvBtvajyp2+h/zwFPCsf+AYSflrrw
Hb6k/Wf2/5bYSivoeLHYSZFQix9jopnOJwYit2wBRsutSrZU+Do5e9+t4pPPBlAoxu5+ptfwTo+E
AkizRSsSPZb4DS/ixOdQOtGahxxUMTbdehb558j0wuJ6jIq9RgY6qt4l1et5wWBnm9VEd0V7tD+n
duqP82PIzMAq2wzBuETEig3dQ/SbUawG6C7HG88ZI6U7Z9Io71MuABuzvymRKnrtDr3yY2ct567E
0DrtzftrbPKKlkwD/Pde6SK5kF1XNvFAFaeJLJ7X4AK/CG/S9D2LjB2cA5y7TlyhUSHxUuSiNX2h
JQ2afUcbrTUinfFciOLgEahd9ig2Gy/K44p1ivUWEym7LEVbSUepuy9JOvS3tqbHmeoP+XPU92fD
6H+6AB2KwOeGOtAOE1HhbkcF52zvsC1ctxYh9+/sIZwImlUrK3xSbSfqA3tfKpbkiR+XuQcpJ+w7
gk/xsaFtcSecxSMW5GFoPWaE1il8UE+HvgM0YQ2bez6IQhGHJW96L2Lg+afmxcuxnG7hY5umpN4i
nEChHQKxW/LCDaVoJ/g5YjVwxBRU4vHh7rPSFGl99u6ScZeFXq9De4L4jzz9u/rUi5t5OIjeVp6Z
NL3RiugXgTmOvfaNgoeFmyNLs/GMJ4pCew6GRH6RsPpN8GQJoyH6lnquvDcSWEqeGTYEbjFahbPY
I/epv0qdbbtB
`pragma protect end_protected
