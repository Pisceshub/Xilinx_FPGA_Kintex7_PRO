`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2432)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9J0K+Bz7PXvRqY5GmnO8AjQFYBhsG9kOjzhUnDjlhbpsP3BEuqGv1GnV
UPBC6drg63N2/+hTfema10++VNpEpIj/3OGOTarmQ8FKQMzlMZdZtHh+rDXtl2/0dpVtjv5uiqNF
9RaqqnCBjMpjnWUTaorOdTO3FUx1+nORlhSSaoYoM04ed1kk7nrt3Tx22EuKRW688HFq5gck9OSM
csTeDeFlfq4O8R5+rLIaFgn/g/L3+i83KtiqtBKABKYeKDlfaiZJSgL6twHbS7qlI66/XetVkhuf
+NU0GR5h3xpv4h6fz87KAg3phC+iqdHkq5G7UXbv5t8MQ3FgPdveW13gtdch6qrM9soNfM9E4lk0
Kqs+L4tKA+vSv9KCwNYLS0pBqgsvQRFvIoMSqKOCjFSjQX8b6OVrhg4FOLITjlIlUqrK6DiYgWC0
7FXBM8Vw0djCp/wPtB9ZNatzdgcxCrrVoSwps0ycFS5Lh+s+69H1DYm2rSXNUXRKUce5sh941ee5
FHhnLXVd6VCcyZQepMKBKcugt1qSaNiPtRJ/oAnos0njHYmomsXtNllQCPu8dqswviaBBSEzLHOe
cH9hl6p79p6yKdxtSmLcDJUjSwhGoFms/oG3lF3iBByu7TMLulPdmYSDGRQxnWGOCxQlMMMVacXX
bTCyt6tfCWg13esafMzrOHhFJpAjRHP1FTkGBXAJmefm7MGVZzsmwuw7LOCkJFNqRV+f1LnwIE9M
A6IdpVC6XsSAzKyZUIOiRThJtUG9Y71FLscfcCLZt1FHrmKhAaXXSam/iMosaJVkTGguIH5xKWUU
X1OEfhf5te5uL+2BRNWTjy01uSTATYKfVKhOzr2CC3Pcta+U2vc3/Sar3MYgNQrEs8MjARFGa8iO
y7Je4H610axfdjRfKFtIqn1AYznlXk5RfGOpiAUWy4Th7Tzdxvsy6XJcSl4IlXGmWBCE6KCHR/hE
DXLprrqD0J8QKA034dsTkoKxzOEdgNoWkkOuNBsZ3AJtGA10W32jzVSD8gJ+H4eb7ioOkq+4wa8V
7MnfrNDlnB3m2kSP4U/1MhGue3tOpszdil22MDnZNjNu2pbiiGhNuezktm5sUGD92KAkS/3XSef1
8eSdKw8Bk3pFoqRDyBaQ3O3VDyE690i3PTBVZNEPBA8xsTVl8rE3TIbo7uFNmTVMrw3Y8oEj1Zdc
ti6XEFwCnd/C1Xb+sj0Q79r8zFBhcWxnLMIN2WWrY+yBQ1H+iK2deLKsCTBBvCeS8rn+Yxt/AxGG
fexvr7uIyW1HYf9oXzFdt7GCV42L+eORimZ735UG+0XT82AizI2lcOUFA6ezZoC/5KNc4Hst8Hpf
uhjcb7OH6F9Ot/vpZa5BapEYYkFan/WoDtBTeTnUw1dV9JZ0g+ryuzW9KmKh8lHlIi/Ole1OIeN0
A7F9YRhErGrqsqb1ubfYNfl81nhc9j+UwCCiVHKdzBliSfiInGf5KUj7pMckjo6XMIwG0PhCLrB+
9JClrKBDbX1S5Rvrtggr4Cr1AYojwLYgztd3a/c8jEvagmsLYu+9bdP+6Lrzw4Fu0zWs930kPJQG
uczIphSjRhMsR73OeHPg8Diuekm1NpNL+nDCa0cR3eecRQTO8NRsRKWhcbSUOF4gm7gApDNLhAVC
Dj2V+b6MQvoTR72SFp1za/ZXp3mfKScGOa7jGJMiUtNTnfWq2JPbnRIHvqpZiQwYcGqf+ps3DQus
mcfz8ml73ZmP7X2SMU0wMAa2+jIZk7tGix/2bq8dnyOvD+RRx1peXzsJtQHiBEIttNwHfUGRRuEu
0LquMvftN5ITJuet4B04D4CdwgXHJqaFD7Ag43vlDOlLdPaWNcPN1XllGbTurtb7EFhvHoFZ8vlh
FociiaiWJfVgFAnHiePAs9fQWHvgAmpdeyjkwKe7ZUx6rDHFNlHM5W18+wK9V3upggepUZNLIUKA
9rYLmfpCATXeC+v2P+Shf6FB5zsCNPQVZ1tTs1vy7sR3Au6b82iWavfOE/hQkoCTB5xrY8ICl3NA
vAstLq9Swgo4Gxi2Tw/gqhwacgVRR2dCYVLfcwSckUzk1aY9th9u9ZVh47GUYSreZgzVXj54ZeM3
CUyjTX7Mj2Sm7os1r00FAX8G1cplKxFAeJoZex5MsG0TcWSvcDA+6ELIxvNI/5JXEW21zF1vgO4A
YEBII3cHVjXTl3i5mKI3bdEeBLHKsxEizZwODY87CAIHqzuuitz11t6qdtZmhHu23dNChszhWVLT
W2GmM5IE6AT5CkmanyQv6UfKTvGYjZYpmH/uUk45dycKZHV8XXkBYZWTkHAn/3ud+Qop14xI1jX/
dW0uYKo+nBX4W3RiLTy28j7MLnDfGVtyiRrrGP+nSZOoSKJEUVCUZjANM0RUB651H1LVwHVesxXB
ME0t2GNHNqxoBDRqQEeo8nAA6c8S4fXT1Or0467A8vy4I4mbtWUjg7RjPtvCakQBUVstCSOLBtev
GgZdPUu2ecIBM/C65k/1Spd46ddpMZpJysswRR69sidfA+NQS0XPiiXt6T73PiJjoaG4cLYEl462
kZtRh0wPrxLSoXLZtY3FY0v+Ce0PC6eu9dw31oB4yhjMPx4osMR5w401VOso7yJTynb/zA9KUvO7
PQd1c7C8mQAAklCtG8UEqfl3nhWY5mGwPXcJissJ9BdBkGIcr4+c55z2jFpKMid64Mwb9a5txrSZ
gm0bE5UgDKd9lZGcSWiYospO5ezDTXf/iT0wgusMuD6ZPhiGe0RkIoIFR304W1NvdihAxeXup7oh
k21aFjmi5TjY/hKqlqlMhD2oQG9k+bDHx7mDMjsZeIpbrLbZ0JREDoDQw3oH9PdSZKtaXESsEixv
RbItlD81sBc6kbVmVtuqm5dR0tZuu73dtGxr3jvONZ1B0VUA4/A6YQ3YMt2FP0F6ltzHN77wgGri
YDR+rB51CDcz6Z3TFwIGZTJX2SoA64GX04ub2sPpyzNj9UCFzG+xqUdQHJyyJPC85+5YDMHPaDQi
2VFj39x5BJRTYZtfL8GbgyLbndxo9aJud29Kqx1r9C0C4+MklHcYo0Xkcs4+JNM2A8VpN4/HawkZ
FKJGanHQQT1X3g7bB59/4AjQyS/r/0SlJVIR6ge3C8Pm9N/UVjLzkLjn9Sck6YcjAJtiEva/zqPZ
PA8w0Cy0ybnjF7/ZogKgcqqR0f8jceLv7lwFgOnU1yFwwZhnAcE=
`pragma protect end_protected
