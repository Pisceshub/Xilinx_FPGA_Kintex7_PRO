`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 136048)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9MVAJWDJHNzPOTKFbvhWRW0efx2SFy7nuVynm7Ssc63NALSTHMOqvZn/
AdqLH2aChUZCWY9Pjo5eNXyKP7OAmVe2wYwsFz56nnu/tO4rwE4qamf2w2L2uEP/mt1Ksz3851eq
AuIMM7taB8szD1NmehVVYJn7HbynLio0SCoFW/AtgIl344XLvRrZ2GGbUlxsKtFG6CUzOgREaclV
x8qP3C3ZLqlX0Vqw+v8LdmXlG5lSnKbkvhbAfQyEzSLFvVjJK/ErTp8Gh9WCN3O8ym7kW02AUL2P
FUnm8i6mmUh986q5X697qo6olDHWqilCyFbF9gK61zGt/qZ9+oU5wo9l1CRab+cW/GStKXPaEx1a
1YY3sqcvShmZs24FbKVpwTDjvEYOxp0DW5yYSyvxKA2L6ajUvScMtN+mN7fLcXLD/ittgSNbR/GV
u/YvXC/98mAwdbggIEEgUMZjXYB/HbFZBnipCBxgC1diLwFrv7dKSH83NdzqzPEE/rCMZqMob+xy
9NeTG12r3zabcHNUIc7Q//2vkgJ2W15Fp3s+PdyOUYeUmwJ+6ff0YjsqBuoD6GRvWPbeOkyXSpWo
GhLhMqGrr2YSKAXmSHkVPC++JzN1u9h+de5GDgNR8tbDPJey/oxRPdv7K0e9p72dpU7tI7BLq3no
RTgkMxbyeiQC1+7qwUPOxGSeCgL3bQX1OaTfSqHqWswObIZxCPRWv3o6tQhFf5Cb49XScjgsKnz7
zY2HbN2LJrNvAJ5joGjxFQ4SYDmDHHeQgSdieQ6kLtfqkCUz/FJdr1gp5J/H6CZdJIxh7SbI2Anv
K642vB9j0/bBXrTMqu5Dump2YUHcEtcXXIB3EOS4KFn776tRN3h7+CKA48uQaW2Dm0nIHeczP+dh
YP2GRG9yKVEJUcgP8vwktibz6OL58pU3b7xUf+SVJNTVZ4wcb8jWoTi5wLgWCP9VQQDl7P6Xv/IV
0yN4hdZ5k95GwHlKhM0Mlchp4bLK9jjXtEv7IoNqrXJUCgSGmijKcz+MQeXJuD29GG7vIKbHA2F+
9W4CpnunQ+8M6eG+eRvdWeQtnfdVUtXdkXJL3FjVs4uprAACzqkSsuOeCDryPZ37BQLCyG9/BQrV
xV5qxIB35+Jq3V6CudJxNEizJl6qdj5pWOmExuiWucg2q9uE1TsvUc2hKE0gfP6jZGAHnGtEi0gr
/bb0kYy2dB94HEdfHzKK9pYkUvt+z3cdzDGExihTqsMsZKcqM6MoRq3M4N7nIi+rbK8l+RpLuq5R
Qz5jZZjpBdnyCUgfOSu4cJ0A1M3+zU2wJasgIBD09J7lAhnJ5DQ7cUjXAMPdSxjuwtG2OoV4oylM
e5yX6UogCKz8aRyvHij18bqVUV5A/RRsWSv1UJ8/wacLJru3ThQzF86tXsUCtyF7nY5U57dJVq2/
q+Qvyw/B9DcSCELuFwT1L9A8JPKjtZfXeXgoQZk/SaKZ8p2FzinpNsMzpnS0WGtXgYWJUSNYT+XE
M1I2zqOYdirpqquTPCn52LVb0bgDWmWpXlJcy/A7yr/ughg5oMppdvr6esOAfxg8PFwLTn/v8X+5
WTxMidZe2ZqWLtrrsD5aZZ7kw3MvTnQZZZfeX1NGP/17m+7r/1EYTfazXTBAeJTFhQD7VgbuBHvH
6wPAGAtjZlAVjka7V7wz4CI1NkQXLFI6oFQ/+pYtBW5VlCur2gNvLa2jzQu2EboJqtSo9f+xv06b
9WSDtgc0rZaGUDkJ0mZ5A8jzKN+4Xz7ztDdr8BWTBG+Ny5ht/pnNsRCaCH257W35Deieq0F/lm/G
m2rt0EO8HvB/bwvabRWzjpR9kOhlM0Sy4yGC0yAw5PEqcNPpPs893wm98BgkjUHJsU7klBBmuvZ9
a3IKD5Ob6U1TRso4hSyBlFOULhHtF5k+/aTSq4xL+77hwjmOZgBnfQ/vM/BPNqcPFaytg59S7ZDO
LVSnmcQCDT9R9LTqUzqJyaccXMeIGlkERLxCnvaHCVv+ZyjfNppHu+8GM8k+neCAqAvmk72WEPXM
0SCF/Wxe5M+ZZ7+J1IGFpkdzJoh8q9wGwCQna4qAnmmsXW/21NmqKbEodS614WXQ8OpAr2YDblvs
LaUsLTYzno7lXzIskaAIqibVMkPfCcQMq9Fe49T3R16fImbfoXLxHdm0epQjWPx69U0G4etu7Drj
7B2scpT8zsHv9nfJdYbrqJt98UKZVUvdbGXgzuKBEwa1iVIzLHCknnuNgG9yNHNNwnyeJXDOZMvt
F+hJuYRRZ/oiBPcvSSDxM6FOAZCq/7HXdyQvZ8F361TKfghgmjIToh5MqLlOqfIEEOpDGeUBYGCZ
drd8X/LEwDm5A0nzjpEXm35SszheFQUSNW231QR1otAdVnVLcWXWlAzJD2DPNbnxtJCdrCGV9c5P
JucAYGLEbEtrssgoH9p9E6ZN3k5tIX7+wjQNuYvdhNypPUEopvi+9YWb5L4+n0x00uE/L2VjZm5A
TQoxfA2GGJi1zyAwT2RvCsG+hIGVsxFXfPeS/fBQ63URbR7ivt+Z2i1WLtEIRYgx0ey6mAlZzV3o
jbMXL4AGliMjPoMSTf8iqA1x20nn9+ci+6g4/ccrEhBREuydIt691aDfd44xnNCpQH5qjImCFeHF
DD4KPIgL1xpDkqFFpM5rUmJOcb5FTu0zkJxDvJBFG13EsMWC70DAUF2kOAZATJIpYE/c1DDIGoZK
RfA6NG2oJW+Mn/UEbG8GJwjqLqnIxnjGrJPpIuHLMm/XQts5Ey382E2iNBiOcl+YkI/qDbbV++Lj
b1fWP0qrncBU1CUvBTJMwR2MqHWHvi9gtdiD5BANe5CVEafqGlubjdPgk/OHh9QlxtkGPqNlfgEf
6lKkZlVyWAyo1hkyAw4XpfrUDsV/tMnxNAw6C13AZFzRzd1Ds1RYEXDnD027bN3DwaZNNNMT84/X
HN/ZrXrEvDZKOsMs/a3nbD1Skz/pPoZ3yexohlK410fM0dJkKEc4FFrXDMj7DleF3rEJvBygmYjc
NRxYtcrgblCCzdrmE26hA2oRaQfbiBOXG7EoOMjOlzXxA2L27Nt2anq805dnVYgbi1SSqFD9rYcw
nmM2UG3uljlnY7snXJJPnQjJJ1YYgAMy0KAmHpWO/F+Tt8DZ4Jblvt9gljjSVG32WMw54Y3ctffy
6vGclnK4TDJ5QZ7zIMmx92u30xWMq5isOi4VIgjk1D3+Yn8s4B1MkAXsPRVN8SS/HJCSTJfyurzO
DiltaWWYI7MUw2pS/a/AAOLpx0mMNbg0NocVpqh8bF/lxuvOBYRSvPV+FQ+wYZT7MJPczB6opcaR
AN1ekjsmDmaADEd9OLOvdlZbmO0HxI0tBioZ9wyaOdatp7+4c3fhkD2ser5ISOXs7zcT2LG1kpti
53LwN3wQEFfPfx1LR4cVNeX9CSO/H3yIZ40/rHAlF4jfKYx/54wbVnbCWMx8oQNp+5Oae7dzfUem
DUWivY8WY9ciVyq08rrXWQHyEo3wse5B8TE8ba/JHtLKy9+aSrjqTbDWkrmetVve4VSrCov4T0R6
in2xqH8No2kn6Ufe4aGGh21qZ2oNYasUJFVFT3sk3/uVyTe+psDl9c7FQ1Q+yxq45QMJNkh2hRxf
dvNhNHBJBqalCXqpK1hDrGIyAENFSt0n5Z+h5FibxldnNWSMDZVltUWVHun6m4LD6feKdnbm+zek
41K0wPHfEthxyLZFlJwStYG69KszryqtDTvFMkIHeJmdooZ8rv4wud1Cn4RnkPH4SLmE+4mUrU+7
1Ss3PB4gUnJO7R9gkUGEV8RD5uqgh/Po1qUdvrEp1C/ZOz/pdGii/6c8DxRqe6Kkci7JN0barUlQ
w/4WzdDLpvV91q2OODSJrb+O1lmPhcIowmEOK6a+ew4LFHuzBBsciFNRrOE+WdlwbEbZA2+ESZnc
/4Oz/WyX7vSs8pls6ucScqzBIfytCDWTxXRgMlIllJyHC/Ozb0PY0/tty2JjesLqsItBf7EBuIWW
tNR9xcYESMX/wreT+FDx+hiRRGldiOz99UCn7XMPDSx6SoQ9RmGjfMXcoRA8Wdem91ds4VD0sXUh
8ZTWyqQC5JpduseUZrUOMMXMIE+hQdoSGvIhSZprTbTsvspwGlq+oj7brzkAM03vVNxVS/AOWlR0
p8WzK2mloVWYgS7xVE9Pe4Xeyqzzye0NYcvcQCVjZyYSotSmTRqVG0sZaIAGzLBpX9Dj5vXdinLv
djy8MfvbQZXzuvu2GF/E80JlDDZrDDDinEGktVDHJzoIzO/Y7d4XVKHgE4dy79GNHki1hIHCX7w+
LBSgRlIGBBKqCAWC7raviwu7MZtGwAMB38Papd32ThCY0XaipXT0h2W5QuaYPg/mH1WH0gTeCRI8
fn/5qSAkuxK42gnzmeVe+A0pQJBHbdedqf/LEEYh5GgnWR6L2pL+bwT0VLSHGNBtRkmGOG59KJdk
ZXNIkNSYIg/p3+7IlNN9LlIo1+KUCtblePvUK8CwUyievM4IuseJjxvaR+30DTSADJkaEqMZ6JIx
bvXnhJH0S4bEr+wBcaexpj/AjNcW2PC6GfgHvyS5KK9LTfIwmF/5XxdBdNj6SriQa7x+A1sCnlxO
fSeKp24tWAOOb4eCwEWPd6IbJEoumuVhxaNt7qgwDtTxI0+zxtsoZa1dzqR4LqXm3h84E5ixAICM
QffR69D0VlU3aXkC6BqI4q9HUQ/ECCDHYmjJ2cTNdCOAJgY8suthaFCH6uOKzma4BMX95a55CniU
fC9S4apQ7jsScDLFKH5FAASa2AkDltUbjqJ0Yqgq8usVYWNR81nEl2UzZgILEK/Am/9BdQNzyrEw
DxeMA7wGGmPB5g08o4sI6h2z4QV20v5hxMFQZlqCGU6o1tVQM5WsvONFDUbq69OZcRDYvyoIhvxg
N3I58eG7htsxzCBNYHBbeX6AJdEAXeaQUzGQIaxZ6LaedU3MKmlXgLGuzX7R8l4sYKJntzJ2aQiE
hphVAES39P62RhCzkbzyaKxFr+GjvEwF8awBcWD2vnUKVFNCy16+CBjgxbaBNY0HWFmqq7S9Tl3x
d2Uh7WKXYRMl8YjU+xw/bmxuDvR+zZIc2ghGYvJzAqMyyvgRSa0/EAlOxTwcrhk2Z4+Uz581gGZH
pebZU5va2xSBvCFbDBDbUvvpADb70tStjk8boUQZUcKpW6H3VW8R8upu6C1K4IhdWVfa0iCNKUiy
SLy7eNWt3qlBlwcRqU7ZPFP7CObVkdGNdt7sadMJPKnW02y+DeJdF1l/4sW1rbk67jWAcaxTfWCo
OvAAawiFVeWCOfUM72wetBPEPABuv7NXR/Vw6iZwF9Ul+1bINtoI65onnqHVG6/RQ/JQz3GxkyZk
0Q4+LYTFvqJmIPIv3aX6H4Kt+tgfvJJAvXaag/IZY3WsFWoC6q6Lqr5YKRODWVpjK2Sgu7gRLE9Y
/USZOipsQaWNqnmsiPirihoYMSKWBYwJ4sf2Em3hO+2lreHu/OKF5G+8p/hSP88dtfl9lp0NnBm1
K1IbaGY0Fp3SSM9FCge4bAajToNiU9jDX+pS7mKKkrfzdOgP1tgh4qH4RdHTxbis9yZylz0vj4N7
zSVPFiwx+IfCs1TB6wWt8UZbMTjiksCiDgZOWoaXRo92VMm5FtLaI8Uvh+FPS4LCItin+DMr6ILt
bWli2/lXiLScHYSJGVmfMmrc67MXNqngnZYzt5zjtSpvMDpRce5O3j8PAGAo7uvYYGOcKE/7egdl
+TH53aUFsAHlpbs0TBbF9hJmuqYGiO6bRg5bQhh7CMRKJktxrrFybMs5/hBqeEAxA7m4dJMv58zr
Nxn2pCYOGMjDhhcN3L4QwZqir4PZczb6RaENWl9QMJfz1HTQovf3cL5h1RRAyLTbFCHFzJ0RzPzQ
VKLRSsPnJAkuxrP8oPLZbbRdkL28rJNu/fRhnnmRfxb3QMEhsBTFAoaizCdR3U0emu5dgK4UK+lA
CQrXvcYgt495jpJTtrTNvREmKGIHASoe7p6YwnMRP3lPKtja+13sxsbNPk9/zayOPVwiPXLnZBB/
dH+Ml5NaiGeofP0dITXjcs9zFMPYunaqFGJY2aANbMX3cS/ldZFFOYS5xeMNy69c0RqXSc8rBuVd
bbMjoFABQluFeU7D5xQjdiXWbkrBZ2fgg2uNWu4LVGAfllxuAlj5Z4PhSMa0x0AofMWeb053J9z0
e6vtJjj5DsBZ9/wrABX56fMA2nGgobYO4x9FrQKboISejtdFOHVieXFe9vuP82xjldPFnE9iUydL
s1EWd54TgKf+I0r4RdBEgg/H623DFfXw77a20esymubGhGgwXlPYopQwwrXr/TjeXED4iTjTatT7
3LGxYhfubd5xIQG1gjogt5pLfc0jcytRh2+G7HHvzw2RqHYwQyYfHdd/DvI6H4LObteHuvzpJixl
uoej0JIKA0CHEVdJXsSlj62CO898wWe1SODxqWLbxEjPEPfG3fK1J8utO6DRXUBcvyAG3DhQLUkB
hc0dw3f0sp1mMg269Uchi245jH0sBSjg/Y44+is2SFx4VsCIgFxqTQ0W7lFR1QnO3jmcv1+0n34Z
tU+bHAO1LQ8gfxUnQ5UeC7b3dUsSy23ENCsvI0b2g22MNO1+vyUWi6udTt6ziXbmNzlhfPkfP8MI
dm8BGQqksqLWQjJz/wPrlBZi8pvUNFIbrh3amEi4Z/LjZSllunPt0V8N4MFJaq1SGbAvNab4VO9t
xHhw43ec53+OEHvhpNnzWsSdJb3RuviUbFUzbKvnBuE1Z6A7K7CuMCR3RxMzXxgPZdZMR222+EF1
6dJIFGaELe5LlI/WGR3F70SMcco9dE1Aj+wisx4k/fOgdm70Ty6fIDpYoNI9u1RZuumZ/ylnH5M1
FanbcY96YmR1DoINxPFAJL0OiNfBuAaeSHGRTYr1bCCzUekLRX+udbOMB2UoZNv3/l9fYzG6pswg
cuPTkHHdcSABU63ppSPV/SAqqPgHs+p47iyFAK0Q9y4/R2D3PPQYQpcZ0Iuk5oql9QgFA38gDVia
X9edkrLAMY+eILQ6AvTZ3ArPYPR4pKS3yysayw5Y1evPNGu2kHMO2MUZ76DcxYgOKMJ1olyBUfR8
oY61xuFbLq9cztvbEhDYHLc6Bm3rkR3I9OVduTJKYc/Fv3P9DOZwiPZBq4j89/Ku2odnzQCU3XgF
dBi8XPn25gnkcicr17X8zOTMU3RTzXJH/tfvfu+lRwbId6IWf7yk7L/+CC90anSjoWL7+4fHmYLH
qvXrY1qIVuILpILc4i4p9lGKLhsgwbvuSETgA6E5cSMCVslvQuftpURlsCLA6ycYtPsrkO4mEbTq
XQm1jA+BClBbA5/W63clWQO1uA9EvxO2g+eEONAOteIWBrVyopEBzLvTb3wYhpw1oFIWwXBitqer
CIqfFgESTLfg2kI1oXUywzh61LcrOvrA+LbJseoC+6jqDwd0MNwjUE+7r360uJdkSyES+so3W7N5
Y9mjM1PPl3NP3dNcdzmGRdgRP6KoZmoF+B5iLsMLO9lD660cmmnKsLxdgLsvyFLhwYGCVdtl/rYH
kpLkvpQ3Skj+VTQy2M9XtxP9p+BmcINPnTHTQHRvoGpvtDwI0hF1D02Gs0AJlMoty6aGv9oXF50k
SUQn5zMG9w1wFkfDltrj+dFdEWv6CNYGrmlaTYjyaGBzyq7s5/tB2eORgckrsHs5/Fon9KgqaW/K
cY/qUZC8vFKaflMD9WMOthuYT9fYpCEpc0nI6zFDZumxLdO30WsqHnKKl7eEL32a1MoZA38BYwNZ
UPjeT0QJUc3OpfcwzJVLdII+6qSDeWZwtzvqz9GXWL5FGt8BWtlxsi4BQQyOIsYEOt5Dc37XIctA
G3yiOCcLGg3ZCQEwMe7/woAF769VZY51ihr5F/ACsdtcbczjiOfjrs4pIhw9LvdkkmPcnTeMAVoH
BKlxs2SJpQ8kix1hegyXOMJok2UFRX00wswSkhoCPYlQOyDcQ365v8YpRi9mFw5ImhT4LZ5u4+8e
bophOiH0OME49/adVU3v/+VStoJd7CT3uXfDpSfkWZio2YmN5eJHTfAqq+zWl1/CmoKsYe3OSngE
OQ4XBYHQGYT9n2iocG5+5sCKW3euFbMY4j3PdnUtC3jUMZLhE5wiBrWOYfrmqh7BUWRSAk3TSZAN
hOvLdFzCnFwNBJW/I4/D9H2pF2g6WN+jdjFFIysTeU4JdCmL2d9IstBIy9Lp48z9v2byi1XV7n5H
YEqytVGN0hxyvgqhCSSB32Pyf/WaakCW+eUZUtACNJZ0AXmFdnPDOAp78f4Qzl3krIvARyLAkpVY
bq+bwpC6z3TCQha2LAXx8YLrCsscE/czA/Bnyn3B8JGDcvYKAIWhRozACQr2VeuHw4IB5fRQileY
aU8fiWPHYbC0cI5ar5FqiBoCwfxr23TrIZG+ujbhn2Lb9Q4GPQv1hf7Q+lEtGnpqLkNQrFxUhS5L
P19B15iqfYJnpKGq3ia3z5axfU+aoflTN6DB4GzN4z535QetkaTMDJ/guO1227fKQcMUa3IjIwCo
ef+Nq846KH3QThOrxA3Owor5zf71cWQBADz9Ag3KzSR9LxW/FRyBxFESC2EN7BIDMK0xS7KI7ETH
PccYVH6F8FG23WELyZx5OuOSN+pj9H5Dtrhmt5CFYxT0IqZSurv5kMe6+obh8HafZgRN4K8oU7ox
rHE3CIZK3HLP++qGvf6omMY9P9r3+WiyTWBzIJjP0VF7gbUV1HGrWdqlL8kFGOudmB+bmJTEOEdX
4AW+axO10rVbUp7LWTiSPY5aJXdbHtaKZZ7d6qVri22lHcf/BiEZTPauZcllQYgCpkaErBmHEmLY
i3EJmtQdCyqnsqiDTohDomnFLQaWtvcrxVcF/ZpWn/ZKZVGgMTBgew0hNbap3+jtRPzmXEThYszZ
MQODFYsFNP7ngehk6fv88BJjpqlR2avSDYIvhEocYN6g+Jp+Pz5tR4pex1OwJCjDyca9iMa0m5BL
4BzgqKilrvrrqp08aHq3vaDRMX0DjYMgNYwwpKhLJmNQaHpfZUiK1D6rvdudEZ6z6br/1E9RznrH
a4dMX7IGL7NLpshQ+W/0p6VWxtheARzlTfb1ENdyYDVWXKZxnSVQDpfdPMXuVubLN24jCH0C9hyM
j5eOurVQ1X+yYs3ffoQonXBLNsQQRf0ZH6wncSeXrm9A05bRnu9Vq/xi1Fs5TZDrD+WqOCzxnjTP
K9keeRdswthTxGprxWW5i/TGnYjLiDBmS8qO87bRUTtSFJP8zQWRzVZfEnvTvLChTvmFHcYYVV6Z
sZRhIyauZz6btRMg+kPVZ7J/JBM1I9UwXinbX82/Rd16AlTjx4uCT2rYIgrdywarSUA/hNfm08zR
hZ0G/iu+zdTYcKNq1e85VH3DFVPzCphbEngY8hGyElgvGn91yRxulkqcNKs2ZUtFEVZd0wjYPwIu
i5ROtPQu7EVs3A+RZ+QbsXCsgBIC7otdsj5AXG/7tJHWOLcy2MU+5GS+hbuXV98lIzSsu5bpUx1s
l0vyxycCkAm+6VcXXpidoMamoR7nJbBi2EmKfgZEWdR4JLIo4YHO8FMHbeTfbXKWd1WoRYqbhMyO
4QDuLyGhP+GtL0isjW2I7SeaDc+gbhp6+lqKXvyl3x6YYTh2ra85bXD0cHNR+rQ+5UphHJeDuik2
ZsSkGw2IRaf0ppb10xzyF+B3/dW2kAIPKrXV4nToemkfZEBf2BfxMfDcOwce0LPSCXJzcp1kSiIL
8mN3AocKxgboEOgK8nMAhic64xyy9u3UaVBtaBwC/i6q2yCfodzKvHXpywYug37tvRVvUDGIPJBq
h5/HE6o3wJnROdk5BJzqch91U/0/rsJIDBMJWK6zcd4YeLPIm2fAIzWoVqrweSYq+8OIPiqBkYTN
brb+7JqlRPjq6sKUQ7LPGBy7vZjQgMb4t29p865+bVbzkjCXJnBQ6JajC4El5mLPL5FkV72MUbs/
YSNmjoqrEyh6ZSX4cj7sxDr+omZWe4lz2HTrUBNtRprLksfEeBFmwxSKia1ekaRTEXkvXlkS9VMc
9pEHbsY89jAA7KVZDNZiNg8zvlH8IqbNK6djAtNu6e0c5f40eJTQVxTo3FTXpQ/Vv5o8ZTTKubbz
wsMIasgQI1pyzp1iXs18OB2fmcDnM7ucKKyAkQ+iywO8uajp/FsFIgQF2anP5sl516ixGwmsQ6kc
DzmfokqSJRcD8HA/i/RK5bbFTNSJ5nA1isSFjwGk0kozswIeaQOjwHLRETpSCqryc54GUaLyB0lD
5XHeRiygQDWgGTu+6gLe9sNCk5OO+FgPFUvrD8fwib5ZM6VVOLuYC77EUNJP39sVMcmPMT9lgI7U
gwO58qibdCTxO7VGFAnfcX9LsSN4pKNg3ydXdVIsV+52DW8G80EDPxdGMzYDVKGaN9tyj0ecAcAP
9SpbkXGt7DFrO4eHZPP0jLif07cmlHIeczw4pjpP9RmJMIWv/u7TeIz8GymShX9d8yQ1o35osC7Y
kCP5Lm7l3jHZflUXM2KaAfdnrxF5FeXiq45VFtDGHHDNRkSgLWLQF+KDz3aWWSWRbTNr2RFv59F/
PDl+7WOFNSLiqyHfZSHUKGf3VsDk90YomRm24IFZ1hGIZ/TheWw4aDQFJb0D6zzD6ag/oThGZcPZ
Vjg8yFLJqL3VLL95vSzZ64z5Ie1buV86/f4/3kbTU+OY+YrGQAkf+q1WDgmlKR186ouUeuUbtIZF
6jHMYJrBJtSO4Um1MDnmytpk5r2YxzJLNdmaqdacfm12iSPEKgu51bXnad6fA9ZRv549Q9ZLCfgx
vPn21It1ROVYrLN6O48OJ98v3ux17qRqZAfX4bJenSU4o9p2U4GCdlqTuit3YsNEqC256TB0HUJS
gKbxRf3LxjbDccGt3N6I9g9fW9f5V8itmBOTnj+UriGaJ6Qr/0I7ibypwBvgbxlvBJMT44M1YT14
R4OU/Yy0S+IGvH+YMkg1RbiMZVt4yv4JROa+xjfSCcb93Dnm0HWQvpArm+WjWwYGV4oU1RdJrmjK
iacHHwGsmkdfBqwMf5grRYBbCeAyrkUKv6YprKXtLLi54uwJFETss1yFCF05Y2fCYx6Qxe72are4
kq/j5Wfme7ab2ZvQaSa5cDSLuAufLaKgQWaNwC4LEv0nmerseXEClPztto7gbPsZ9zvs3cyzwMxA
cDiaUw6FXm5v3p2xgsIpFdTCUtyuVAU4Y/AMlYi0y5q0DopW/n+8sbva70ChaYZmXvOKPrc5Lb/+
i5JrnoafdoYlrqrIfVjnsxL0W0ktKaLO0HnfAgP6/AqqQvARcxVPHV5sVLIYkHV73mxT6xSoloIL
BUXkwXzYq/ror8NU7drM7Rd65zeBAG5q8xacqcs7eNfu99u6cjjIaAq4hkdU4KPRK50PtpKCEZuR
wbaBwDT+Hh7tGfhj+oAa9KVycda6iVc1HflbxaxUKg2rZJ+AIgjr52hqJykqWsw7HcfgbY5RTyw9
cHuZMLjPMzm//VkgmbRJIYQEwn9mGi87RLWmxTiE55kONDFe7RtJHAOPys50fBlc/EIWBRjIGjgS
CRtXGRLDtA1vJ6HOUjukn5ZWzeu492HXjrBea0Rot3cU9edJ6//1tUgksfhyMEFwT432piDXoQXG
vp8SvytTeCS30F2hE9LRVDP82rcvuTG/qIsjQPmhZThWofUTfrHgy6MC/QeTAuCOihLtFVQp0+Ak
urureMtRqHuBJO2CUVQUeUzrYS2ZawOaiDRFr1/7S1GJyrECH7uu+mwJftcxytJOBQOb6QVGocTH
utLSuihzDCIntLVpHokAmB//Q9fq210vn/XtrS/mwtkj+u12Ro2et81Grt2P78j6+84DRip/nB9h
eo1oNV+dwx1hPRCPLsu6uJzDLkv9up/STnn8iSZIVrvSxMYTddkjDL3mlfkKJoZ6KRaUynZ5DMKK
B7URYyr/olf1JqTQZajc1y9BG+PwKo0SNrVdVZ/30FqO9/VCgu95lNJ7whrAy1u92Emem2+cv1n0
oC5IhEeKvxSQp73avnU6YmQpLztJkhxB/1usxyftp7/mbIr89WwmY+ud1dBEwDQ05X6sleCFtxGt
f2j4Co9dWinFY9uAIla4klCGfiGCodoKGnKrfFwSdhEnnD6cu3WdZ/J3Zm47JVxCQByYjhGOI1Pi
uchihGOvCOpTxAsZyWtNYkKM02+XqXMTnYHamFw0GaGIKu3xtlYCtsm8zlFc4xMe0vIUHDQY/2cE
TzYjGQYgDW5DvvvCVJ+2HAeJNKvXqy9p09fBl/Evj/ZsmcdfODgwLxEeDxB1x2BvmhSnk1kSxGcs
Gu0jLtidQFqqpZ1bL+UY+8XO54/lyDXVvuF7fqLOJSuFlDlsPNUUvbEPllN+AS3Ozgo2UbUtITro
CVps2TrsqIz3I9andUAuBSNKTPylYMPSYAFier460YtvqXTBUzqOGLLgJ3h0pCnoTuTnHUovoEvP
h0LwgOQPER9uvXjGnpvU4/xNiuxToMcvfClIY+r3u5pLOKqJt8G5lJe4ZQknh/iW8yQcLjGh5B3h
kGgBWOsvOnSPD+ZPN5GuDuKhblcbvWNb5TJYh4ClsCtsj9aSI5AoCij3SJyb5Z0AikFKm1wLshHP
VaLN/wNEiaaGTtoqyOZhs5LAGaRHx1e6KIh7BxHCmfPg03DBIjh45H2ottXB69rG4XsFhngdvnNg
7HLvWr0l0IMBCFoDmiSfTZhuNJ2cVs5S4opwv9EZ4mpl+RFE1BGs+LmDTkn0F0xv8fpMweLv6A8m
+57CmXxut46ajpukTUA3cCSj5KsOZSD39j6yyrzIdMQyDib91qPkXIXyP3SJuYtJ5T8Zzzouhar4
fKwobfvEhJ8IjPFJS0d8qiTcjEJdEgivYlhGlgqDhODm/AHJaXtzmbsSHMZlpUfAhnI8GGkO/Yzd
m0xxQcfSvMQYqX0hyZ4yrKKT0Kvyi1Y8WWPem21htxqrVXZV2cFu+uqX0zv8hTP7LQ8zffgjEZDJ
Wvfs5pMRXXIl3Ax7nf48MDcC19vOUk4waHDbs4zq4pAp4L2xviyghdL6RK8pEYTRk02C+iYwHOjx
3hmdNOI1B63Id+5eP5a7NSOOlvpjzyzOm7IeaPxjs2+/Gqfiz/vAgBq6P8yU+iR/d5S/aFJxG7VP
RBpSWnyZWIUCI5EOqFeLadEZohjRS/HN3WBogqSyISYfcp36yL8ikoW1dqDzAaGuKfmCWTaDdihf
9B7Aqc2m8D71Xdhjvd94QPfoK3bBA1iZPbIcAj7YdqvR8K+w5FCv0IuAvoWnJihpowyF4n+aFksO
pLifuFgkRHTr64NEsb/IvT35JmsIS8KKCVDDKKeR6nAmx2gdDcxPl6z+nzzlk+icVYM+nHshZdvP
gVcsN06UhFjZQesuoh3PBf8u23dMrxvle/6W3K9HiqugR/rZFKWwPRjoT49WKXnoHlU46pViHRiG
KbjHieO8UBzAJ7KT8QqckxE1ZuN87uJos9x7gT9BV8Gv01uWku82rPxRppNS9OYHBUjwgBF2V+F+
4GLd4FoP8vRV4DOl+okk7jRi8+AO2h17P55szJq0aUcIrwNXAmPJbA6LQf6v3xn5nn5OFhreln5I
ic4Dngh7BGg4P89nZGVq90eEI2ZGwHIugtqbYK1iGxP5ScICo/mZsNdUeA27QF54Af/fu8aCipcm
lJwduXFibzxgHp0sTDRepRL299ulySMnxsP0nu2LvQPPszza0kLfG5Qm2RixxDF56DCTFR+MkZnD
LKJJRaG/QY8y+KQk9NdYraehOuqlcIXgNL5aLK5a93tRVcItAHK9F2Hg9IL+Axrg2GoaxZ9tlJkC
1r9CXbSDGC37UyYD5GD3HRvvj+GgS29xUvIQZg70qkFjqdawU/MN9mbtQElVempcBkCC/6BkfQC2
KPcPy72jJpXy5HP2QgwLo3mG7usn0OySVVrCVyCt/MSK5c2kymT+rU99hhjMeKXV3ye0NWzE89CW
XuDYpc66oV4aYh+THfWbJvT7cNBJdFAERsL/c3KXETbzh1jWsfsVtP1maVfR0vVl3KToNxkAfD0e
LLOV7rYDMnM5bV+pS677NiJwXTiiJGXb77jgFCZl/NvV6BPMj2HqUiqqjr14GHjpHBHcfdlPIQcB
IdZR3kjxaqW17hzPqSRDMAWf/3EuxTjKij9OmP8S93dGHpY248J42D0jQ/mMzGHzXDMndArZ41+F
3mT7jEaJIm/Bx6fPh/JCxVcbhOOirFWD0wtJ5/3YLvCsu83djRcxYyWkWsSVkEkrI95IS5oXDgFP
qKwNRHHLY1hxlOuEvtxuyZEWHKWxjJ81FnhvVaCjxCUGGVxWM/6xfhY0pn4hLf9Wwg7VWUrLWIJY
QgYLR1va4jDohI1mvo9K1ek0UosquBrCipb3ySvQFqgbIn9LKKH7zYm75/WMAKKuiK21q/Nn/hGn
xDsRqB0yD0m0FENqxQDIQpGZiEul+uX0OBdmPbCLws2jss9971MZkZ+caE4AicCeSeNRJzurtdAm
L8t1begSPtCdoW6EUCrRQK/h1WEaqW0WibDuhd4uKc4Qc6MthZCH7EJQzLJUS1I+T9LZxDHe3BxO
7A24gc5ZgNGUK+iDW6U9yNZ2x5c8Si90GAf9qFP8VvsuA1Sxe5KLRdc7Yb0d0DNb/YLfgEJpxLfC
25EiWEERY824b6JaSRqA0Osti7aUh35ngZSiJQlf4qrkiq/kbdOg2cqkDqH37YlRtJpBVvzjVk5T
zHdwcReHaICPXm8ZSLmeUvpuN2SBWOEyFcnU6xXNg4yC3CdGiD8k6iBeixTAv8lRuqDo6VMYKXxF
XZtDAg/Y0mcqZgVqTZP5Bp+kzWovo8vHWwG7UgRJ7FZzVXV8BYPC9HgSpTRP4NJLIvkPxqgXG8Sx
FuWxJiTLL6ZhJC+dCyQ8mpl41wlWAFD5YmNvDxzV1RyEp4ni3qRgvfNKLXKYmGddjFeYwcsqGKD0
seD3ORPw9ktst3za4k7qm3pUjg/q95YkObCDcvL6mJsrsc5y24jL8dnMCNd6R2H5QDB8dzEEh/Ox
TKhPnMNZ5s/4kX/uOb54qDtluc0hnKY4MHS2MS2jH24ruTYBAUJaS8sazGXr08scHm/lO4zWlbO/
GXMi40vfARsuRcxzHoAGmmfkq5TulpgBPyTT54IN8VCsI/fgZQ1I2EQHoGTxZNrKRmggfSPdggSN
LGFmu+drnN4xb0plRMkS0pZmmJXZlSmVPwqlmASBfiufALdHDA9/oMTF2iScrSLvymEeFyHUsyMx
RlhwzmB4ikVSHXPTYwVztDM6pzSoEkVXgITCvgUl8+LHBAL3vofcdyn+TRXVNEDCJNfJd40/DpD2
HFU5Y4yEFXDwYMruX7pE6AlLOgenI8h7nxWut783SpTI25AY2lmpFN7trHUlIT6uPFx44/lkjkkn
2koY1i7IrgTW50faArUpjDna2P8I2+C1kk491zxpjROhzlNze5Tx3tLq51Iye4XctBwYgEQ4On3E
3rgJKHP1HUMG/0B4vUC9odoVM4Mfh2R7x2+bu8rZJT3cklRRRfh9XDNz0/Vw/sliGWM/IrPxYtlh
3xHAzqJv6AAJuqs4Yt5OdZg6FmC75pryz6G3Fcb0XbYhv0VPubI2w5FqRM70iAWr34timfg2wnFN
dNZmF9kHw4thrAGaBTcgWZIbhT4OYQVYbZ4ZXO/N5WlEsXp5I1harWEM7T0Si29cydG7V0ggQXjE
8HcHYodOOC0mDxOxeXwE3baMPZtWtzTpAM7Kph0T/+EW9mIt1T0EoQUK7Xxc5EPIunhpS/VpEUaq
ATJtVIZ2QhlCDGiG/VYxqRUWJbMUIHI52XOmnLD+SY8BMbHyQ21LELwL8wxZ6LP+k6GbOioFbxHs
Z6mk9T22kx21Mfmw500hLBKHeQ2l4uEkU/V31UuAWyuGyLlbSGaAwXAsboBN7ngZzrpgp1pUX6Nk
rr/VWiONcIXmaqbYRso+If9HgYK9NSYOes3kf3fCMDBlNlwrOXpnxmLTGdIEfxlkuc9v6SZvDgdg
t5/CxYuBRYgGSNSGDdj7ShQFDOl0oUnzI2YE0gsBGw/z+sLdcR/gqXAwHJAMmviQa9JwgSvsnBkN
Xn/CBbny/mzWSOKbxhWN7kvL02ECg7zyEorEHj7FnZoZpd61WOe4kmUdQLOHHU8ep+9sQndON0ta
szfBOX3c13oggko+5nqIJjaRO6rojrbHdkxhddlo9ImjrUdz4BeSLujpvCo9whZ5666lwwY05VoD
sAsR0gbsDnTDIE7AnMXXhJ4GWXl8FwzX+makBumYyY46iNMb0yIZxJts/sg2P+Q3fyg6sinudOcK
DMbWxNnFxJQ9aDGbdqPJh/xuKKOUQjl1j1AoZFT3xdRb6hNUlGMmab65szd/FiXf5Y4nslRBp+M9
NBOuTHqi/TM4DE13N073I+/LYQZopS6g3lvK4uycIi2Q2mWfubeTpKERgJAUikiPLM86/LkZPg8u
b0GynzjojeAHh9ESCYtq31TUWmOcaWY0OzwBcaPbwpHURVbizOxn/npkvbZNVGz9Xn0L703DES+3
TSScJE7gO/hJ/+Q1umNSLBO8yU7jMfyIN+Cs4QqJh4xk3MdL+wzwjwzGek9BLqCdUcE2Ms99bkh6
Wa2ILSEZLW2C/rwSDx4fU0GEa+z+QtkgUzPCQSkP7XAa7ornnmUA2hvFmvkVLlMdAPcx/FHXE38O
WuzMfnpNWw9z/UR9UhAz1YNB5oSxkDjgHu60qlOTwijimUTrjeVouherc1aBitQ6featF1GprS8C
Kb356ZKHUhz5Ji3IXEpvRMOnox45c0ZiEIRQCPojlXfO0nC41vzAvCeKtoNN0zt92m/D5m5WFYAq
3AegyovI2i2/OFL+dc1ktnWc/blvxXt3Z1VobKKKMurA/mky6lEmytjuFDaS2rSXshNI9sUVpwFI
MCS1Zj5SjthP5dO2EG/qhDylUqMAAlQ1rpxWvQJO6ZABUv2WYAtoHAwv/X1J4GzZRDmynm/vIYvw
T2mqZbktKd5P4rrZ7qE8weuzU+WnybUdyglET2EtoeY7V+4K6W48g3i53ld5cn9553Q+Q4S5A0n+
2PY1219mFhSmSeRJnpS/pZVSX8a/+skwOBCkoZ7CxFigxix5pIr76EoK8ovaI4llqH+4mXKlUKNQ
qaHZWy6I7nX0yxt8MS5oGxp03xEmDH2ex5KU58cipLNj0DUap/FmXEa4cj5BpErpuen9NkmbrZmH
7jF11R7IrmrKfuul5P4ZM5+p06EZ9rGSVdVhAEBWc0B/Zpxxni5xa5PtXHR/0Ypm8bCpaBKqBu+o
8lA0/eDrYtyzhYFjmCaSu2sOqhLYfgVxoiminonEiza8luHUE/+MV4nbdjzYqLq5dQ4PIUuHcDMh
+Ga4mnSrZN759Hb1y9gEhdjmkZfZvZebHcLcRJ5xg1mzVHMMqs2WeDbtoFhZWPYqn8rlgLJ2yGKH
uGtE80kXcqOousQlBQWevZl6GP4n00NvN2u8fu05NEZJetb5x76Ewlazx5e+hI8pDb7zZqZIN5Hy
VTowYBBiaaQR87L8eXVALlVhNdVa0/qTYDthyl7XxA3c8sltvdxtoDbxX2ebWTdl1Ag9Vx8uT+aZ
IW3gR1hlqsELRupwGEQSnGf0FQfxw2sv3n5rAwigcP0Cpyh9qaKGAE6ve25jcBfpowmV0RHKOmQQ
5f7iban2Dgwu+9l1UET+z3LfpCuym33Ge5AEebRNzY3Abl7FbPaBCfX9RW9dhW6Yj/IxnnXcTlCO
iDCgyxd6Nu9Hvq32ghgVWXDWO+45Vjtt7UjSg4lvCSwa7E0YWVKWo5D15Hd1PYIWyTSyWvsg+p5+
WyJwnh+00Aid6g3AFCE+CN4xL+JrrofL9kttP7TiE3CYTuQieTjjOWA5XWQv1dTTGAC75BVBy7cc
3R1hfVG0WEhzuQL1C7SdCp5MayljJO2iUWjxJ5XWWg2j9DnjPhiS5110G9ZpO+hqn1E55slV2hVl
UcMtG5JOWWj9/InPt9PYVPtVfClu55YW1dq3bmEGpuOszPd5hTUuTOoVi2fqqS/H0nS5eO17F/Qy
gG7qb7nLWTS7SZ/3PLlMP/HsbwBiYX7+7/Y3ttxie+djDh/307VoOr7k1aRyW2oTCM6hry72GVeW
N0hZ6q+4g3CTDlIJeYmw0DnoWvIOi9OKltU3ArblfjjSUezp5JgP45B8WehWCpWkAToInnL+Xy5i
Ya4kZFrPrcPdsbj/KkH5e/np8X9s2mvMVtIbXq8YfMaQiY9mPTLT/GUo6NZTgVMEsyC6o+LggU3P
0Ix3tWG89o080VJyb4D4f8VvvtCwHMcbZuqt+UuMR10NiaLZPuyNOqCpKxERrfmVOYJeCV6fNEgZ
3NRSDrcwRw+yKNSVSLPPV4Qk/iHp7UXnCEW2Rg+N+usOTDiTZHzGfVhr+y4pBUY/EzpTX/ljqKzS
zdBHOH0PCVj9Gmww3Xb+qb8gpEwcmWJEA0v0nhggbB9Bn2vbeTnPVrRA2WMOKBTeIjApieyjMrM4
cwdCMZ8r1+93sSvl8cQ20ssMxvhM0Pq7ZJkCEZ5u4Sj3Y7RZ0cHHefLmsqznkXjI+bpCcKUViiWM
I2TlE3W4ryVFZeQN+ZGI4ROtzi7DjBW/cejwnk1LlHKL2p4XfC+iqF1EVO1Yo+dYo36X6Vz0OF5W
lyYNnhw5E9eyNRoNA5QeEqHs34jv8u+2aFhcSHcOp+muT+yQP+wgQXlMD46SFi9+jKCLcWL3yp8o
K+fhb1dM4RDX3qP6+4cW9tw6L3adB5pSXCzdStjvSSQmSiLceHsbd/f0i7/UiDCpRgyCldqx0qJQ
c9O2XNIkqrrQy9RjHgJrNRRmyekS0sBv5MK9Sq1WFiCcXEiz6Wkf0oI3awrlvjjLg1u8ikzNrpvK
CwWR0avpH/fgIexzSAJT17HDnVKzP/B3Sz95j4eaRft3Sx+7A23mplh88HvPXB4XYHboRJGsCevk
6FqEC4rv6ZTbksOi1XwXX3bpDKXARB8Ir6VkQ0HJa1qSevsHXLOcIlTxVUogoZ67gqDoBlh5iZYk
gH0iaUBDAl5SLlLP6QdPy2GbC3OPKgB9B3/hceZVcOoor5adWiQlFZ1L3xSsT4CN/+dJAT0YY1g9
7MJ+/4jSqlELSxL6Ktwk4zZjEBCtZ7DXbtGc8oEe6QKj6ZlGWiGSLOcLWxTqcin7/4p05pc22JEO
uyChpCx0eb9+wTjHulFJqKBeLhPRCXCFW6OWK3TFEhQcBI8PP6vjaG7X+qecglWkHHql4eQNtFrN
VNiEBWPSola7eTAC24u/ntXBqDu11qzbBKtcwzs3kG/7Xeie6OHInSkQa0Bz+gx4yjOcedUp1LDz
Qgq743V7lxR5KhfEdLv2V76cQyMdyY8gJ4xzVuGPvF70lRHf39mabCcICIGUJk7U36gnHPz2zki2
60kX8rSryIIFaLSWep/Wjt3xf9Bky2TTK0OUi5HhOuFm+zhfyIaQzhgOgLpVyO7vbsEAj+fWkEw2
J/ReklGDAblqqunzWVyZ508meMCmkxIBwVMY3IahOMYbEmKwOIaLjQxIKu+DG5SIPRERnJI0OB99
qX4mG6ArAsRr9r1cRv3koFVczQ6BbPAhEPEYP2efd6sXuK7NyAVoaWV+OdS/OGi2utzk8tF/YrZq
xOxi+3RkPxOzr/y1CX9c/05Hll1EPsCGRT/fuxRM36TkbrrdeC6gJL2AlxzPCUgYayRLS4WEfSrI
LMaVUqwplRw2BCstUDPWD3qjkrQZLPvVGm7C5WTqtEzdUI6KJqX5c3qjoiYbtjS7z5IMtA6/h0MA
OuJ0ml7LFLN31XIWBLwITfgJJvSIfBJQdjg38GpaRr3fODckuAIsbC0dFCgSW5Warb7a7GwTTJ3X
HlghWNU8DSZVK/qG0HbhDFfg+I6opaVwxQ7OZqe+NvgIf0pVmZDgJtRB6X7wyx25N1qXrvXN7tQB
l62z/7IIRb0k7liETo/PGngXy6leTSKDPoiAxuM0gwH55k66tMDNC9FelJCinI22Ri4HorllL0N/
9p0Nwk2RRkpFM4UVIp/LWBZmO8AkgxcZO5uehiTXnLUsEa63topGsWfn25quTzAnBV2bwcLQWFnt
dZhj9Xd/t8Zf/1kU+TqJSgeNydyp2W3UXg6goDuGO3ASM+DAOFkbIaqHwJs1UzZ+u8U94vNkCVZg
wda4qsN9vHodfUsEZeZjt4yFNZSqeaERTWWGbikWWTQ2GZulxARVt++hdyjkXKDK/RqrKkdQTDDG
ehYMH9jyiylCkYWi6UayT0NzXd9ajlPX6ZFvmqj2yi90cDNCFV/sbnIPYlccsxVMNBMhsgE0UQ+F
UZ4/lVfnXIEktd8qIC4k5KTNOas0CHoUVe0egDKmwacFzQtmobxjpYC/fcKNJFmrgK4b02mf8ADz
rKncD3mmxbuJqJDPOP3n/IHL1005tG3CxeLwRDMbxKMG/0SEH3u1lsnnEjq5jD30XCJJNiqy4G+z
dTFEIMjSOhKN6cz06D7Zat6fwQ+uehNfoztINno9RS5g9VxFqMIpUC2PMqTrvFkkqymbp+PLKkv4
auLd9M5C4GAOOfsSocqINyH4ee7jw60BFVb+klQ36yCK1HaNTDP9GX2GBNxT8DkKrKMn0wcD7SoU
2bwH5yacSzvq6vocaOLmcIZ7/fxztZbTIjslvoUwGcjyoaRicaohyMlemc2qkI8kFv2KeOubhrRY
q06lHVRZbMOqX3rPQr8NoJ1RjV/ggrXInMZGcaM4xkr0/UNo71zox/k3n1ow3xzraW0vJrIT5bRX
Y1oEFhKARcEZFD2/pekSxRU/wDBHwSqrBefTohH3/NRiFI0iYrEQqAsct2GQqAZ4qtQSCrUwTQLg
Fz7IepqsUXDcM7tVpwQK3NEgOQGDYqgbE5qwjS7SFVV/h3xtahvRac8qliLtwu9fz+FpoljX81dL
dJS2vvC571E4m0+OsuwVIWqBQC0ilAtslMD1Efad1ZYCYCySg2Kcw4OUUeHJsPEkYIW57fiVciBr
gWni6XfDO31P8zQtQVvBdd68xuoIXDllEFPBckYryElIiz3FZyhEyaGc+BSFVuGH4p8Pny/wHcSx
QVKG03a7cGEUsxfcT80yNJW+RKvt1SiNFcTDDCebTxzQW2RPf/2cGASkaiCsfyY23I98bvCYg0RM
aVyB+3+xbzEGhS23oLbAGNvWYANI8aQGr5BnY7ho1+QB7CT8mfkmk53mJYz8mEJVxZABwq4KTac/
iaUurXvtkCW45KnEPFSJfd1xu6eW5fm+tsD8ssTI6pAD9QIVooqd5QQ2YiqvQeFIdctJLd9/+HIO
tu5rCs86yZ8oA2Svij294dIHbapowUjaTdZH7+uaFHKc2JKVFW7G8efeS12PuHLgFE4+FreFMEdR
VabKujqD1QK4OCrPXu+fM5crCx8pU82OJYB7mUJ2EUNcAo7cVM7AaIexJwtqIwnzFpaVBsevATV/
GaBzRX4U8y9EU8siRmdvDg7nsmkCFaqJ1sQfCa//NNBWhdlDGaP0QZghp+4TO7OCMZxO5aRoPvac
HuTloJo6mlZ+8AyYOPzIs1pTFS9LsSYKg0rK3RFakw4YH5Aug41NIPrh8n+/eaE6jkSmjKURYhtV
C1VV+5rRnBmw9LyR+iyZxoaM01aJ2iGNyZuCoHc39xUnYSIU2MigUCcp905lCTiy+M7LmOOWTGBm
5x2N9BHMSRTb2M/sgNbJVVhBtDlA6fG9UYouSS4k/GI4yDdgmAmaEu4UFQcd7WQfhaNNARFwA50R
T08dMAruy+b/kuFmxdTysVCMWnssCvzNLZA99CaLafq7TJ6jgElUBveVM9m+8y2U043f3HUED290
6IOxIvKQ/OjoNdqoxCbMwZnm1hcxPfJUszDaup1hQgTUO/740wxO/Ra19WlxVS6CjAEybbXfXrpM
H2j5/bOEfpwqetmq6jifKNnrG4cObTGAGtOYpZRZ/3EZMXpe1OyUh9y+Qv73tU3FfJC9ntrQiwKq
kDK5427IZbqWzaOoaQTtLjpY2gxO891PIsqGCPW+GlamPGMMwVzbTvUXOBsdc7iUZoX+U2rl84/Z
7FI7zmL/Ju34zVU5tjDQfVaNrzxfUefB+VCkr2Mgk2Ck2nhMw9F40EMkj2KHtljLuOzVDx8Rg6w+
/1CVpKwtL+hyj5QfEGIwkbm0mTdF/YmJ8LTHjG1AWHw+YbamiHohitYosAsFgcOufQdw6K1qkOJn
TOwAgK9Qfbp2oK0AlvKvt7IcZ1hnf9+ubjFDCLEjZhdMsVsU7eKaID3oBxnOHUcjXBFiUrXs+nRV
2P+hqZhbWWSuZg5J2Nxaocn6P2VnWameQpRy2qsxGO6FcRoU1hh7+80gFkeZsJhczGCVeM9qVZRD
eVjaSdJ28JSLaWUOuri7GTFFP7Ue10oikGVnfMaF9p2PnPBcXfmiXUN6+7IbemsFBqyu3qcxJQso
EQ96urf6icWBs6gockheXYN6cQtO5SDJddHkd4Fjz3TkCyWbKjyV5l49pWVNsVtDgRPCopEZJpmp
Qxl9/Y4MS/K/ubkCncIx/3y+8Xj/XCbY8GME+HSFXqDB/BY0yfGxDTGGXugxukQU6AIsoSI3F/LT
aBsBW5J8c6UyHPpKN6QcGPMTQ855SRtrx+NMgXWS/FIm4J94dpjAw6SfIRVrmSvwvAIB4Ik0UmKB
fbHXI3aAIbH7qW0Jw7+67ob0qdvQHSd6GXVlQIAd19XtAx3RzOyTRtBk/NsP6RDO/Dk/0LYTenh1
4Ev3IRvduLg6jG2wUTqdvM+Y6pETZw+z4C+WGvAxDxOmR/aNHu6kLymyeTHtn9jbO/4751aroaHT
DOVgtIsEgazImUN0b/ZExPfK3RVpamzRGS4SjmnfdRlRgQv7oWbZJIN6i8yP2xRbeO9RYBCfOg3f
Ao9yxxQpf4VdXzSb+SjvAKR9rD5gXHMBrziHqzKoQ9UBc0YbUgqY9ofo/+xsFShw/1fDdkmXNW56
XyG4H6akW06VgpXDiBi80ijolupUxzVzGuOWpFjztyhcviBqXNaCVfK2lNrIt1UHVlEQQtoSPdSN
MI3PSdvvTVylmp94ZJDVVT52LAwdh+Fu1o1O8rmuuQF7aoN66aBdKqg4oDhEsTG7nxi+57KSYg7q
oBxavR35QxlGH2Bh+yoO7c/UbsEw1Bbk6K/NtFcfl8QyaHCWtVa10aypej+qjW2fRFCcgB70HyWf
knrL5G1RUq/RVRgWJwC6kUpx1yN6f0nFgmb3g+gZO+wtFM6MiLyAiXPIgbJjL7XCTJBszrmpnpCS
Y3+9JKCk/xMfEZ2DMgsYFTxiyIfCnRCSDVTB45dNLXRgwo7Jgst/J+1kySMPLSejyeWmTx2YOVI5
Bi+6JlCSNZiIUfpql1/NBcsVu1UmnrpyLuJWmXZrVeBDUt0xIf7Bo7eVTCMfQHXRlY7E4Ib+V5Vf
3BtlAZCc3M6X5oEowLY9QoZJwH7jnXxSjeQAt9LTAp17T60oiPAUUebW9fnqp9VRZ+QPtvYHvFRe
R9huFycCe16oRR3tde67dePY/Y45aF6PNp56YRqlkOJNgxuYUIJUskp4U4KQm8zGcEntIACTutdh
0glcjN7hHV+KcvzzNRsynVkTioU6bi2Zbw/kEa6qiyIQdo4mu2mwPKCLvX2CR8W60vIUvJIlVUaO
GpKK5/9wUKA6mhYWW2e0qclnRvoOJ2KnIVjwbYUOLl0bB52M82+a5nZHHKNLoSEFkYVzrT4zWgJW
nHPtLhVI0Z2VRxOaL8buwZFwbt2q9kEw+BcPFNXuPnjwoChzAo0J3pOvjAREdQwi+YXQfotoa1nu
jYrYKY9Ei0R6X3+4zIRvxWKaZzznYS1F2h3jgT/sKlP0B4KKbKt2mxPwEBBbamVCmoCuUVdS47NX
LRQjTh8VDV+ZrGewnRzbwjsEv5qUdm1OnLywmJ+4GfBFz9QAjTTzZrxCTNftnUQhZpFddQ7/EnvH
gLBgRvEnvxO24I77HlUgn4pxdK1x7WNIcCufdrwM7qme0rZyHb8GrKwopUAeWl3IEAyfn0HMBTwU
zH6N8/KD6Ska275SEfejpixluo46gT1U1JxR1YbTmKDVrDPxtxkUiFxu5hfZR3oTh+vY39ujthty
2AHQ6U/zYgUWV0ynhH8YdMdOSOUZZC0jl+b4aQ4OYo6O9CyQSzcCIdi9zo5V08J9jlRIYAkfQxGW
UzkjUlR9bUcM+WxsXlX5o56WS/ltZOT4MmcpJFlwz9Ax3cfUcTsP2Lt//9xH44GH7lMaEt7VhiX/
RM5aJf73QmTOdnkY2MgWgf6t2j8cQypYzhbT7uxw7fpCej7kzcuqyqI+3HSc9lMfOE/yBQ+eIe+5
hQywV1lVX5RWkRIB/tR50AIR2BfD2S3QK5sL3IK0tiM/Kdb7jr0M9LaetpmFhiqaM5v4MqV0C1Oc
rkyGq+/vThmF9C5iYpg1f196SGZMaUwZO6U9akmgtYJk1I+gAzPn0QwNeogw/JKzfxrpF4X6+88b
kXGsue1B7Z7iSx7y3YfQAHrgOfSwS/Zz+L8eD3rTprBkvI2IE8cbENOg31MVHkXt/WacVUG37brs
IY38lRDWUf3xAgnZKw5AKajDsCc/mYAKtXkXJ1vq72V9V2MtV/lDUB3NgUdM2sbbrUXA63hqoV/z
/Y1unl1T4N50G2m6aq1FojdKzuwZZABqx6edSotPi+HwSfkXb0UJEsEghepEoDZ6bgOrqXCvMdds
rQ0pf4+NeyxU9frrc0eTS+chayyDRImPn+tFXhIHmYhOLM5+o8McojMARkWHcfgbRIhkj1u5pncq
AKt4Bx75UJ/Yea8OHM5L4fhIVBkCY/upekVNi/lCsZ7ck8gADRnrRtJi++8atwRZ1doDCdb6WS7u
cIxEK4gGZgVW6bs+nLfZsn7tiD5t4Mz7CWy7zvoSsBiJ2rTkWOUOVbng3mO+JSnI91jiR+bwRIfS
3XWdwy7wjvTMcuOsQ/FWqDENv8V6ks593w6fVLU8FfjgKy0RlLeJ4I5ngrVmyIym/AVcRQu9hIR2
9Uv6tuRx4D0s20WkfplcNYiPi2U/NDiAbFvoNJBcAJ3Tru8hIdStE4dfKciwSJxuIrqJ/IZvnTUm
S7FQL1zplZeeMqF35j+lHzzhvrrGlqPfqej0LcJ2Yp/eeNyPBxwcSs5wguTBFgqU5Lg1IjuZtkUw
hCE27I4Xh3W+Y3o3dEx0jhzfXjcaMA8AOjIBiKXEe9b7lV8h8YXwLITeGubE9QlKwz6XSttSZq8T
Vbr7klBPyQSekmR3YyTWBP+gYOhwc5TVO3mfqS2RhmkMxYooGTb1eOr1B7516svScA2XpysTgBW1
EXbUlGIehqyEJGHADFt/K+Zb9s/Kdo8ckybGM041OHjMO9jEwLSewSDQSeyej8SYvj04MdYj8GBH
cg/0fjasNWgGXmfscjvZBf7vehfgHgahmwXbzuXre+FrSW/WCg5rFHjjgVt1BXhzAYFQfAigBBc8
84htOJIr4s9Qd1rPQIfTJ+Yo2GWVVbefRpNoYEObbvk8brcv3OMlBwu9h2e5HZn+akEs1vvAZAXr
xcfZ6Sb8EEcHem+5NskBOoN7GD+U9+G3i76LeT+vp2zb3agJtvYf5dBlg9z3Lhjyu2OLVc18dfHO
tnCxtksu1x6drjBWWYWb3Whz3fLE0K++qgKqlo4QaeGZxWG6PKSGpUKH0Ll9EC3UlUDz8QNyYSt3
UxoTt6vd5g7uJFolmVTgO7BymPG8HE78xiL+5ZLgsWuMquaoFeTmBdxFZ8OuFh5F/ppn8tYQc3dm
ySy9UZshG01Bi8Du500O4vi2dht92gUEk48+u8Hwj+0rSjmaIX3fvsMtO5kvrEy/LZx8qDngTsvb
7w+PkluZ5cnATFa1uQWxjg48QQLNWXi9uV7x6IgAIlsLTKufm4H/Y//aeqFgCSKg4Et4SGf59zr8
YgqXShhi0GAg7Ma9bWM12kGZ7e5G1TdLyp/V4anDu+AD8XhRAJiybFp/Fbc6/ZKxrJ/EvZR7Cmdz
QRxC+4EOWUAvtEvNk2415FD7um4n82qidcO2kMUocwU7JVhOXPCL4J2Dlk3St8yQAdGbFmIh8rOR
jSiHkDe7F7blTHSlcwGE+FKyHuTyur+xAbwxCLavyl3m72C10+BCz1R51jdu1jAt5D2ffOl1PyXb
7BsmI2vefstfnqboGaaDM9Qk4f/ZFdzvp6S4m2f951xHIdeW/dGoLf/cffccKk2RAvnZeU0NyznD
5tYx/jpQozCxD301K/Yyke+zp0O3XjyVrEn7i/XsywAvZuzwasHIUSvDKRJ51/VKfix8i0ZUaaTh
rrm8XjMJYDRkYmPQ38aFaqaK7Rk5YDDZdMckCeSrpTRtYMrW5FXD4gG69GjdJvM2qNaVdI/07RQ+
ZX6gC/FSSfxDxcktnF57sNcsa7JqlW3gv9zzXHdUIzaT5yXt1FsmuH1142v3s7jluTXz8OhqNM0h
Q2DkQVWzTa328Yy1xrH4ZDtwHfUyKn7lxkVnbARKiEtmlJu7C7PBPiuerXEsTVSq8Ud5JL9EoMC+
Q9TWa4TTB1H4wXxMjbgkmIPdMjdy6jp+h3dS96AO20IHXLjlII8rxALktHhedfCD5B6V3HsYSGY7
LI0Vp2q8sfcpD3kpdx9n9zCfT6WdG2HJE0KlWJ0u8+5hWBwxpgD7x/E7mFCRhDuQe9xc2KIlTL09
txlKK6l41cxtRg0UqnYgfaWBRHsLp25my2uaKlaHZEM9w4BTVJIzyKOrADLNGIr19GxXWdBpprr1
R7j5/gW/M74hHp0Pio40rbJ3TJA3OHkq5nr4hAZzPkoKL9o+U6BKDTDJ7ZIrZVUmre/jrnjHPfu8
lPQ86twkciftG+rTVogtWc8ng+bo3bPUUKaOuqhIHwqvT+Sm+oSFlABP3UyMJTX8xAtWOzFreUPZ
oITYsnchB1os1PJWmy/tWEJj54j4fFKnmOuC8UHECVXDYzmOqILmtbtG2s9oKV4F4Q4Ap+ZcQD8T
M/qBuxwBv+ouENivrZdxMwLjgQqQFr6HrgJIg7x8A71gtKFR03S5PEV+qTlgJfH/lbOKXJC6lsqe
V1paBae/oR/pPBu/vOeRzM7w9bst6PyFnzR4CgfRDD8KqAPaWu7tibWLbh+nCr2FCdbf189eifkI
+M2ObMAolqekEmUt1ulpeX1owfXj5+g/GF7k7hs1PWcF4rLcJXUv8eXMSiEALl368D3MoedB2wC3
dm4gBEZxw74JMRhIrxMEsrDGWC2jG4nHzFb/JCm5G5Bi38oPAaYrmP+5Cs3aSu+FakGeU12yu9ez
9/lL1CLV0y28qReTmbqilSP3I+hxc12DKr7zposctfm71y/YA/dMMlzJV2BCgcGzEyy5Nh+toz09
aHIk0P0x3V/SUxeWCoBfofMECCUWuXob2fufWvsDTxWwZoIGuKFza4mEDUhBpMeurup2IACu2SDD
FPMeSgW/rzygF1pDB9Pt7NXMlb9/p2xSqLBW15JhgaPIvRovPMuSvU4eLF8F2sjFgiuYa/92oeU9
ql4vt7+9AT7FZPxGWjKMpAs8lxgjyQfGan+opA5KbAo5JPXeySNHqvAdT1++cJzUxZLqDhhFEEQF
m0StTulZ1sVd2nJEj/T3gFZ09J+IKjsra65C57K5twAQ1h5hHZh+3yQdhjULJUXrAM8/nB94meOc
2/WluEsMcBbnGoLZfMQKIRljPRrjWHSEqE66HGT36Wzl2KHiGoppGm4NDY7ziZZ8yP7afo/zCByy
fHmJcBySFvhMKUDXAb6Am8fHG3gyocoYufanp34/pxns+sHlPRfCudQxCafozOvY1KHSwoUpM/JF
dyaebW5Sw5IvyPK4wBhONFWGefUYRCXw9iD9kuvAFF3ceq4eHQTSXaNUkQzpxU4JbdMvHwYgjTaL
VF+IFXB0BblufbkZMgFS0adr7TIFoAp4ZLqMtIdHX3WMkmEd7TcZF/nspRwbEBqJhMMP27Kt0mHq
alBWHLnWgusshq+BRZv/8+d9SixeOaJrdQScAKIQUhLprqmyoAvoPYbRhh5IXoYiduVnnYot3XPa
yJiLWkI+t9/cmV3HqqrPssH/KL7XclgUoT29/DQ/4zK8waCPZO5mbne1lHROPNz9ilDuSdAOxiLg
6J5lRq60uKt0E8eFoUNOrEvIF/S/LQk+St9WaD8wFy6GMgX9g4rE7lUBZOIJ3IPzkajjRCwlBVEr
dKsx60Q6WxF4fuaW4r3yoSZrecQYKJNvht3FrXj/N+tayki40RsTnptA10fo6W4JubSz1q14igFe
wriP8PalznW6FMkH4tiHm1tuu0ISct0u06cHYkw/VFLRvwFF5isKHjYy8+YZame7uf9bSanETzCl
lNxJrWx5fLobhw1ZDcFaNM0i6j/jL6KXQ83EWaFEfjTVnwygh5i6igL+5nPLBQCFO8nX/pRqDeIs
xvhr8T3LooFzPs//awQqwBKrMDShQIjWtVH7KLYNw6bqy3mnIl1p4GqW8U9RHU2VZk7inwTBaHMP
Lbu5FbJl12J67PknKccyDJijp/psPOkWVMUq3esxBA4iyrAT42R0bNG9GLYysLxikfEfUcW8kv2i
1K8eYXouUFUc5pkZFmwp1hp1JhKS387UveaqsDR75SSBh2ooFEgO3+vPL5WEPOk6aSCgJNce8/gY
T1kqowyTgN4fpaw5PX9lC4tgigCEM62JdUhp9rWFmukjcYsHRnGy7DzITjJgiH2mhL4MlGXgUsqW
2vNv5KiTPL4+PRWupSwmqeP5lwQuWDXJ/W+eecD0XbTQCDg7NWOpqy3dbkQuuE5pYz1Pz3HtvYRA
lCwBCz5QzK2CbjmKWVcrRS94hf3qyaEfgUKUbuIGEJjXmRvi1vBAHaq6E8YIHlRYp272+5FZeEvR
lEKLFsbPTneYOdMrnoXLPYCNrk98N9RTejEGULLJHD0PX/rl50ZHs+f5Qr4bvMusyBUBsWY4ud2L
tPYIg9o8xQEWGOCGHzxNzGTwVpzRbGSZv9MlKCaDy0lLhyIg2SkAC/umh8hZPpTLJzI+xv3i4D2w
at3E+PMNQavXtOr/OwKNEv1di2vHXWxTkGZzXQMKDl8VDS2q5qbOOm7NBqbEhyBw5h677jDfdKFu
Wz08d/A1t5wZHQeohpXnmXDPn4TL+avKg5fcrARF01JMe867PRPjC8upwAwSC4/1CTvDsUDKWBrB
bhrwaTBZ05ACacyrjyJpLIxh3T1E4+evNY97a4UKTPAxVTe7Z4yjhxEm4qpVN5m1yRmEvvl+63KI
525YI2/QSmjOTpONbEeuLahTar+irAF2jmzv5yLa8UQHVyYdZBtOzt90V39oHD8/5tLgXukWa9uF
Af0MSbDT4FOIhW03tGLaSaEI2xi0t/mYj+9b2VT4OU0p7rm8+W7Nl6N0eNduW5Kp8WsWc1nxjx6p
JyhK6x7I11SMwWkdybZ/ppU02Ezw4x6ocE/v0J7dngdJFKiPZq6azRxk3pBCvIMHKQnxZ5Q17Ut7
TlVJQGzw7zpIiN4k9SvbAWsba4fq1ImmjYTj86Jjpk2ORIjE3C6SEqAPbWyfMDmt3czKWa9zHjBN
5T9pLZiMLppNjlk9srF78W/HzEI3mmRRCM0hFxWAWjdvTiJ26lZOScpShC5eFQ29w3s7cJxGzp8n
TEhk3ff//PuD2OT9F7xOSndQjPImZGbsirvmsZJWqlblTQRbcvjbZ/82O0oQJUEhy8PIWS6AsWof
w4z63ml+M6Z5NnFv5eH/GqW3UP4SZ0sIWzcJodu7pdKJg3djhjkrPrrNyaEm9QkPxaTy1ervydzs
sm8FnP2Xq8HNsUy8g/HS+LeCIJPlJWk85vYsP8GgoxuRegIrRgi2bYR4DN23sPnpUJgOMGLY6n5c
63LwSEkXtxWWutpC0KQU0SZP9oVY2nXPu0ceaPjN2sfI9phNE8lvGT0tV1RHVuBnWrNBqKFKeHz9
9cPqH97XGeU0Rnr1ivtOF+1vkZGAgXCfR6c0/x9hDatBs3ozjnzFU8bscjbhC6yyCQqGFeLeRgWZ
DU3jqR92pExfweZUX009qOmPF1O7y9eAbw7BZGro2w0laPJwWB8JNqbABzU4/Uv/JhlATUqcn48q
5lBi1sPEhn1t+4rTswiyxm6LPbDxye+wTtkJ+8m7aVZ+GqFTY1dFZqZl2CN8GBEYM1BGgru5wUQO
rjIgYEAVgZSYHv4jp17aIGKIGxGcyI+72TINFoCB78ZhxtJOU2ENKI/ZmLH43u2luwHZUMKO/cnB
kH60O0BAYSaC7e/VZpqUir4VUZ244rzfZyrvP/7+R3vCxzKWz5pcn05saHRvnYMzVXZkkxF+F9Qd
RkLVtQrTznaGHfkpt3aDTOKXSbfMGZbMNyYzz4/ZImlaqJymVhjiSx2CiS5hkNAlvfFcZ3QQotHt
UlvjZW9oBNJ1bcKWEhKAvoOY6hzwFpmFiedRIo9TWj1jFJAWY5tPwiZXD0fcyX+XVWZlg7tbtVBk
y5zjTVQ77M/iP/mtifWXd7TMC5jWekz9I3GMgr+1xzb0nSr8LOdq+pht9ysirC8JrzuWk68OvktW
6DAYYcIv+bV85UIS+Nzej2MTQaer0f5W1DQmuClRWLV71H5B/kE1GDkH7xrYshXEPHO5OIRYUHaR
6O3SBi/dn/Ycbpt6Y1xDh8IadYvc1ATFAdzWyg0MueYlKf04vjZwcUF4B5asXFXMhDm8zqquPoo2
8yHiLiOOyt8+Y8WuloIvjhlMkyd/Bm5z7ZDeN5hQe8dzXVmkrezQ5CMXJjOjRkATZq8sv07J3WsK
GEYHDm+irMZBZx54B1EbsAo8xQ7uPZr4wHFexu53wiT152p65t4RiX9TbiYacoz+KWujqBb8kGL6
y+NnttY0sVs0fCUINQ9c4k+yCiMHsQZbWyG/ma8rtqQrVQ2qexb4K147geZdfazNgyQErzyrbZ3q
Zm/VFLE1AA0Vz8weKPqQGBBdqQby73EyZa0TZhzmejZvLfcmyUirW/yCBKd7SF0JpiCMsfS8HWXl
LPNuhe5RwfFXMlxzw3/d5fDiCrTBl2E8RjkPfIwBwhp//jYEWchQfpyd08sIDWhB1EpBBgRcsK5R
7hhUNJpxqvuRptsimJSuIktw2QirtGlubJvW4OdqRa/ObFb1KugOrsa+L+Iz7mF5FIw98J1wnDHi
V5gQUbJ4JZONJfjOXOZgtyvdfnTe2UBzktWbWnjuF9Fg4aJ7qgdSTovafOil6li3cnBZhC0FdaQG
qrT400L3+pd6URPIKT99AF/R0gLdQ35N0EtPhoZdEhVYjl9GcUJvQNK4rHVi817fU6HPbP8FuAVC
PUIQsE++fAn2BZrzWPmWb1eWHYVH3kRjMV4oXZVvYGorNorFj+0NXUT8f659jW6dc4ZgzUmT1eFA
HmW3RdPEpSNGQ0wmsB3z+mIm6+zSafZDcVxtIyiZVbn4jgvJJ8IAxp5fK3n7WlsrICqcgeMRYx3O
W8/z+r4ITxKZ71EjDzPJpHW0sn3MgcvWBQaqRpQ+A0K6c/Xk+GomHNKe4dT5uFOOBfF1TyXTWZvp
6GUnwQrStWzpJ09LWjwH51kKNJhxxU3q2FN7YEkF9drtNkKgXcAsZdvfqlrJTTPw3GAc2krn4TwY
uHAlfXdvTutUrAVwWC6d5uR+Fjn4ZMeSKXTShDekYhnrG4nenFUmDzLeTRIG99ygUQC/+3+Frm+U
6z+QrE+2vLM9pZ8cq8Ze73SwLKLr3gQydZSGTWjc6Ucy4Dbgxu7yssjkJ8FP4Ok9nJ2TvNPz/D4U
pTwOXyicd6iQDcOywZzj2vX3QCXHy8DRkyGh4Fnw7D1XPv6e4oelnrpjyArewwHfhkuVuJ1M/dZh
Ba85yGjshVbybKM8pJS5RHG1RGqBYFV2jOfiBhrmWrA80do/WB9yD6KBbgYj7lVOqeNCOf+G+sQZ
HD4VkTJnsiTMn8MqA+YtoPnqqoflxd7/2M41k6p+ejOnLgMzY0Qi0KdU6EBkUGCpuyjonwAstCZU
sD8a1jOOIuBHEOy0izi+UtB/Yd53ml9GEjRwsyWv1HLT2DgPQ16u0apB+SKEgPTP0XbNM/PaN3t5
+pU54MtAzSszAZxpeqmrxUjpInln/djjb+9b0BkEE8IWBI+9Tdo/UK53dt7w0HK1uuOx8GNAVu0Z
MVElyo0/6l0p2qbnw8w5cWGl0FIaZn0JfGgdyKFeWuyftIBxiWyhYCS1sY6qrI0Z28wkTxX90ege
2vTsUtWAElegSonsL2JrYxa1YxvLuCC9+nBVPMOdaGUQ4xKR0K7E5qTMfEGMWo3BCRbffWmm05iW
kFZXDB6pyOCSzf6v++XGrrsL2CB8GxB8TCcQTtWEqlzhlRc6Pm9lKDnm+vnU/lDLWmuDfg/NANLr
w4MNa6pGsvPiF12aRX0isoAmXLVGqCIdxYlz9bcXiyATPlTUMT2tW22x33HmiZmSaYs/MofCa6wG
TqxOfdx88r9Oaz3+GOOX3VlMmtlPRszioCSSelbH1MDFebdEMp2+tFmcGVbo/QN5DBhdHcYahFhJ
VXKEkD2mgJ986exYNJSYpVk5B1W4Vc2p6+U+nf6nqkvS4QUp2DLUuCnUWX+gZUiumLjDEFuF8fNK
kexYE1LI2eBpzwR0+VYdtl7Q4NXg79KfakzepE8G/02mISge1jQAvTwrDs8f2AeM4Lt0tzW330zf
MptQkCLBdiE/JD5yiFh6TKwHc9A0Kf68yEotVc/g/rglnVcMHDeE4PxHloMB0iG4+Xbdh6WdlOUF
qnuRLUzoDoodMfS6j8EcDkTJu8xjBRcHxiTzeh25rbJV78PGF1MTpO6WbHx0lLD/5Uj5rchUYSVH
D/n7LNIUVXRf2Ee1ZvIhKuk+5Ihq2tLhZgUvLsFrm2m/1ShHLbwa2Q2DamO38QLCRxciWJo12F0V
t4fp0j+9E2w8zQXBVTemUTtyzPbcVMd1tubZ5y1EEwid5N6tfytzeNBooWxNzaEIVMfl3gDRZ8Dj
rsTrAwy4bEF8aQoJca28quCAhbzs68KZSjEBvB0Le1IvaZK/HV8qj4WRNzvlifZwqMra6QNBeafH
QzZxdEYV0579MjGAFq40VELhTdVu1YYCrhOv8gLvKrXFuvWn2ETsFVkeL852hKgslUsT9x7sT/j8
9PF58xlWzUKyIHNFb4dZLYyCyH+aVV3ei0XKNSMYzCVjjXtVkm+MYZJagAulfpOMZie0mu/4IVwj
08hnS63zwTWFErNU+3+CbD9pY7jJyjuyxN3uGeTRAVaJdu4bvufrlCCTbq6CejWbZ9Fnus9bpkCZ
ZzQGvJ5a25BxT0xTBRNkIWmFIZgjQYQLO4M5OU6BTIJ++B2lFStqAi5PTIrmAkSAJtIi6Rs7dNTB
0IOLqBIn8D2g9SWRQZfhV+0Tl2PevjZ2tbNMKkfigM2wor0e3kjZaF7KwEYSUaMO01MiM0E5TmfR
6PxMwEJniW5a2tk61iKZuh2kXNnIcmjnLBdG5FGvCm+uVVeorZtfcHYYIliN+eGdh+9p9tdhBI8z
JiJxzThOUS4oDE4SHTk8lo/3NpI3i09tufn545rUNUG38SSbfNIgmewE9kf1K2RGyacWPEnCygJY
D4kreVDtH2egOxNysDrUSK/PHoSpO5k3Cc6teK42KHyu6kvoGWA04CYeNmWHpRLt4aUDmMHgyu2A
XX+GnCxM2rMUGW4GErnFAsdCMqB5rsr3eqQn06u072GNbhPtsrZVZFwODn1b9IZHx7obaY2Ym31N
Zc8wXGwhfohGsC/0H3Tj8AHNhvM1vygdUeJkeay8OotBY1DanwDXfOzMmzikgMByKvzGT7mmu9m0
diq6WjVzda6k0CQ2XkNOaG/iK0W++tZc3tO+04WD+dWA0/B6TQhPsfX/QQRRuf9lhY3IOXEgep8K
1a45WUI5X1b4hj+84jtD5wQXt4Mqro4fcg+zcjaJ9UONPYFXiXtyzle4wCiS9yEAUg28eB2QffgG
T/yZed8Jbsm0gIyoqe10GaaaZ1dDT4gwzu9YzE1wwKjIYI06dvkdtgcCAiJJvOLzk2098jpujmta
ZymR2CTjNcP9Lh6R7tQuStQU1SUHBcGjr/7yLrQ0WQO43KD8DLji2xzA3ON15qXghF43VxZD3QB9
61omnSksqCtMEQ+m5mQTemkvUArQkj6rTzk/46K6COZu18vtMC+uvnCXu+YhpKbN29XeXyY5bBkN
4INIp+A8Q9YZi6FEmeWK8w3JGLkvP8QQLhbd8jD/xRCVUe51I0BU5XrX/qbPLrtAdUOTvW8vFU6O
2t2FiGOjfFKnk0I7NDgZNsYTyrHkyTGjtRIIFPSRl4R2nLsQe2Ij3FbwL0LJdX/focvS/AN2o8FS
F/VXfKR2nQRn8CRdNgzIscoaVyFImk8DN88Ow8hHJ14zi70krYv8cbbwCXHXaoswhwuE/SAZT+JO
vX3kzPtmTaYcQVW2dLl+XV30x8tsGFFiMuAynyU8RbVC7+wDwmJRIwdE3yPld+F0ckR6PBA8Side
DIZ1NbW7XB1jYgucAaYoicrrp4AUq91pXVYhxJCLNzWdX8EKSaANPJfq1S32n8k2/I/1k6ATXqAt
9/1sT0bP2lcCGc8OGXb8N5+0GHrUL+h3XM3Gig9bkukr1ngg028O2bV8ovN24VHiJXEypVVwIxFC
MPudZ5wxiRtGD/MRuWhynKqJh+KCR/3v/fNeBUhiDrh0/ksWpbJUFxi6ocsAXbvi7+2JpwRg0CL0
spzFaDh17EgbsPuq5PnxUYmqXmur7fcb1JU2mlq6k7i1faLhi1Z5uZF3lNEW+4UqrRmVqyYVkF6V
2yFHekFUndJjkIZUGyMqeyMDV/IFdoakUG7fMXcSay1/EW3gMlzJht6tckP6rPfYHbKve14gu8k4
3YuyNXZI33OXKXpDOsUnMLmloMRoVue6dq4NYsytTJRHcJPxz9t+zBu5oU1zBNIjNPHPgQlNkmQB
INl6E8aDNQ5vf0jw0CNW7s+Tq/XtOD56kndVMxMlhVrlJqvUhEcU8B4ti1HPnZLyfEzolB8G57rT
TIUJHmw6/9XceHl/z2rB/x01uIqhMCbTnLSs5tgywiB5OpinV/Kq90EfvrzhIlEKbfHU6DdjsbSU
ET18DhEdc8foEr9gD/SMscDhQu68O1FrzTrKoSHmSVoskFrGKRch0JP/bnJww+6sq4Tf1dxH2E7F
xbI7SYFE5zngVb14cijX9T2ppbQNZHLIQ0Y63mr1FDbKaofI89PbajpdESDJgX0+TXZ5Usbaukua
OsM4eo5yzwLxH/rwNjpBXj8U4ALfHjq5aNYyila4BVL9szf23sEHsd6AnANEpVCGtPue9I+7eyhS
DgyiLB08x6mYaT0cjJ+JionYItaFt9ejhe3qA6vtJlRsdYiCMFHgmtSg+i7CngSYAp9NCVP2bmty
ErOTaTUd+rrmYU7uiUrvQDZWj2IdmkDvTCxzRDezRHWOY1FCncaj5/PQ9fWFPZV0s4prNPyJoMHs
jFHOQQbSDYakIFlyAfcp16N2LDOC0GTxCYjkGEFelCO8H9yl4qRSKBM1vATsb3xowXFN5OTOc7lv
GGLQ53UysMCviXb8RneajX2XQvYU8ejgZUoijxZr5iAmEltAsvy/A0YOkx4VsVY5DF01Opi+Jkcg
tTooNYGcuyykqY+ImKALODzKPl5i4L6zq/GJOmqMYkaULa2lKvcn/QcEP4tOshwjhOXj4n5zG3x3
U5CW3rUQtPc8bAnBwyOFwmj9BK6DzthkDZ5fK5yYjRusYHNp9vxNLLvPNEFcee5ODTSAOa9uuGvf
0jMjhJRZ3HHUsYs9vm6g3bB7p8Lucz8LKipbI+bIZpViUAn8zwjTr84H1TJkne1o1DuqIUB5iZIu
Z6vcri/NAOpEroN5bRBF7nk7TbLhbQsmW4MWALcACzysQ3SEhFSiTXpbN0Gqbj7ggFF6Y8P+HgHH
JtaSb/PFkVf1PXRoeo6HTAxnQkakAKqSTKB/bh5Rf+n+0W1UwTIh8AStBsLP+9NBNJegVNVMmjj+
/7nbh6MVwaoGOXRyiGKT9WxIbtuHLWOXuIlSO2E9tDFHEWu22IUSrZx2bqEEEAOPFjNQaOZWWTpK
ulJhDZop44J3bZw+PM1PKOKtF1EAoMQt5pHawqYm4whD+9F+NJuGrUSU1SxxRHH8N5NsJp/Zz8qV
5rDXbnHXMNuDYQ+gzD702qeUGEKJTgFYZ925+apgMhhtuUboxSVJxsipKWz1/SrQ09S1pGOk/EF6
5AMrbXXcMi6rei7DgU9FbetgyhBY2xBecAxAb7LjD8AvndPeej+DLzy9GuGzsVVy4DwY1Amrdd/b
10n/nhNZnzM1KcfAeYzEwQGgBvB4MnBgFPGPrtB1/IIU9Z6hqm9ByoE+Y9oqwVNfdGsx5G3KoqTS
act+kYiwwF/kHDVEynOleXMdi9vRJxlVSdpZPPOg5hxVaaqjidSoLhI5PgZ/E35iEe6oz6bDIu7l
Vef/UM5bPLLOljrfznWceBG4cqjnUdKwetBcNoR4OM8sO2pCc6+JCpmXsT3s2PuRSI3KrLRTtnOq
tdZK9axtIqBhHUfeEdM7PaxEnEwGcA2bZxQxrhMXVcUVZEzMN7hbcWrBJ/dpgu87iWIlefxAJgw3
0KcmZx1OYc9Airaycdq4d7A+uOmkwvaR+fAxc6taSvcmzMvrjRewOpCcrfENDfU9oUOB2SVF1qH7
4wufTc5LF38J8+gB4dr6Gndo0YAvEoT8uCaqhzR0dUwqHqEtkBgd5YLGNJNPQFhMtjY1HUfWldz0
H4F4peMh8CgU7r4nKHqaKVM2hP1+pyzFby9sUOyjkI3CGye0LFp70gZnF3DuRLOB6sCl65DGibrW
Y1B16W7YrCU+3c/PSxoArhGfSTNWGMQnhVpTP4FA6fp2qo0wj76YF0SdPoCmg4THOBisdZ8QOhvI
2n23Mw2YaaIXwWeF+X0Cd7nsc5/au65AJ44awt3oDgdH3qIS/DsUEbRO/c+P07BSqXuSXSS41DlV
0urdHknJ8X4vSQOB5ohhlFJRd7aL5Id3cbVVi2m/y4a76bYU2VWmdaUY7WWYb5z4NPCM8+7Geb5z
qJrSuyNMVWC8GFkTw4ZFLTa6lE8nj/dLwliZVRSo7H+suqvHm+Z+JvQtrpPUWRqt8ZAQRYJjyUhh
7CgGlwNSgqgcZAVIzOnk/3DKubbiPWLj5QWxoCOHYus8gAJHyOxflZsoV9+Apmj8dBa3MK3cP3NI
b5Es2JXNl34MC8ggRPBLv2thypCzzoaDGUnTiR5IuO0J22ybVnY/LZkEaZDVlq4cpCNU70lDunlE
ti/GQpa6ctRNzAv49zENBO6zQZDHMNf55ISZq2t1E4LsnBR/9OxfBsOBWYXA8N9ngAFk56QpQLpD
NeMonLDDT74BfZRHixf7TcNYD4bzptIhEivm2SMFWZ8DwI2F28UuHnSijs0cYHOQmu/+CgBE7icw
/gZsT5w5AHwFUVioK8symcRi7PiSayN2rvhCrdNc6JUfRmb356gTmHjVq2ryrfx9TvnOcg3IeGTB
kFBFwr+2iDTNg7nsyh3l769DcGXI1pcApyfSb6ZHypvVQ5l7n78Jf7Ltdmj7uhwdAJ1FoJQXQxs7
l/xaBORyMaGDrx/y+NE7zfQL5N44fxM/LR3mTxiVajguYnwD792z3E3OjFS0EjjKn7TNTThY74zP
JWq8tzO2G4hcBfoSIPpWqrsHI6jZu2PVbHVZbPp1bmJJZhXD0tHgAYB7OlaW5cqpsTpD7zPz3ElJ
zA+xTJmhGTrqWSUYArbNYWV5kbVjbu7nb/J9jXk/KndNrcp/QKhM0RNWc1jwfnOlvIty11PlHkaf
FXgqp8wWNLW++U7gct5FYOcu45urJboMp2S1onx6VBd/RbsN5q5BszxQRClmN3Peu/aCwMXB7ohD
Sh/Nr0s3SCuu2DTiAaYfNttZLB47wGzqFcr3xANtO2/+nYHmVaCLPt9fVdWeKqntcBKJI2eGHbcX
PCuqp/iA8Ow/a3a8Le+9lesefYU+4NJsnONGXITunaSwEWOcgXpwnjDsgrYLApcBo9eOfCKQWBFC
5Xn3+d2+sKOoNTfsQ/b5xBzpsd0SiCYIfMyuAzBovYgUOf8y6WPt8ctAugYBbeH+bcZP+gYvwaAZ
DUaMudamZCL1kbiqqR/XjR3oiFP+FaRw6UPe2F7r28J0wNT4yE0Ds4g1sL6wGGac+wCFQn+PQy8u
wKVonvhPCTzQtxyi5jE1OeRcGZ+FAS1HEnwRjlyr44/ODx8IFWuH5upSjsLcnncaTLUDl8kQUKSm
j02b800yQsRswEKsiRNiCM2MwDmwVFDHtoXjC5GXM+iVgyGcyWj8LhQN5HZUxgWO1jCiQ5wz2Nns
y2lybuj090lZ0i5MkTnx9uTLHstwLXUjd/hBPpxZVadP8GDt4wAcbx+622BF4cd21aGUW97kdbrF
zvSF5VTsiZ26tEElGitaY2hz3qV/SymRLZaA5L2tXhTtBKlIUMpDuwNsoSKFCoKh5jGupX24KGGM
CAYpWSU8HCLakQwIbSi/GYVNBk2SppXmTgcsoFdXqflvN/7it+hwl/lYZfW4yC7U8RI4BxkSMJhu
spnycj3suhPAubaVdGioMI/tul/rpxFzrHs/OyI7EHJQDjDPNkb/GPA2cfqsEa6B3tRGIst3iDy1
fiMbVa1dRgYbc8NGbabQ15vhGYWwmcAjdndLlXFY85nuSCQbSN4hsgKfPUZ9gE3oPMuXBqvp0YGc
jUT3yUYUm6SZhQzbh45cGozb62JQ+DIoADRG5Wrkj1Bk9qLGt3hpniAS+aqg6ih71SaaALoroSQ5
VBxauc1Ff+IW4nEJsMyNn6eYtvU6Nl2pCZffIW1jESpYBwxoe1ezlgSVSZhqT7ammVVLtdG9p9qd
mCes2HvB+oWTHqdRannhHhxkIRqKygt4bcGfXYt+T/Dv8KYGsFEZ2Uh0t6QR710dEGqNrbbeKC+H
HXoRka4PXmu0J+8SlUIYAVS5PSmvkSGt8/fNWl+gkHTYwXSwJkGn8xgtbISYMcl9keRDdFiTvTi2
BUh3CK9PS1tbLXq2pBGg9Qwe/nmNxcbewqGbRI2/+4IUai4IH2Hr+tlWmEolGuSsL4VhBYd2MEAz
+eX4LqdyaTwIWDP7g6tGErdheGyHQhTN/FzSqomHnfy+DTOHmoKsiH0kj9pwGr9oi/PGOxGXlRm4
wnJ8tKpVdbwegKx21gFeohbhLWkDwnMFComV71/SptNy0IJPKyGW6bCsGsDFwdF8YUczCGWe+cta
pg1CVN3xWWFx3zMHbwj4vd4//A21H5eggSivE0VtBwTiTYCP8Q5sFW1kFo7s/L3dIyNi7a+Xzlit
8TKELlMeaVKtEBTz4190PxenXX1d+9oIBwaDgy53p3bC1uW/yMSsArUxoAlPh3/sCpuASn340QCv
X9BzdY8ehMB/EYNGTrJTyVj9lR00X66PTq61wKYvVr/KJNbXFBzsjndGZJPaw5/qOFT5p5xfxef+
+oMKs3/HrdWPOKzH8pOMrjMeZdsFfWCGg2OnlPxkALTrNQ+FCpDvY6P93S0BKwa52KtZhwX8k7Ah
OLKNTmTR3Kv9HqEAB+4D30iaVqgDNIUT8JpvUqwZvbApTGgWhbjz27rCzO5YqPNJ78kNlO3cDuwk
E6Dzlpscv4Zq5xnvJzc9LCMdsQsSXwKM781FCU5IRO+F2V5fn7o3xMRFwn13wEzC7KZE9TNU5zJ8
3DANeOa63BFf2RUShYAogntHUeELUjhwOmZyY+CEMF9p5YXMwHM6gNzVQI/w4FLDS0OKrxAziI5p
RcujYdHzZN22k5puvYsD50HkDK9y2dNLsTMToB8zgqYXU58v5xCt4jdxGioFOhoHRMW9JeBGY0yW
MkNRmUyK+K4KPVhgLCRjZPOs4aYPdkT8HWeDfjiTtl4Ss4GVDib/yNLvlNhJSWEIuTWidc0Pa7+3
F4aCSHSh5wcj5N/Jg3dM4tPy3xqr5UoPU2sI6/YEpR4i/M+6igZkmFwXKCQbQTNELiGM6Df9/SrO
eu+eX9Qr9FMjYpqKrvbNwhyR4B8yIkf7nUWyLuKZx7cV62zn7m39IXt1G1hVzH10sbwcy3XMp7ZY
RSwvq46E9q1lpwoNA7ZPzpWs3VTA8p0Eae5XPnRJeZCfiNnpM5ElMBHXj9KR+WO9m++mEQCM7FV5
7XYglHXRBZX8SJccOfr8pHV/lZTprDh2eMNTTMCBzmqFLVBuFZjgzslDNqw3gaet3viA3CJ7DOB7
qiP9KgX095Ip65lZwacW90AcJohF9dcbJkSQ67JfnFyowbG3Q6S5EKrCvslwdlpxAuAJkL3waBb0
uko2oP9QrA15ooJVsqRhQwrHh+zQyRs4WoKkEdXZUrOP1Jb5ZWbcSdglLuXfq1cjk5GoMjmIWPa8
FOQyeda/O+uyCu4NBXNQ/ZKQECZc8rixAbUL2bgbgw1eEc8ayXOUHk7ZTJMGW7uOLjkLnGL13Pr6
K46vGguMfXN60ePiFvM92FrKHqrlNK4+UVirpus57hX+h5Tgx2aiXRRFmb9iTt1kF4jaTiWwXpgc
G7KtWTzvBC667tMUjHw2zmOtQvdRNOmsGHUReHMZBT6G50ihHUfAdUizPCEeloCon0p7JNlI482+
IG+cSVAUFcjUNGo8O8q7Zxt1D2Uoy1xEHkIHBXpBkr2fMotBlKojy/Ex7l504gvWj7TegDnuJ4tH
mOskI1lmy45WROzpBw8g1A6ojZtyET/SG8qak2zkEGtwtdy8uaG+22aCnbHV5h327TkW0Fw/2UsS
5mudIL71gQJPDpNvUm79qGRlavFT9DGMqZIA/j3Y3qAfbaXp/fbP6INO5mR7yxOLCk8La/f4KrdX
1gctBkbHcOpkY94xKMuWUrXJXWY+R41ycdJAiYDUg2pGGhxM+ohWlhLCv3GgW2aQF4AtLX/5UIe9
RwagoV2MlZ5PwugCwOST0VYoOAECu4tmEomrwBXt1H5uV2BfkfTu/mzS1D44PaC+fHId/dNRuGLr
aAPHzpOdaMDGak+L2G8kyvamw1SrACZUd7tf+4iH2Pah6BRX3ssupda7AsWW01e9D7nj2G79QqCZ
xKWSVKNJWOHlrLW1Bi7+70YFRS5ot7yeAqL7RtRyDL6ENR/DsPkBnutt5CPzCYyDF40ptnr0vXpb
p3Biu6nG+wnRtfrU7fou7W/p2LYItLq4LgDp/NtUsvhipA77lJgEOTrudfytXx3ucdLAI5jV9rLs
9CCeWsweN7OrkHevIva0Pih5pO/YuXjR5hlbq/z1r9Vj8diZNVFJDtIoB6uIwox88nytkJ5QW51i
XtFyy+xooBK24hDx+bn0tC5kucAMhBPULJcKup+vo0VrSU0NQfsuzklIx3vK+CotyugzLtjtug0s
j4/beQDqmhN1qFtjZcWG6erbskJKtw0GIlOrPaMEbXbAXBGMSXcNfUfE+oCZXGENTq5ArpB8WQJr
6ncmhqn9LYA6T5xcxCXgDxMOtBQd2q9XoJTnVg1U1QLqtiMcEPCamfffLuFOU2FL6Q8sxkVDHfJ9
TqsPhBWvPRwY4OKMrqWiCNn59SXb2SrCOS0v6/5lbdXt5JriOvO7qoapvrvkfg6fW1N2Hy92icP4
q+aGGAxYi9kvWFZ08kv8/SWPeI17gVAare8iHiSCkUxRehaLhBnvhzchl2PYSAcSib++TDnAFMtA
Lnr+MB+4inbCTlr/XRzs4d9JyNukpJak9BjLjCm7aDEzUUsxmUS66gUfkVZeR18q2n8SqcMmsl6h
GYGrnCpL4NGel3Z3jQjP7NuGzDvDMl6Gwxe35MJExAwIFJMP+uyTvyVVRmI3MnULk/JGnQrOyALz
jcojJTZVK8deQXLy0HjK5R4vQmxkF/a7K8ytKNzg8XqjONWa6wIfnBoss0KHCnthuISjvQWAnfYM
VDEn5ZYJVJmA5pDT21SbvEI57gaIP6aV7+1sI4Yqw0pBcsnDdiYpApK5vPLnSgiN4OAH/3PHW533
zhytW0/1OonoVIlkV87b0jWAu+TRb5TaQ+T5H53ZIoxngmxLuses7N//z1TjiOm86NgkWY15G3PD
B7gegyV7CrUZ5/GEPTE4AlwJE5sPtFaxRysr/RerPLpGgKwVFCxV4uipo2PCREpzAwigL619q6aL
2ILLZ+HCiBX0OPc3t237AFKJAON/0ROEfuWawgUOyvCKwxYkxIj0G56twCFgFSMKgg3DuLHcCmi2
Ie9Nn9WV6uOK86ffU5IFrveXVJYVCmKaZMhGOUPJDbXwrYV77a4AmR+sGuTHt8eBrXEnBSA6toN6
pbef5sPISh/vc3WUWflmCiWYj6QRfSvWtb8t7+uA3o3A0XE3PHasQD1W0IJL7M6U5ug/zPIdQpQK
sxmLrfQxlVY1iV3s+VsTh3xvES7BkH6dnSHVL6udrSzYjtmBqepSCy+CisodItFqnw8HGjBcOKnc
EOZknzfwpgMHUJQK9KhahiIfED4mzi9H/7290AO2RM2E5mPSO/IC7/spcbdb+l0IrYpnln7m2LXx
Zi0CVoGU+ud31/hcVdhtGUlAsz1jLRtzbiVDCGRLt7jcSHnjUx1YY6oSEpR9S/V9KHPoOvhsh7rd
UZ99o9dJRSHCK+l02z/XhRIj/URJ7iTUtMRtaY29W7tYyEqJ8GeRPtKwIeyNCQCtfk082qF2XCHF
PlwTHmPo1nnttbe586owZMpIB7B8AtO76GinujMiFoxZ/Gm7rWj8Ra4gW+ulAzQ3ucjcTBOs+FJc
ZCgJJO1QzvzWXnwVO3j8vcnrm54D4oZUxkUfGk78Ja6/qNieXnUPkmHZsh7sCLrzB8sd5vcBskgo
Ui88OJyGrIz4envdwOPwWJlUtkIhJNYnvOyxRDwyRsEcwLRGPDHWQboCdKzl452ntVQQDqpdC1ep
kflWzavOlqbgmQMEsAnKYl97Z9sYfQcidV3Ba1lEFS2U4k1GBBAc9NaqpjHTIP72DuWuwbWN00gW
xk2WplkTl+vHfNMQW5Sx2Up2gJelw87K2OQ9i4LmmBfGtk2wFoCM8vVQpeUPe073gBZWsfhaLZdV
vUfqYKbqaRiwjFQ7xfOZ7t3nFtqtvNwMKylqdgLYD/f9yWSOYd28sXAo8zlG2dvMJUPSym+M9ZCe
En5ce6GjyImGo/I/kM1ZLrXSeX8LqJM0AeOieV7E05H3FtJh56rz9VORWa7HzFRF4xb3tXF/4o0H
3WFUul0AM8EoR1ap1DbboAO/ndqdWWAOn5IRL7modYucFJfEtu6uNO8BcWMGbhQDcQPwWGDCX7Vr
frkF3FXHde5zN3durbkmtCLxejYO2e81PYbdJWxfI6pYEJ2yljkisiCZ58sjUkbehknzREc6tTC/
Ir2fN8yfbIqv/LBn/D44WdYxfGNO+N6HDmMSFNK+4EPYaHB8Xl4u3TqMLTOq+epXuPTRQ2R0H7JX
GXsEjT/VN1rYIFdy6hXJAfW+HY6nyO3EiTL76uU1OvqXuDenfZW2UlzYA6mIcC8HtOqV86yBKJHg
1xPod0OL84Nsw2caJxDUeeONwJJS3EWb1OB+3Lxr57eTi1T34Y/eZ+GESXmAfqcl7tRP+vNOYLdV
afbUfQMQYWF8YUM+zxJyuS+sWFuE1el0oaWmvVhbBG5ESsCQ3X8Pw7dtlIILxj4jsuvAGZvQooAB
nYDjOy48pRvn9Es/FOs2wGhruAWmGs/1CYSOFIWK9isKw3jbRHK6y3OYzsAQZf8Ei9rRU6LspVAU
GUvp9L+4y5raD6PlQLoq+wp0sGAb4r2ofzOCyPJ2+2PLs0tN91rdSh+FVv7PrBJZeSuXjfmBmrv2
eFpUlP5eqYig8kEpp8ZKEgbBRsJBxDCl3xVrikbfK7uLtHw2nbBjRbiMmqiXpxzNkUZFdJv/CV8w
27L1Fkj5lXzH2F85bvnfIaP1i25fuxj12FZe8+OuGsURC6OFSsXQOq53Oz+7MCEbkPUsNRrkZmYG
L7ohIhJE7Iz0/wDgqJqXk5ppeBxcnDJ6sP4jNp/RooCB5lSWothflkKZw2ZeLcVDk+Rh4gTuZi/+
H6e843fR8aq/HE79DxZU3ZgnoX/cl9bsPztKnWlL26ofRujmjYEJwCZm+BKIdbU/qSZNnZ0IkylG
uvjOls7HurMGBYq0RBWfn5FqlUQiueJR9B1UVGKVaBSu/SEKYsmO9GJ9ihLWTbDLDlTfm+zxyE4z
ExXdLwkqSNkWnzjbjWeOa7C7lmNhOYndjCN2jXTDfzvzUeMcMxpiur70pnYdG2ej3Bd3YWqsnda6
+Ufk28fUSuGchmCEwUuQJZr9V7VrU5LKwtEU5A7FqHcx7ANeMEwMR+n4BlwCjZPIuCkYYk5q27Iy
7H1rA+vey+03jiWF2Gm3+/rBtCAj/ZoPxQ0lBRftsgRI7jW+Z7O11I224J40tSMaEHDxPoLnLTYv
rwCSlsG7oHn1NS52cJwPOQVRMJmvuwSc3why+MbaAbcM4kAF1mPZ0Vj02VNWXXje4hh1eMwWv0Yb
t6ICfjwgHkV9PS08m+cfE2UQ1rwsaxi2VFGbcZytI5UxXrknL/GbGyWHL6Nkt/l6Ylax9gkEv9/Q
/ONb9EQJZQBnCkk6uf5nAm3NRBcHwLtiT9qXru1cJAttnpKTWaaIoEguftWlWLXztDs/7CRlP0yJ
985J4dWfylvBq+VCDNiRfQ2lJ15zs20ZIfCGui5m1sZcbsiH49mn5w/ekulesALqN8kuGbhK4g/C
QwdNdlyD0Wwea6OOAnjGTc1Ttl0PNHHq42DOc2IZxwjrKfx45Bw1y6e3OyZnlLMTAXSM6vGyjoye
7h6ElXmAZOxXd7mB2OVXmoWJp7uLvuk0JD3QnzIyFmK9jonG6vN1vOls1TnDnl8vqLQmXOYJC5cm
xS4J/pE699PVw6tyuBbHrjvTBWNjFQmi3vUlsU7jCoaRtkbJLEPteTalxH0b1RSFzgsBxKUpDAHP
ofQc03DTLu7N0AZ1P8CEvo+o1dyfWqo+OyVKBaoOdoXqFZNjq5WwZkMaTQJocOrF9aC8LaSh7rGq
HWzxJHapKWC/Vq3N1TtgrSHL8k6xCSu+WxSsortuYLclnpxYVEluWIZSrctNbVI9ZnoRYAczx7N+
VDM54rNz0cTF3uORRKwn57wALJJ0ZUhb4i1T8pdY3r74RXuz2I7l5WLtqUeWAr5b+2CvRol7FYaG
V4nxBf4DYjNbQmB1SdcTcfdHszLj81FH6cpsGdh5pc9hgQllv3s/Iy5BZdCJGjUyrN9k+a36Ep0E
37xSYloul5tWWR54G1lqQX8iM2pYEIdhm1rDPP01DUFbFW9hrIPHt0C+IgoHRRDSBFQfLruJZy87
3vZythe90Llht2pnRVLL1e1KaeZeNKzXxGdc958eQQm9GxpjvIN5p8hTzo14hZSfEWjPo2kSAClL
anDgbh32DL0zILcgsSpdkDK9NjMpR53hEuTmzg53cMV3L8eR+mILpznKUwB7kUtwwdxlUkfeuWa4
KPF9qHJB+DWxYMdF7TrNE2UMJ+YreTK7lcHVEnnJz/BMp9KrZWvvEOSsOwuqjXTrasVPLoD5rdIf
zv3ntGE54KEflrqTFZCkjBAiWOvFznMTVZB7ubmd4BS6vuak/rf1HepXqz9FNgGW/wjynRMRxWYh
Rre10GDyL3HbUDp219hIGsg/v98/5u0zlvJid8LBtEAseR4mYuF4Y4dYqBWMCcVHgkMslThjDCjg
38RxLMG6wixKNKiQPQ+Tjmbxtr+BKpGxheVdRTSq3lVVRiTw/bse9pSPO8vqhhTySHZADQFKhNhX
zA3nvc4j84NoiGv0Mic4dUZ0htJ9aqkFiB81PRo6/Qgh4Vunv61WFmav7EvtRYDxD02s2BALaX17
Db5+drcYa5pH27bYDyyo6kB6vvhOaw3zG2i5U4YiRxQYtKZe7cLhRPkpjyS8dijzehwUMXozwysc
IpubDa+m2nhXisCvp0YgMODxnDTtRUEkl4wF82uR1/PDSoCNm/PIZyynFNAuOAmkjAE0G8mmb71d
HVoilRRHKTJEe+DpTrArc9D3MfDYlmyBSEBatKp0AptZOhyM0cgWCoMT8iHNLEQ0iGBaC2+nC8bW
/FWQKPrgWa5lbxmr1OHfUjon4wYNbqChJLT2tNwNUB/96mrJzaz5lAFu3A+pWNsjAcHZg06TzE0P
2TuCLXUbc9DuKj5wGYPlDv73AfSb0x+fSq1VohInJEUrC/Hw9Owg/rMlhIO/NArjrTKkhDWf/x8g
l9lqDTNEU+t5myV1TnsDAypt2hDcjwj8x0iZZM8nEU3sm9aqMOEYVePeN5Pnp6RgbFvFvFhn/JJL
KNQljQHL3geqAQYy+9kXo2cS7iT16DykTa3WTaw2MAqO8bwismPY6WzYN18gcHf/lsR2LvzgVUim
E9zXBSniDCo7Sd12vx/Z+huvVTEQU4cXg1Tc9J1KFDTsl7Sco4Qk119pp6KaSDEAloTVeG3He3g6
6TJZ5IiM34pVMhRyoOdb7qvIdeTSuhT6o9BWMak/s41boFtLzSNoeAk4ZdIo6NfyO9QcAcmOrnE1
MkeXYkGpRmW5Kv991WU0zdGvZIedTM+hx0Z6SwQYCJO5i6loyf45D2HdCba39kCH//Rkrhmx38Jp
0Tj5EXlHkLoIMIEMji59XXZvvd4KyhWGFFob/tEli0hrkE0tTtO9T95oHbluKUaP1U1IBpGPOUpB
MK3L5NJvQEhJQYp1x/3eg7Iy7Gk7BsAaLu5kndjCEPavON8tNFH5UtUknPEQtuHddeTV8abKnaZP
1w9MzuIAlM6XxX+ZPjF2sHGkBGE0u2Z58mzX4BoOiM8Ok9xrNnHxaZ62L9wz64uxoPvjygW6gZFI
Ig2Oebxbiqd1YJYzwPKRsl093t6hte7fan63DpVyHVzcwwtoVpgMPcLD+vYyJMg1YJGrGQFvBr9i
poHqeorNBNb/TWdYWzRmPii7nDBjas8Su3Uy4OVCUtl5LZoLzmqhiq+7+pSvchgH1Na7+NA8IBHl
gkupXuiIDelBraAnXsCRN+pFmAewkSCOJ4TyEl5EY2PRg8d9HCSKhjVQuicTScwg56HaZGQVos6O
vzc9ak/B0tuy2lCAXT4F5J+n0uquEQL/onhToNrEPRQPQnk6KLMteWbQX3cNtEyVazd6ldZ2uLw1
f0/s1qcOyuOIPV8QnM+dd7qrbZp7NNi8Az3R7svFkFgZQC/0BbXLaYvlqQXbb++6mfLPbnY65IB1
98QTKuh2e2i+2BVS2VQcJP2zWaemMK9XpiuJ8IM6FZ7tBFlMZR3yi67aIbkcsqmpC+A+DN4wEd08
doM2TTzMGBCfZpk2dglqaR6qslsMEPa1snPoWwB5Cekqp3W2SPoI6qgUnbNlkcUC6VBVOpI7pq88
seunnuO4CsYr1a8gbHtYxCCYiDC4gOt4HDgBXOmLVdhstX/x7yqUUezWq5LUXBigCD5G9A4Bz6Ej
WGwp3Nxzne37+UzLeY63DwbvbIgMIXeL80lVsSFRPv1KdsgJaDp1XxyQyVgB+rPqmm/m9PNOq4yW
jCexW9eihqF+nFvhy8N/zELajVthAhXoSoXyntI9J2QHKFL/K7NsIE2Jl0MY4fotte7s89aQeeMZ
mJ3Q1iowEjvPCPKDF2GumND9TbEnt+QbWC0uKIiGq757gjUsQwHpXlrnn+40xc6KXQj3k+LIkMAY
XC+ZS3kyUL3Qw/03TTk0VjlxfhiZUeNxSZhiMKLffU//+q3TmEcQuwlSnNhcPzgCkEr1B1Nq/m9y
poWm3Ck8vWGkN51JEJ5giX65xt97RQ6tYQHt2wWsc6mJlC5tgDHoszqVNt3DyAVSjYmxw/9Hl04v
a3+6lvuuWmYGZgEh9i4Q1+K/1t3jtX5tlTfGvSFJsewpwZrIBinwIrQrg5UXkcj/8MTZGbQwhyTd
tPysrN/kzFvD+/+M5fhndnK1davqkw2BOyMcSEDy0H9ILzYApwposraOnTeU95Y+NCHPPrvlNxPE
6QnNtUcFAJjuUs8W7rvU7NkO6unnl3Gk9jchYdg32YWUVig0MLGmXfwfjBGMoMhATsgbbDUlkww1
+K67ScTAVD9gVn98ShdKd6j4QFYUG3yDSGor83jMOS0yDWC0YLxKpW3vRpDSOcV2gVoaxbBTfd4H
m3GX0Tye3Q55pwlAuhw9s1/ypX5oJeaOH6R9rAjpRnRPoFYZJxwVZ4zauCEMfp6t7WcjwtJCV5/M
/uM34+ryYkPTGx+sdxPn/d81I5RBy1npP5QGJbgJZc1n9zUGLpkrA1bJAXPF9kmuwkZOxhndphXI
n8hOQDnlMCZ/KIfUCE10nq8yenfH7odOm2sEwXsMXYJH30uxJgj275ugejE7ABzEKv/mN0sNeL0+
vWvlFAR0KwkhNoXZ2VskijlJw8kRahb/PNr3ZSF7phx43UEa8grutz5fCTvDUZFXe2ZGCcex7GGm
eQn528C77iVCSe+NGzxCJzFnWWrhomayKXaQ+xH3ie9uGp7yNMRGQfpNiV6/rZCfTulcucDKjFd/
r1P2ovKOEMVoTFyTskl1l6c72Q89LXr4e34qUTTszFAvjsRnhi3l6o8trQb0qKIVKMNS5h6dPgDm
r7LliVdxpy8rRaCi5a82gj8S1TBaKXB5OWW9USTBuKSC0B/SJWZt9BkaQB3AVQmH1rlRxit00TcT
BBoZLc+ytUXTKaxUq0wM2PF9KC6SFVsD7UXF7PTHj98qVgssClNTfHiueEursxfYLnGddq3AvhiI
xiHdxNlNEAnbKYuWXykPkwp/MOCDMxBZ4oaDFCb5lz5pEao2lolOaOcD+vJ6SlCaMaoAUcJnl6Ye
GUDEF5sGfV/BG+i9LAJE0rUBT2O4tXc1KMsaj1/u+Bz2xmYMZhmFni4NSPqHUhsTHTbZRP6no9MK
EUE1ZY9I8M8Hvt4foQUB7LNwu/LCBgGwLsAjMFa++qyfA/NcREPpafwRFjiWXu/rVhM/B6zylCA3
nm+SP6Mh0lEgGCHXOatYIa17SmY6ivW4lZYFnIlAmFxMj4H3gA709Jqd0cUXtwQ2bWLUQ4B1XR5R
lTS4WxMJGnz2jHjlwycZEdHll3XuqVO37oAbjkyaljmxSaqmWc8ODO+gybchU4vOVkiMT/N2GZuZ
R8PUCHzPHq9onHjtrJbqoO08IuEMA7/wUM9yNysYjmVSymw71UogW7GSW9S8v2z/vPMKcAkGDC0x
IBJXzlDCKhne0/p9WOFgtxbzHKpUSah3fejMeeeUKLT99QgrInmGPxAS+uk35f/2nT6gBNuiNloT
kYxdWvkIzVOYIYWoqHFFtekQMhgBf6d8nEzOLKsENqjvga1rCb657txQfpwNlhFc2L7yo5SJembT
dy6uzQcyAzMo10HCixwEM/qygrsUJAMemuvxkbH7M7HV8JoRW//fwao5BqswD9kyzr4O6/y/fEAq
dv2muo4NNw0vv97SIz7hS86YYT1J/oYrp3sbP34ZZxtbqBmsrw8jvYgrTifPmy8B89j9Q9UsnhmW
8jWh6atoermlt9dp5DeSPHh5xc2z98/O0A6Y9oj2OM2Ddh5hIxF+0PTfkzyrEVqoSkstfwDop+CN
RoZvngotfspIIMzG2jaj8E8IZqjZbY5QIkueLyOArqSko8b7r5vwEIsqWKbZhRdiRIZqPgIg2Xpe
ErLLkoOiniZAoHJGuNEkc3LFNhQgORQh5CmzKZkC/BJ47iqq9+8ZJIcebhGfgZOlSTBA9AHLpv8K
L71+KY6pN5hu7WsTvIYiXlyAHNLJp103S5uoHy3g5DP7ZWJnn5+EhfXWqTeJbfC8MFAcVsU80DRu
94NEt23t7f7VucW9U6lsYCqlpHyiEOKeXkJ0ESC9teYBSzbVaolUOEXUoYIzSTiH9D4nph3Zys37
sH85Ez12oC7ZJVSF1KtdQV+j5GruFVqWfrI7psoULn9lrMAP6s68dHwURqeIbwE4b1oKMFK07w2Y
3r4FSLA0WGpqrLcQ4RewRxdaIKq7r4l+zkaszcJntX/So+tuNUuvHxWlKiuL3Ss7sXUNgwqk7haB
SaWkJz00iK5kolzM6ulmb+JeLwbbANLTmgllyP+SOUncOh8pkLp7vDu4YhqRlHzMu8quYKNfbB2j
XD9dkH95adbzw5MUCjRk9TMc71F7jzFl89OD4e9iTBNxi8rtYTF15zVPUVuqQFrcCLsN9q/EUAZk
gBOELZNBTAc32o62OSVWEjG1Z5Zm3bctEMnX+FFBj4TfyZlfPa2MsSWcvZH3U/hkRnUAPCYsrGzI
ahR9WibFFIuW5rN+ShNH+bTPhLZCNGeUwivps5xpvHtAVqKxCRJBG507as5keBvL3tw94gybGZS6
uBm7ZrdI9Phfo32sMFk9Z5Eueq/77wBRRDVCcvFjy//gcQazs9KE87ySzzqh5W6bZSOCWlD6LLP/
1A/FNz/unYbpY1HosVTXbR1W6WcyIcqIAi46CNLuXz7WK7iWA0DFTqO+ZQTn0Zjm7I9eHkfAq3Ha
eZHNmqLCZo1rlL/9AloVqFNvQj7CbdLM7VoMJ27218kZLtc7GmQix0dPSmiGjcGFrqFVuPZZXTjk
6qBnqRIPGSfnTCThOtGj2y4PhCQp5F9Rwv6FhMNiwS0JyaJB0KRBYnmi6twpQ5wS5RAXsn0JaWu4
8lA8s6EcDMQSo+60aAyhwsfi/areVM56Uw6dm9GE7U3ILFa1LW1XfBbzjeXy2n4mDBh0AAUYjK4G
LKkNSZ4DfkVNerT+qNG6kWYVb0zd/qNWqEUPfX9hpSO5jf9crlA4frtMn/QnFiNLp/nbyuq9Rlvb
v+pzm8EaEOSRMfEEwAZrtgMzR9pGRwbULmjKeATbUSvQmK5c079mejhtiDk+n1Zn9xtnAgyyI1EV
ZjuT2RP/em4IKPa2cR7lDs4Vqz1W6qxy7whks0vsua0seFFF4hM0ZAaNLxivrJvzsyG7YHwZKnJM
NedmcQBVVDHDGxCrOvccoaFccMAJvUM2fZ4VUmRseVvFfRVHuprG/DBsVtixbHLvrkRRKR4b5RiG
ZlJzbJw1R3lCV/W903XjFeEh6m1fQGF4ktnlw4Flpnjbqz+Prqq/UYNkoU9eiFfDIVa16n2uqZDJ
ASQKHNcuABl27Ftlk2XfT6Fwd24rWIsb3vqt0tQ6hcGi2T7+rnuKDnaUzei7S8vqug6XOMED3zy4
Jr5BctaHnXuT+YT7AH5+PXbaTb7WsScGI7TFmHT1dJ5wzjlj8tzulLv0hoNMWR0WwBSu9lk19J5L
Ec5LjUYsFVm0DgPmj6N+AbIrybgFwZtSQmaXNOHptRVyFMuTB6+boODRyH1X1RvONxAMinaL6q2y
yLYkxIOyfeTwo8+GJt7SDr2tJEfU/TGT5HE2h3gb0Xpd5HZIBmb4IHitt/hthiT4OuaWQRfgYvpn
KnGirdjw71hijjoEJHnnPSogGAoh7VvlMruwSahxBiTcGbAqsCeipEUGOl3ZtsErL2XDoDlG66s8
Fdwjgtndg3nafBwUuMHAzxjsYQo9S85GTawx7TPezXuHVC+hbk+ZAh6KV2DfX+XY4sndKNfu82Uc
nk29IAlYnVawNWG3rkCLGgVZg2eosuJNcTRIntJjN636px+b+HY+WTlrWjx+2RRUorZZ6Dw9prnI
zg8Lz7Rfl3tGrA5n1lruMYDFsL5kML2dRfRW8KfhJ9i3TPwWUL3kKZQME69eSqw8hzw1zjmcvThF
Zu0ewGXiAqXQHgOxn3Fd9IskCxP9m0nn9Tu79PphlDL4Bt8SRvp1fO8wQ++BwJKfs6aVk3Lqn+DQ
TkwQHDD0VNXnmMVlJzFCezYjPCmAG0q3B6ausiclEUfg1sNRxmvyj1DoswhERGxq+BINxoX5VR6H
9ntag88nHAeqoyqPiTEW6OJtDc9Vsc7qXKzVcbfJ7wcDeNqX4nBuEuN8ThH9CDLKsno20Q6C6pDk
gt5N4bd9wyTxL7w/G2X9/xbRTzWq0jIyGD8vN7chFj2VGsHauNlKHTgodgNggijaxQodA/rn0tkQ
O9oOOgii0z5snvXpLPCiL6HtzaNGde+6ksKNfD1uKiepTZ4bZdVwEpKmRVd2XC7be94KP+WaWbhP
xXmBE/698lxorwikTt0t9NLAE72bFDy9FYDzzDkbvTlwkxoJKR9viSNmEyyiV/Lct9g+15HG4dmb
GSbXD3KpJSAOe9ymrW1cxGKB49m6ACXgt37rhkc2EMYWaJr4CXYTaxWAIl0nvUYx4mIkNMYDSqcv
L1pZ9uEf5PX95e4jkab81jOx8OcZCca9q68YwlBrB6vxFl+fABfzYksMqf57bMt8fEMIKvx510mv
Z5DkITrFYMxtKQ4K9rOU852E+xLxQiuTBU4pFuDloqIg/yzqCvgr0JZj3ncaHPNsJqrG05N5e8I4
sVBLkAC0PuDBHko/Nm603legkdhBmx//6pMlc1mTex9k1Ih7nGwIXcnqEJUPlXO1f2yRoSPdCm8V
0gVMFVAuhDmZokNUgJ2fDfAGyrKMUjjBloYfMxgsb2Go5XnHhipkVLpRPfuh/BXi55cHDVh6b2mH
QgJpGHWEA8LVRlZZy8dNAAoH0o7ql6RNwt9eLNwRbkiNBHwZVpTLpPcK+WGQUG0McuIGBl1ka/XV
tV/hn65SixjrYf25GJyN71WX8vy4hbAq99C1NER9Vnlv9xnVDAOb+bBRW4JerSB//L16yM0nO3V2
N3c5poZ5sFRmrHRyHxw8qQz0bYQUt+4b5FKr6hP3pLcGnklkxBdhzmUpTTuOWktZG2Ud9g2l2MAJ
TiPoX6otirVtK8uFzP4giWBytTYH/Xfdf8PDBXJDtUq49sKXwbCLayPyQRPTrDSJ3kvEiS7W8XxZ
MU9NB50Z2qjV7c1WhbiRC+vFbm5oXfUgkF6lUasK1BaCeZXCNpkASR7Dvd9fpUKPLHn6Wan/zQSU
6tvLpRfNIXPBgTEhfcVI58vhUcukSyywqUkGrGCfg9hJ4BOdY+UiYTsKzp+t9++sRGeWiD7CIELC
KR3iA1mn7py+fDAeA5rL475stgbj4oBbABoTe0cwyYGeI2svLKSx0dnagSL+MlqOsN+Eoi6a7XMh
G3dq3fonikl6BH15hPc13AOsCuwwHkkkIdeBErqdrzzeEPelpEXSRJtXAUpmAdWlNmZnvWsFUOIu
W4FY3elnhWnBgsXW3PzgEf7cyjz6JvCvfJ7ax9qrYa0ANZKNs7lBtbTB3RKHEkPv5JwGzqHYZzFh
sl3w6SYzQcKoW8gPcyOpdKxFAfTY/oduKIwCePhXmFlA3UxdlMeQJiMkNP8tw3zAK9JrMkmK/Z6C
A2YRDB6ACuKqOkHz72fBYlkWH8c0UQapjXtBiNkzlAqc65TTLNQzSfQj+K2y0jdQeyq94DPSrYYW
kGz0wVmK3lJ1g1P8LkqsMbnovB071GNKd5DuF63dAtb7brvn1w9zdG2XYOwiFvX2NKNeDV5UNkt6
pozqJUUBcJ9IAbx1HEd5BDOs4KDg5N/WmThV5ZlQTgY3/cUGc44VsZZK5ZhyBMr0LCBJPNZxigKt
utC7Mk0VCn/UMCCwJfEZmqZ/1FEAD1Z10FSqIqaWh40U/J0dp2nNrZ+t4IT1kn95VXBAcNxlHC1M
owLdmdlMJvAupfIQFse7u5lk2A4KMGgSSaufoU147iTKtiZ0soltHEBeYDzUKZYUQPc9HeD89qnH
E6jMUPx26vThzr0ZEiTlZ1LIuEt12YV50NWbC1cmJXYjl/iJOF67xs4RbnNLwmY+Io461b9VOnqh
0Uzx9Lk9RatcwQdv79II7yeMpesYsprafmUX1rpO/DktqSY1I/iEz11fMNAxdjp+k6ikt+8vT4pk
3xiAqjQTNZhwEzIPn/pW3zyCLMRDepUmY7gOTIN5ye64wMn+iq3QO4KTQk0EIUpEwt+iL8Iwt3aT
y/ylMo5lsQhMmq1vdv6Ef+pvbKcw4ChXPnQPUKf5gBeXGYXIieE07b9FeimTh9VhBW/aUNbBWLNt
nK1QLmAd1qH8VxEwdZT7vOiOm4LEzDjTcEsbB+Ye8jJXAN5naucg5Ey/ccCTYVPQwm6OS76V/uGc
+ZBdDqXi1za9j2W9zfaC5vqKUq8QJmdi7LhYwWB3D4DeAvbyXcLpR4xxDIBFNpx0dpy5RP3fhWQA
K4cSpo6drtTMx5OsgG8GTevahZl2B5GL5690SxTPAEaAdrk+JJ2YOO57RtMwA5ZuDbeaQKehyVh3
WkcwwQcTpPgAkDzlhSsee0iaz8HXRx55erVlwupgyBg1C3ChBxOIkMvIKAk5drYE+sC7ms3tCvTG
fjRulsRLaXZVfzVrvTNDer5zibEBHrs/AWheWOM14jb/JwtakhJCdxugPx/n+C9QXheo8vp1Uraw
FOl6yMM0SyFxh3CVH3SCjhlldEJ0PQJ9/f751WHPpOSdOqsVZGTuxvZ5sh3Ck7xUPN6YRoSP97ly
P1DYKdoON728oOCBWMoBU1ORZhOpR91bi1LCHOTEgzzrglif7qje/Kn0a49y4RfVXQ56YgHXFPaG
cCCwwTvKlE/Ho2lQ3+1fyJwOPnccgQokrcfCeM6IOWyTKsfFlbT/Gx55zSAvtGwddIdWsrctE7nS
iXHqQJlzjRA/asAMaXKz2u5pl2mgiZHBWxnrpJhVNO8KkArY6CNpNeA5MLZF1CaJHrZqZkruRqxr
VnDc8x+XugxRS9a3oX1Qm+HHvUCagE7pHh2hwbk0wLXDqTiEb7nQ9AOugAaS9YX0e5yx1JH3afIb
jnnPneOk2KHuzD6m1S1yFwL1v/rvVfvC0KUOwcZzMUYRUcleRwi6kRJl/RoCE58+G0u4F+cekpbB
cF7XrzxGDl0Fta/SSo5Am7Skp4Jk+4UVEPiCvjm9frBz6U8Y11FDnXrej8uSpKOYzIaMcxbUyxnu
OYAzmVOQs7L5B1gQbWt2Pw1u2gnA3lBKmIi2wpT7n1Mo+4KH0ShTQ7ls+zbKdt+HvxoF3kIrlrfh
9Ln3jpD8o+Aa6VgcwiwOtA1K95rWYhyX771I/33fc1i96VIJyAMW8DmUsgn96fLrrqwJHzhFf9Ar
FbDZia2+UamoyDefX/qXugOXsm6XaLAuucWWNvAOHzWEWV+UqdzPM9COvRhB65M2RI5+TQt6eu3z
ZUTMsOkPImekzesnl9Sa5DFixrws/UwoGfszBHNlXhL9GXVhsNgiFhredKQhts6G/wJfp4oUy6Rc
USW04S7DMi9fLFId8kfo+KKfsSNFGvDvF+ngaB2rsCaHJW4SJl0TyAW5G7gCw9SHnoXcP2utndYW
FPUpUbSIVV2ILKkerJ0fSAL5U6K1kZBt0EqD4rf++j0O3Z56e/I5mZQ81pKqJPKd3jJEvRaI7wpw
5Nsd1XDgxshEcJSWiAafAwLOhE/fh8fwXMyWveWFNrAxb0IvtoMOLZgUpd3Jg60M0FLfuaTkbH8K
RZbqT+qA+XqIc5ip4vw4vXuEZcYPdrP4VAC+tmL7YaaQCbeP86EK0Bamw9mqwAJ0mFgduWxKlEYQ
qeUQcW5d05RVzlFnEmOmrnsvYTMkxefyYYL0eG0M+neYgybklbTRIx+wZnMXXXEBs+28G1gLKLP2
SxqR531CsibfJpChmgLmJEgEuwCJwidT5XQ/vMMqu7hOIdMQqe45XzsYx9dUFAEZxketJZb0vU2q
o48FZajrNzpXvrFtmeHvGgIwmdAzSMU4212UtvQruymlH7dnb66t8SIuDDJsD9/tMIWm1Y8jYsWR
5OJesfadTSQwMvbOxo9FX85Wyw3ia7knaP+ooLAFyqmqSSMpJ6MI7fOmdzJfFEyGU/5RzA6t+AIY
BN2j2zlAy7OaSfoxytKYpUpg0ZaNmxD61KndR3XNXcRybGae+dSG2Os5suItptKWk+GtCgczXbKn
DF1pUwmOldJY+TQYadf1H0XfGRRXV8Xt0r3Cb8zsNauKqrLZafsdUWPXaX5ck9BexVdolNmtLP27
dEiW2MyqFxT519M/hH1xLCw6hHDeztEhZPC8faV05IJLd2x8Cv3WkMAqyZ26Qf9WoVtnKjg9ztr9
w6dzI1yBcjelvLRNkegAITfvJLZrMyjHmeY/w6SorAT/6OXS4IKdfNq677UOCMC+rxKMTnSjxIrV
dr+Ho2IizVVybgn8yIdIrk9ta/vqIDycdwD89G8eNRKSc/OSeuC6rmebXEhPY+TvBN658T5bUM2N
7Kd+UX7TVW0GXlUXlCPhJ3rl8hGzWBk8tkcx1TrUjV550DlWVWku0eq6+dzsgSo3/7CnDeQDuHgQ
8OhVZ7qLG6n5AkBLBEItZdfKo24MBklr8rcsI38iIDQjKnvWIQfTIVBPKoWk6sdgTg23/ualVzwi
AX+uQJcA7cy7IVmDMXBWn1lCnFYB5jrh1yWitt3txAqzM8aNHjv9ShILtPxUrrQgMnq9I7QJjAGj
EEg4CVGOGEiWxjIKpHDOaVbN/1BJ4eKorrwPz7X7wCCegmjBrZJwxcfvxSXC68mRMgAr7dAoP7Ic
WTLH2MF0bAMhmTXdEDKfKriOauNhxub47oMd823g/Q4L4HZBaJriRTg9prK8WSGxkDaqiGuZfVAg
/B7Fkl99xTKajWrAzdkzgONS5EvL4B3Z6GA/ZF65CjydyA61eciKHs2F+pxjTtR12rH2tHIB5PYj
p8+nnxbLZKhx+P1trwzOOxweseuUnaLFXll//kE/fbDsZmfZEtO6FHFnxXNLCj9Gc8svWfFpZH2D
4ShQg58VZjpfFnr2pH9YDGFI1iWwrDW9AHgfz0ZVqKXonXpqcMn/92W4QVUvefeRVjj2Q6LTxe/I
HnFDhJYVOzde+pT6/W8pHVQsInVygY9PrpeCik5e4Hmw4T6Cem9bNIwaA2QnWdYJnJJIczjLOZGL
h1zBr6la1/i3aUgblAjydDV5ruK4XYPzBxWZByZ+FMjVnzYkATTMdduDn9kocJcxWsjkKpaKCFFd
msUfEFj5Zt2G+eOXQUGS4pKKZJrxmmgfz6zkCpy4sp1J82n90+msbPAauBxOhbJTwsb7OukbCzfN
kYXHzHMG1Vs0bSAQrAVMCTH1uqQKiHlKzrppVT/CHF9EFJQd7VGcz55qmfn/p8c8AR7ZmfGF1+Wg
lqDlAzrh5rAb/WB7xsKnBeIystNKD43OOzbH/zARR6e/A0yUrgKtYmmIMpSJkDMvngzvXcdvCfoE
Edxvwb9rBH11lxv4MJgj/LBa2xBxQOGV7jWwwkADvBxgEbkIhb6xK1ZhlN+7k3QIXrAKc+Q83+IM
xU/GsEewK7GFr7xxK8PgYL5OEvxETGVhqpD33TwCSax40s+zWQXzhZkSIHp1BLMJrqIzSytYDHdJ
DkHXkXeB7BhQdGEyBUOPosYJx+Sc6e+8rXO4He8uTYS41wpxdlyQUq4sW36TF4xgx3zJDpOyccuL
9Du3/+OdQvUDXwv04KtD+Ld28oaG48xJccenW2nYnSYrEWlji7BIL2Rt5sLHP9+W3xmqu0tZr6rF
X0A+sNvNynM0jn5j/r0AUq5RIN7uwwd1x5DmvgXhYXXcxAiP8uzg9u86IE+upUW1yAwblTvX2yFM
yz2uQP+mVIJ3y2iZg3hb5ukQhJ2ICK+ByS8lyx+dPIScO4XuY6lvNn5JqPP9Z5YrGg6iC4dSmWFE
R/zAFLGy/HJ4wSuXpUMmIrBhBA6aNYGyq2temYbKwz+UY8Xwrj01O/zya5xznVTC3L+TBafLOFlA
KVVdycP+Vin3dJ3usLempkYa+PJJeXJ37rmvUIpBejQBddFSL419EFYNaqtAgDbu8mU45HjJJLZd
acr7shXTN4qw5H3T6cRzlrHq/EHUI//AUqGnmiY+GuX+GB1EXF99c2B6wH1d2B+sde1As2RkQHv7
bE/aEDeDckokZehSqfcSHiuFjmMNWCqZftZl1bwGXOrtHBHE2ahirY2VCvtbyFGG9L8+2UHGJ1yf
RpMqXLZTAdwNE8txZcpw0cOIJa4QRkR73gTQJazilvAVQnt9z4hBCmO3p4wtiXDCSwC28klTYRjQ
ZrsZnH8AUKU76xK9zmgJWK7Nb3kitAMnw6VWHnwdCZBqWucXvCnRbQuSA6WDOo9Z0CBj0UpzeX0G
LXBqZ1KSYogxooC9Wf5qk1bCunxFIvkulXIgzbpcDTzsZj2WoPEcRERkg/2+Z730l2VSo/iIQNiW
nc/gwvJRev4o0/iDfYGDSBTOOO1omPqtNfCiZdYjnAgHBZazVtjZ+dz49S9eaaN4E6SuhBavXJhL
V0oOKJlLZssRKWO37ZB3GtiR3t7MN3S4OOwur7pp/X62fRoUOeX6bGlfaW1mjxB1DhS1X65boecf
0uX+gw716nE/6Hjngwj35N7+0bjhbIrPwjfSW6ALI4tKWtp3KxtRUUqRtrkOP33XUym2n5BIwDc9
LLkjA3qXyP5aOW66i8G9PNTZKfqtdzHzhsZMn4J95ypNPhawfdeNQf/ev4XNwLK5niVl2yBBYFb9
KZ/Iow6sR9ENvGfTutlhmo8kLudB2h15yfakBn/OOOUgNaZR5TkcvkeI5kPpXwx86c6Md+ZLE5u0
Eb3QI0r6htEKP7l+OTvN+66B9MvxiENKc7UcdUEBsdst7f1WfdfMIOpno9QRIXdIkVhgDO6dqvkt
3TjWLi1mnT1NqDAAvqjsvvkiH+jgNa9PPcs2y8YsKLp0iVfFNSL0JcEEut4c6dqZVe9oq9sJjUbX
R3OcP1ciThSzSCy5bfDZ0ioGb+bJJwlTQPMSv8ShSCnwjO+NC+4msoCkBBZEhah0JKOz6TCUrLDJ
DCjySAW7gAanbrXwD5X6pVRmaQsvfKuEfrgupjYGHAOmyu+18Eqzx5auNDuIfjjp77TXySXvRHUs
4ROpbTHgM1DPSPOv08wf8KVnXCvw5dZN28XJhV6/d7ZuEvVbDLVJcoYPVZI9d/0mZ9rputTy6Pgj
43AH5mA3WvMZSa4XssUhw17a/mIMR6TXTFzWlqTtnKZq7Aw9cUXXJp4L2z1RZ23PMVjZAy05C3+9
jbugzZIPnIj4Eptct/oeRStnL92gJbSkg6zvdEaUgCD7w/hmdj+AQdJ3ypqFVQQujJfyjXQc58w3
UDUIcOZLGVKqzTu700L+TsyHRKE+zMnWAuGo4U1Fr15AKd1RWv7HJxsUKiX7Kyx499FGG6kONNmS
gWHQeHNcoz+v0die1eblLZTpcWWXu+ScLqQonAZ2jtT5VzMH1oftVv2kb6lsc7Yo2bLpVmhLFMER
P4SRsvSM0fXRI6hscIX7z0hmxYQ93SbPFF16OKccXkWJTFe7tVfe+7WhRAeVPgRgBts5eAUs2PI8
GeZbjSwixtnKqMbzF0ORxYGo40GDLfTMeFZLqemr3YSDvWD5wjVeI7san2spv5ZWRK3n7opoIB06
IIcg4VT8cPaLtVFoFJm+SpyRZI+/CdQsad0FcE33MRt2/Fm6mqFjI4oZZY+cbC/vw59xK604AvUB
MHliXp+ipcjiuOReqb2ZSY8UmdT5vwYTFrcWfayJQ0qA1KGQJOtlpJmDFk+a/EhNuCdoAwKiSzi3
evNxyUZfLftFY5eOfuVfeYdjmqpox/VeaWmIfMQfTHuUUh66IBn76C0QYJHDDbZ6y98XapAn7BiF
OyufYOIwFYvfxH/i/Smm5pmBVUHVtzP5bQaHtCmjbsBl+gk6ZBXLVdIhvjXioq7cJkxjTTfz0l7d
EJXYYarpfOCkQW3k00VUymrqWAN3Pw8j2vC5AAwixx+Z3uQ2yFNFmUfHGq1N/t2xRUhjgMit5bTz
Aff/xjXRkVEU4xEatX58ceh01yEOH0xvzCZ5PJdzNFXOExGE3lf0nhOwZC/1AgkUEFdTEvmdAJFr
zI+xp9Xmq52te488h7nYNvleKEp4/QbJ7OEr1jRovdKUvG2bRBhckEuwvhE19SpN2PbZ/j78Oett
3Mgk6wg+0EDS7oLF74FHluxAEEJAdVmhW//m3iEXYX8fXv68W9AvnSZBe1Ahu8dGwEgbNqEDPscY
ZMWL1gn6N9Vc8t+kDUo6xBSazL5ZADlJDB/6vMtD2h0c7p7OaUvAdDT/XaYcgNp5jCCVQydLlZBm
UPxpPQh38YaOtcx0j6wh8n0CI19Xalz7jGu3UP6DYgfP/Ejf88NgkC09JkEhMbh1nff3HsJmusrD
PVg/MFgkF3jpaINEpaYNzJLjGTNjUWUGiFh3JpaEDDWU/i9K0lm3YVzAQrWxo3FVWUSKsHNM6lDs
8qfZK6AbA4AOlVI2ef9T9J1MfZVfJ8tcyI4RI1dpWocIlH+Or71Bct6NXme5+tfXjtpmnjupa34l
+l5wXse6TY1yM4bSpUlOxRswaCp2i4CabDNE10AEvlztgpuuFdxWGxjs3ZiMpDXFPQSKzMtXGlFC
/sHTZoCLMSnBzXKd98vivFnLkCeXCKjjbFR7+Zmkko5wBXGLulV3NOg4/QdrJS/ftnHcJKX2pPte
BqdfB5spsRQtCsITLIBf92Nrtd5P9M0NqJ+GemymT+sCe6U6/wEAwqc9sQq7kk7yldpGIvIg22+W
bv4hoVo6vkoJ5Y6Lgd9kAxlj439/hkawr4mLCH8DKn/WQrvfuLPYI2OGYy2c2ye9hrpCiQfKbm04
iWwldJNJwV+2GKQ5CwkWwqsQS3Fh4htQuZOEUZzeTfG4aE96yv/HYtEPMIoOsf7aEl5H/9uFoZF5
gdqcRPj833VZIvJGopDdforTZm9mGiw/2bKB7BcxgrGLY676JnPKxiwaUEI9hQ1kY1s6M2NRaeD0
3nvEUKLMRy2P+RxMWIayLZM6GZHGOnIMU0iU6KLqBPquGObEgA4pEDkR8/V16EBT0/Dklb0O2tlA
DWwaDX0PxJSFhH5vm5d1BuVLN9HxzWdRibw//usSaWz6pNBHWJpvS++XW7FTDm992QTw0a06leO4
6Nz11eUdz0hMrLTMDO6caTBOEYtOTUYCXUEgrS9nFSyErwAkp9v0vYJHaaSdtjyVYyggox5t1oYL
zTA5JoDE7ja7Ynna7BjYMNNEBYvEF4CyPgzIYb17jJnmaAPnsUzZrjW0mD2h2bW8z1a8b9Htpqrk
05oOsBP9zNUzYFuaiXqEr7pYkcvKbCRCMEads90CdEvYtzSilnpAR3Y2R8S8O8gEs6L7NEuRjD77
gjEYvkn3Naiuw2irP5aymfSQTzbcpBTt28aa4IEtq47bRvWW1JaaJ3SA3NqOsZiHTJL2PVQ+cO7f
52hFYS9SNbu9bKjtLRzLKgPpG4GiQ/Wor9e5IF1awVfnDHzz+hXIrDUAeNlsM/ApWBJbLPaktvJf
TxtWllJxumZEjfl5/FtFtO1rzqS969fmiStcsz6ydfgWeF2UkLasf5LbGdl/nmjgAO4v1cjWQfCk
nuGfKb8F4QKRPOhoEjoQ8Lz73vday//ZGzyLY8/JEBcLR4pcMVsqPcfV4G3kkP4N1URjwyLnculM
BdYOhr8LvQ4uYk4GLS28gM98etjm0E+DW/B0876yGbO6qH9ore44lAIrd1u3JWgOyCGA6btvAycC
wMHuGpg9Ma83zvGVHuG1piPDUo4FI1kB1apzxEseI+ERIsPDgnQ+Vp59lJKfQ7c4Gw5HxIhvOrtp
cHOG32Vbht7yR8hriUhyzhVO8Dt+zYzbKCxb/2vkKWZmhBFYL2rEm7Pw+ob9+lRkqwEfSl0SJRXQ
0qpK5XvyF+NH2CvFCxuFW2r+o6fbvnb5GYtX2v9nn4y8f9lKE0KZ0COq/DGPCsBwyWyQQdGnmEyT
wIPK4A+EgcnT0eUAnsro6dPyZDEwE0m6HcLs7uZ+I4exH8V7W/xtsfj0KEGBT3Gct4VH/J5byvAy
b8J/tH71n3Y17N3KPr3vLv3xR5vfz2RaxACku9cFQXHxzhg5mHYZIfuFyEecebPBJN2XSKIk4eVE
x7xhn9jBYTCUnRUQR5GlyNx16VWFqAKmOwVvMoNLclWBCs5MspONN2UE5kgWtrI0ZSDsin9iP83G
IzAQBe7r3LUPKeZWp6znPB7NhFtLsUZJJ9qgwhchFTqGyx0D42Eq7biH6R6NTtWQyTMOhr7tidNn
WUrgaal+bbbqv2s1SNDXldFpO83kSk5/A4c2Lsoa9yyLwJ+1XlzdOGkmzsCR99eQh8KK3Fv7lqCt
iDvypX5wqcymoFCycjWvvAwKDG9ZZGlYGxrSE+L1sang5VhNIo6SmnMWSZE2vf7TNS0ZtTpxd1Al
FAFqOqJkyfD/CzM1/EDvikjHULr/a21uqRFl5nMwogrQy7Lwlnyvm2QQBuSUjuefbFBIpXMvAMrW
IADePW14ws6ivxzOCx/wE4YlpTy5YPXDl9oQV6/s3pJR67G+oKoM39Np6oX/4UKCMWGvdlVIT1VG
4SD73C/lQLHx6Kx+OScUBqT56sBi8ImtntcV+O+5vy3HXzK2pY2zyJC1kDPJdMDfwtAGopYBeqjR
Y2zq+g0MA1mdtUx1XU6XrIXhfdpnzJhCtblVEbOsvIQNa3Jth554cIPYuHT3NP/bwiTsJdUcmzwA
82SLrAxudW6dbDRFKxVOg8s4T27n+6UCWaSbWGchdXGuJBGWUGoUPgW26Hf7sYJeSEaPtqaNnf2r
KTMYYKbc0LK8nzmWu0a7mbW8snRVQXGXu5QQki+7HcyOHQtDsTvMtUx7lM3oYHr/YvpEMIp912Ig
D3khbkapbI6VFjOc9H1ItL7QRkBjp8Em56nScbk4snGELa9WxYtJOOs07J1xOJOuAswQKlOqAYS1
l+DOJKRWGv+vs8vluvCKk/ELIZjDL0DBqAe+mtt1xRETe7guufiL2quU4EuRECxQCk5s6qS5qGLQ
fFVu1U08GxccSjvT8/DuuBlEV+Llgf9084YPfCbFqM99ZNY7TOkToXmkb5AImvXfbGUeFNQoWH+4
JuSOH/0zc+535Vzngu1ViUHD7W3UUvBAC4miqxnpEONQIgnRbqE6/QFAZd4jzlgoiDbGO4rergr4
xJE3oDvVsuTXFJAShO8nyuR5zQn0gVXbPA4eq5WaAqK+cvSLis0xyjggarpLsXohIC6dG+eZkMXS
ShFRbU/7+5+TH9T1sKnn54db8BDQxgzyUuT7zDl7QbN+tl/NOS11uAPYlbGA+HgRkt48WdeFwDh2
15u9iIv6noeiMqft5C0AcXDvPRQBsCLCeoNbQUEn1ZQDx9Pg0CwRFwGeHM6sH3872OCRdAdOT48E
dG//gW24YZ6gJTV78E5IoGxMv5ZaKHMh4ARv8CdEGuoWcFf59zxZvk5frn8CKKuodRLJMjTmEI6e
kmDc2iaSaBvOsFbGBesExUQQOnhMSpluimZyNVUa7NTDjxuCHFrxmARtzFu/CB0OBd4Stuu406u0
zc14NwDxCZEYYFF25n4ggYMfVLtUgH6R6L3vWJqNrZZDq/1417Lvn8/zC+56tFsO7kxRnXI9ZP2/
4ELmgfEAfCi+KUHBafhPGFUArTt57pKLKEYP+KZk836yjy5ItvHMb22aXwRY4unggJxxSYqojSRp
wLQ8+16hVQ+2G+RCvzxBJ7gxzkb/x1a01g1iqQvP//SravBI/CIGxPl9VcyO5bjXB3Lj0OawgS0k
i7DgDyLqVW3OTSEUfXfcJLeMsGpThSAQWLfQ5O1PfoVS8pTVp8xxhC25mnQhXyCJfvyqfzflEliQ
1oeAlCmFlVdJSYD2Y4DGmRVusboXGFZI7j98U0K+LW6stWeRGVzIidYw6mpTkOcT5BH4mjDoVCsP
5i5uaTcXYKACPQjpFKjndwbB1dVdmnifNNVh5ifLea6L7aPnu6hA1dCoH04S+nDow3AuHhvR6uCI
u3ovozU4y7wiA/wPXx3Iws5hvOFnacthQXqkQNgUXPw/pFlGvM1fOQmK8n3+e8lnHuIritK4ruaI
Ox/YAcZF0T+VVosIZ5GGhWWfwc5ydCoSn5FhVjHaLDDa5BlMuetDNIj8EMOkxPr7iOehrL2A4OaE
CZBGe3LnytBFKW98PdLG+F4uLw+tDtdm4jsEi+VAumpWWFpb+Q/mFy/iRyqSwlY37RSTFkJZuwLs
s6E7z8YQZ2LLVdYbN3TtGa3v2q9h1dfxAMcvlJNAX/Zsh4mpFARMGGAR9vqRcTjhXtJN/fPIxZRm
gcFeDZB4krpSl7HJSV1q7HnOCkwUQCcquw9adgRsxOHd8YmCxI0EUm4Fpp2jrmV2W2pF4+aTq+pK
tjolAY6F8+Ic0SZSs3RzK+HXHoF78m/XxAUA2vr/Bgt/szU57tffkx62N2mbH/CjpQ7ghwhExgE5
steJHd1s+HbvzvQqfDlSBv2xbLSd+XrJ594JAQbZVdcdYOpDkL+n1gH1YRlGxrukyTjucYsiUs8p
GKnaQfaWOLH4vcsSpchSzmjQk3YqLid0NvQEalTmNVAIGCGTkARxvqf3PAehrVB8qr7stQkFQPEL
1dudVQrYf7zPQyOTQdMT9bJp6M1V+UVSIidKVWMsjcazPsbAJC5mLinnmtMHt3vCyEVe5fOi1f/T
duyw18WwMoJA6O3mK5iWMEdNkwBmutozmCgnmOLThriZeJNAGaWd4mfKeKQAGXeMJJh13Avp5bMo
BoZZEso2odrBKerbnsN6ooAj5/i9qx+7Z4Mdexofjo6aKeHMsXEhxDGlclAr/CCIBByNx15NSe1P
15Xe5Wiyu0pN29ZOJJ2ybqnKf++9wYxSjr9KC0uR77WkNOR2jPTnz8PFt+esju+GeUR8Vi5BaFBq
M4nU8HkJ8OzuywN6CeE3lp2I/8MEUrbx6IZ/75tmpUECJ2RgOWdBVWeVo9Cf2jvKoZ5ILpncPJ9j
gxIBXgSZVtai99tR6Z8cy1hQw92xwejvI6Va3QGXP6pwjzj1LdXym7oYF0j7N7h3hSbWQcIcZtkT
HMfSlOWBO20mWPN2ZcLoz7dQr23e5eGbx9gVNhaWDnPw8za7rWxle7pkLJuE7Hsw7ouzUkZGyHhU
Bl+1NpX7Ts7dOW51emmzYCTK0GeQ9Lnd7uUQa9Icyq9klUQxHzkwj28I7/yisaXUxdpYneOh9xkB
PeyZC13CmH5P5FLl1Of22HA1RAV5pgQ9L+DMZy3IA/q/eVearos3TZx8jhO4rhMMf6ddV+E0Kukn
1qdtjeq5BS8xf3VGpIf88q+3DPIK00/fWR3GRj9LifdXFxg20k1EU9wuJh6Oyaw4UPRJPFqGkDRX
UW0Ui7fDeUjHlxho536gvsR/2T2fLPRTFDxSAmXGFEhMvUSC1za5KVkTMBH2UTlWnmamPcaDixnf
zmDg0hiJ2cjpyPimfVUTpuAhpG0TJmpyKMQW9XKRaum9RehPAixMjH+LWUtUE9nsOVYVbDvczPK9
nZjd6oSakfcFI4/b9ZbiQQOnzVD7t/55YvRHSstbsgHKnftQKKEZTluPD9gCDmv6u9z7Hw3GcyZW
PehthsqfS9lmv+fhd12xsbafdKn5vP1VharTLbuH+Ba2pX/fQP6F7vYZS7Y2xzhELAhD2TnzHSXl
3pRPJqcqgU7A+h9FRe+uSgZjIoi9p5aIrIUM3dtrVB2Ewte+9fOCvDvJjxgxlwKRsqWa5De9eHj7
bqkpjjaxLNCOrGUUmRh3fc07hxFWJ8PAoF3BBiDU6Ulm/wSvsPlmwvu1iNLEswA/Dfp5Xeiir266
BmBGeo+eCkfBLlVw0D+lBDN33FWjecmuwSKR8bE8VLiHoUAHSvLEegkwzxzmV/SIDOWw94+7oVSI
XeWIteQ4Og29IYDWAH9Fto/RnIg+j9OlH/pxhbRanOtY+fmhPjTlSWxZ8Pl6HbcBP7qEhzwrfoSV
xVkbqLuwrYSpnTj8gKBy6jhn1SkfIzspOLcpK3cTxd+PcKYdiZ8yuCqvdpgalS/AN7W4SVU2osv/
sqj4nvhvLRPt/fETcXkFZiSkO5lk9EnCJS/vlrYStnc4dAgtJCZTV6tt6waWYO9ORgSyOxFNXHPS
03F5UcMD5xuCJS09uCVDPTGj9fsqUxRu3lhjN9gv9Q3+FRm8wJ3TkHS4E1/sKjprr5ESwDcpfYMd
fbPc9qGU/qLyX44sbVdQSfzaI5Fbu/+IJoZgd7+/JDtvt7BP99Hex9H1Az2x79rxoK9lhyUt8zzf
akKwShzfZ0r0sNxijB1m4Skd9DgPt3uFeA0NNzrhfNfSHqWAPHvmExigFgn+lQbCp+KTfnkBaeI4
L0QOvTRz1iYl2av8rkaFnTuSr3yajjSrBH/WdtPnWdtLc2f1EaGtTCeNgFmbuJJu1lhKRfxmP1Oa
3dCXaDSbp0qbz334mln7vH59zYGXtqH4NYvMbtnZiz9CQqgrcKDe/KpjF9ZrsUrAD3BwDx61/OG4
hLpXQ5K3dzsLP7AAM4uRmgaAQgrneNR4bLGPssW5FBwAl43TYeM68dd/M+PT3tFr4oA5rDed/L92
/PrL8Mqkx55ldzX3y1vnTxgUGi2vNahr7uc87Eu5+5RSutcg3Sb3tuYnAoY7RdXf3fbItQocNx9F
D0BWIwee0SEJIMguVF+5Rwi1SdAEqofFWWrgPXdFPOyK4/W3Wghjhuq7YbMwGVIJRBcHcqkAcyD7
aThbGwuBOzaTYCCssqGlu9VInNwUMRd6N132NJhPabKiLr+82iAQ+QhHLFu+XVLCv29FUSgMw/Yc
HFEy2riMWFmJrV3o1oUA1rGKxfYWtfmHU66fqNSEid8l/0JPkI+4FQXCsyrop0DlUCLnPkSh/qky
4d2Tm+DrxJ42dT+rX6iy3NfIzF3jawRo3caGC8IoTqFf5PWeFm+Wh3WIHeIa9fvq82kNh6KV4f6x
kk2ggZrmGYYNqMQ6OWgWl8jdsu9SotkHphI8XAz4YNVYOe52dqZVR5dJHfiyD8iKHVIQZ+Th6gsU
f2GJ5O3sKp+TNsfhGUd8LZHaRyp2sFQ9W+er86WBhGSzarj0g7qgrQYbu6r3lUGZBCqqYcqSPq3J
5jCdhUHAKzjZf//wTTUyuH2hcmY7W92nr0zjBRHVdw92icGjWx8Uo0/Z3mNprEHTxr0Lwqnp6hzU
NCAeMqqQAQGUrVbPjGGC62QdeEgc4UiNOoOSOH0CYXNcY6eqOeYR6+Q/DlFPzhLWD4jPKHMWIa7f
+wJsp2Mg769K9TQoFMWzdprJiH/bUA1yfbidosRmI6z/FzT5B/AmDGcK48LLYMSg6PEEFQu4qrNo
9jeW5ROVyKNZnhtJlKN/4ZxbwCUEoytv+v83zzyEq7BS02e6jHTeqQi/6keIBONY+6EN/8DvcSb3
uJV7OzLVusa8WTgVxnj1aP/DUrPJyZAUe8ihv8ysrU8CoEKxdAITT02YhUaNBH3Ic6e4TAZxzP4c
PrXPqwzW3a1GFqGiekB88m7fgGDhjgpZZUH5I7ch++n8OwzvkqxpFAnWw6KaJQq7BHj9iPeV5Kh/
lXDkQWr6qg1/T77sUfdvkuaiEpQAFgRQY47KUpET7K2JbJ1c3YkB0VrRaDubYCRbvphdlitz64Zk
Zmgj3BX2USnwQsryP6GGPH6nzwWuj1kh7te3PHUmT6XSjDYiUg3852eCYBkLksMxC4XIDqZiu00U
Ivb2/0yxHKLV5JOKzHa9ZtEhSDDkhhxqkqAhkbA8OTTGFNNUBrpQSEtAwO5TuLXaT5dLgwaoHxyP
S/mUc9hyxnhezi8b7Ny5XD+t2ZWUMdn2b2uRsDbBjF2rY98xVk/MCb6AKp9O5KhnSvyQo/7GW8Pi
0Tb9P+BOY1e/RyYdNW6oe82bfXAm9hyNV1tHwEEPf9IlDrsRu0STHHRgqr0SqDKzBRMdMVhymGrT
wPowUAHOTl1tKBJZr4epX6Wm/TMZ6acKFAZI54RF3atVNd1SzOVvuhjbo4h65R87Lr850xkBKdmR
PLKqos6CFq0JqZpIFk0rK0dKz/l59x3aDwoN8Muzk2Kj5vQahA++Vnc9t1lOyDH37/q+WhsOSlhA
+anNCZ9TTydaGDfCFjhTW6Q7b023Fg/AEPh07gLvbEfztdhY6y9GM83zXTJeopd3fhywp/8dnBPm
79m4GL+QXeJ3DpWO27+GiZjqpcJpUNK/tWIXjj98WBG+QWr0Blj2xr84wMf7ZFvOUOE9p2U/UrWy
6lzUhxyeXIr0FP+SiamEyw7KtdQTb+I+DsOBa9dHe+BkOHoElSZLJAjmTHs/HixEURPnikWnfSf3
WYhukc3n5Z1gv1PSgONV7miyhDkcjGkem/PL7DwL/2HvPs2piyF4UJ1P8RPYJ21rNrfRJNiGduNh
DnRBeNL36a76CHja8BPMUQ2mXgyFKsZO5hdDoeoaNHh6CQNZbSeYUJKpTwp10/UNxqAuM7BZ/lrr
IRPybVRZ4gPUTQnEAN9uwToCDK5ju+5NOel2J28P5h6Sfv7K0Nd5iPiNURpdWPvIygullyMi5uRX
NcuTyxR57aakXGs/jMWmWRAQoo0s5sTIDr3+OpeDTTeVlURPg4hZqTNn5G03KbxQDIYSP27tPrW5
ALWZyRevrC05QEd0eJ8OHzQvGT9x6keJF5W4pGlwyLGg6OqqQGnV2QiBx+8/F0gpFEmApZY3MOnj
hUkY6i64peFGnW0HjfDg59b6P8g/NhDjGsKaAG6kjBYxkqdB+pt1mq0JHX29oxY1R9l5/7CcE5uc
Vr+ZkmNf17jkunD7uCgZmRClytr3TJ1pLWyMfk1+ITrQ5fv5bgLGYDbPxFA9TGSecmZziOWfRWRf
h7ie/u0L3908ufNNEIS5XGZLiPyX1agGfqFT/25sdNbephJlvbBIZ74cE1S04f6kkInRy9XgE4eB
HErfetuVDPWOJHmdaETSalJ8jHdDfbZkxBDGgzVcfwQj5kwKsRMUQt8Oj5HRywGs1m0OSMHpAPYv
Joz5PUr3OZGXobWiyyhqr5EjkW4jC0D8EBdzxak9Nr5KC2arsbENj7UDQw0Hkqns+pCprrmqlUGs
8+340hb5Hkr4Nq2r0mqf90pNN3d1YRy7OgBm5t02toh8WY8zJIkSLpzTYHLaVBbQCiNRnLrFfjud
l5VOAOUKc0Ec3kpd6RGpybiKioH3Z2THN4l/45pfK2Q9ZDtdYa3/PiPhvFcgqKmw3FqatNfe9V3y
blkH5lVJ7gefkH7cv/8LDkO8+pBSTesMc0/ZAoCtgNnEqpGPNwXysid5+8plHi5vUsNJH2OK3yHV
x6z8LU1vuYAgMn6US3hr2Paq3FANd/Ocw0k54PilKZVnHJRV1RQol2RhX7cqCxP5PatGPy1Xp8We
I2idQ657J2wSBgtvtoTGnkgIQbV8umPJrOfM+NamLmR+xnD0ybWDvX4xTD0rWZhvGUQMFAUtjO3g
WGQ4iLcYKkY0R9KiicI213OpWmUuxAlBs3zmoX1SksLX4Ghn+TCFKyhSgQwCUmN5rWP+fSazcT1B
WbiZ2FKzDWqH9K2DhX9J6AnDLBxdmdwvlUgnRlBM3NYN6HgQLfRLYTrj9sRvl692IPWI9PendxU/
epucJd+mXiYPArjnax1Vt6H54wL1FqykAwYgV17oZjpra874wyy3maI3LRI61IjIJuuZP29acfwY
Gr2BUa1cCcy/Xg4/7Ok3lyYf4x3ywEyEQvPjPo6RF/81j7bMytOaJudeHjR5UgwoDOA9/PUtxV5c
xZ2SZJxViBdDo3/M9iXR9zfy1n5s7S1JPWboKRZpcidMBV3fXKhx8m/E/zlfbS6RloGkPDnZKfty
jVl/hTqn+xHSf776uuJzm28NVr8pcGloEyIVbz0iPnzcyegB5vvrcqQNYnlE7vxJqMbnYDr9QwRY
8Z+7Rdu1rOv0dMdmWG5IQiEQIpkX8+2XINQrFs3b1rs4M9S3vIfVe2I5OZTX8RwQaGx88PFX8iL8
ddQqTK7UEls1jCmSgrBWsobuNkk1Rdk8FEC2fTdYNCgqxee3tZuBanKObY7II0e3hQYkPyMmUYnT
CG48gp5NM7yxfyPeLo0aCy9JucszdJ3nl1W5Mm1k/ywMyo80HM2NCqheJyCJsi8qQUt1wIs47BkD
V14x3wd5gvc7BbN3N9xjmrNYzvihOUuWF7skdlTu0M4r3D9wEeoH2zZgmv8ZGuh/8yOmPD0G9pXj
RDSR9Z5SUZBXNDYrZ8Drartpt1Ml1aQ33GP5ILm4IXaxfE8Ns+2O0awM8WDlLDyIETRz1GUxxuY7
Q+S82sRDOttr+nMbxJ1kO1BlLA5Zjukeb8/Mihsblk8oxztgRCiY7LDOMCDb84ikPuS7J/0LLcks
qsWg6r1mZi7fBSynfAqqlaBIh+O6aHceREeTDV3cPKbOWfdtk9/yCUL9jZupelAesRi5QO2gZjI2
covsZOWQpb7YDqZyzPx9pot7bFzPhVFd6WYOKZq0tkZhO6CwWLVio+o4OVwWBwrMIjJOSQz7EC4w
BirM4oJ70jCauDShoSoMc32jpIhfEeuvc3TMVDwgvQOJjKxpsyeB1DPviNRWgyyeM9nBt8v7cKWW
+Hz4rFMVFc/2aTSh3tqFlcZsSnjrcx4ZPaP9cuKbn9D3BUL83lwulqK31V7xm5AFmqaLVye7Ih+0
kDAjW6LvVnTBnCpk2ZfasLR9SrDELIYgBlti1URVpHlKXwHBappxfEx3g2EvTlT3PW4NHMHM2XXh
rT8ELu9x8D866vsWbYUGMvHF2IpgQJSs729zIX2qinsVvCqEIOe2wnnLR9/2rMspIGQDwXXqulRb
ky0uRIwVgVzt51UXrETqGME9pw1/hVdjFyxsWQWzvh9xOCZkCxVTw8DXHnpFRzctjuDwVZfYxu+3
rBIcbiun0OrIMOFDJXXv9+mEO5Oj/M7TlY+2BaanncuVq9FYj65hBQmKMjxQMgsV7IXFU+Vx14aV
W4gv5Zu62/uBa7R3rlrlDyuvkMneEi5Z+svL6NAtrDpJVut42MmCUfaD+YLF+zEVEuiQjNHKZxnj
mU9rX9LW/sKL1zdr6VCouSVncAx99iCL3DfDGRlS/7s7P/JvTU5wG8o770vgpMF/b1WnqCKNhNCH
gOxxhF4+UU4vRXx4ivVzLx6Xgd2Nij4O7qW/jd8gi9dj5eJ/79mfFZlAWRvy0JJ6/7ZEd1x4CkJ/
EhckjThHRMJJaGaPJZ+4x06x1qWho62AfX0+Z6TqHXXjQ4VM8wWKC+4Kxlv6aCCjHgY8GYiDTfiM
TOqBMLn1B7JaMsoVYPjoOXs8QhY6TVSuzOqjWZvE7TR1gCT8mAHUCxla8sh5o2eXMu+Fiwab1abJ
gH0S/jxod6NlPrOHk7Sz5KaXiZgILZbcsFW+6Z+LLuLiFRFQiN2Gih043x1nl9IlnA30By7Nu3GM
U5K8dm6+GGy0HMSaaLOpdrxPkX1NgTlbUOHZ6dGM747OAilatcUxU2lUv8dZ8B36k4JP3DK4rtRi
mPMw1EgpkRYEZjUb1C4j1WRfRYVdgYH0WaHdrhLS53SOC+61fJqpqJRJTiSdRglHdT6qQShNhaXn
vF6RnUCKlH+Mp526FReFrWMR1bBi7fVTv+Gcc68WMqtqVWQFt7IKVRYC+Qx2I+UGsfpBoR0jLnq7
5TZJzejTTz5Sm1c/X61BYTN753hU0LWTmaQNPLu2LsaqzgSsxvn1amQwuQMrzL1anQWDaUI4ZqB1
BGd93+fdPyVgc4iRf21L4XXJ0Qj7mvPzGl9Veki8tor/1i033f/7qyCKwG6wy8h6YcMkptfPLvnB
++dxu0NA1gMP8PB8Xj2kJ14yeHDVS0KHHBDGU4sYtXOALINtqJel1vQWg2bLqAKQiDlqmRPl+IYw
IAxritzEcqcRhwtOIgeS9fkBWQNajxMUnyrAg87WyTHW9TMDtllE14hdT86UIFwn+W6so0wsKaKM
Z2hJAnmq81tcOXCThtDcpdFvaxaL9OMDvGonyCqJuirHgmQidbsH7m+E1zQZGjffPtnPOu1jy9Mc
KJXwY0Lm9fPNdj83zyKb/BpkYtZn63aWdqiKKmPIfBuiq/boCNHWbyf3tJVdktEb6FdseCPl/vNX
yR5N+B+nBA4SvjJ7SAsfW44CUbqSicxy2WQKp1Dr9spjtW52R1gc4xnUsF7KkCnK+/UBZj7B6uFo
B6sTYCkKWhifLEEzfK9UW/ttS72VYQFL7188dU9u55FPTYnALsIpjyWoCeAaW3ZcoQcwld2cA4hg
uJ4LCmIO9wNnJKEOn+EHrJRjLm/BOd2Cq7BFLIPY3HFWVMThKrblmxFq+AJcM2N1MlJIXpCSUC9w
4DxK+GRVsSTHHo3RYKPgJqxWCFFwM3cMnUcm2FKLLRfBFNoYG7o8zi6wpTiE0V+7J33rcwyCkZXn
Uq/kW0jhGvJqT/6DiYy5vr+iPfUY0tvuZ8TT0NjCa0J+hF8hb5M42b060VOcWAptYRwl6QEhZsSB
1993UXtQmzEnFv4MACIUO3AAN9CCgA8uF6YIeZwnxEDGKlt5ve4tTlG5MnZpHePLl2rnOU1ThTUV
aqjvOsvhmDhVuc9OJMosSDRWKtPrvH8Ohx91yHRh+WkJWnKKd5qEpBeRYMHlyJGCIpzD+hMX5f4r
49zYsMaoudoA1tHBXTcbezH6oNwhdNeOcz5OA0+5JtJKso8hIYSy+hcos96z0R600hTjH27iCA0A
iUq+Gj+0vnReDNdITpU6ZII0CLT0oaWt4p8DJZdrARgDb40+BxIu6ZIrfAfmGhcDvfTnixPWtCco
z8zo9bWXoW2fSICkb4goUait4wnAXjTiFhH05PMxmrdgaw32BK7W2H4ktQcktQyTtXqM3KRQU/PG
fzYjF6b/xN06JKhVt80IaevCeL0Ej469OHVhIHE/ToOuHyZFamys5XW6ZHuoXHuS4kyeGoPFKDmu
Z8e8wuIKXUYr704ec7GBBQmcFaSB5YLXbOcuMBzmj3lPqOLwkxp2KD7hOOhJao5NHaimgKAyQQ0X
e5ipyjDHft6ya3mLMH3Vd3PbBo3AjVs0orQPzQ4rGWQcq4iwGlHcvX1IFGG9nvRpCcQQjXWwpXUi
QbilG1/dVUdEQkkNZ4nH3/QvwDgsgXOs4/46kiPAHSrZDzE27AvIXZmvRIRXxiFvgjSA6D97/tLS
OBQVXiDfVlSc4FptC5/PnOqGqnVaq+y4eenNJeB11H9qOSKaEP7qwFTLY7MnjHN1B6m+oP9w5esg
RWyDsZMcpVVNVcJg0NJtKoX0bSOuw4qqgz13IRSDDqx/v+3AV5TzeDBS0XKie2/RRGtqJmFpyqbo
/8jlCb0yZQV5fTVmrwvtXHSihgod9lDPFJLgmzb7g3nFM34FpWOu1mTXJyf9AwcAjs8G3Fj5d+IL
9Vj0Rw4q9A3GRA6MTkwIhOhIIoWcQ9j09a6Vba4KA4sNeNQybqQT3WwzQmqvRSideCc52TabOtDu
Du3WG5aU8MmR6TWjDqvRrUf03rxXNgnDsvm4k9W9KF7TgO8MaEH9vW6LpQ6SKENSM5ALddCKhgJf
LVm0sNrHPZy1+GrucHcS9t2k2pTh1vkI+ZaoMfXLkdcCGrQJqcpi/YxXwPYV2slk87lBZ2tJctxM
WcJB+g6wgMjK4yc0reRYDa93UkmonR7u6iIyEb32sW8gPoI6dPDyYwKhpitpRUyxXEBHbGsM+OOK
fi/InGGuIbLJYRT7lwbgNRf4uflcnTg8gPrmCxh0S9tgX6jjPNwe9PVLG55stLUdhlXPMwWIpRvH
enEjd5MFq3/RRUNHno9mYUVqRz7HPTZ96vSm+L/TyKKm/noMfIJB9Ff5vwxTp8mbiPjbOHL9iyRE
isulzrWSURH41gzavGQIjT/MoT9CBGuLxCJ+7WtEmby+hvWt0/zlD4bmlDo77rJiHLWM9DNE7lf0
5MITD6mxrw66O8pZdDhv3GZHlF8+OsZtXwRf/dyGWirbV/LC9ROHDZusn+I6X6U+N6Drf5JfFj6W
6qx/Yd9T5pi/3pk2ZTY8VnSVqKj/TGkuADA1HhhH8JTTrlE2u2eGOlLAdt96T2PX5n0YIknDH5Xt
azf9eqKTdD7/nEs7T458wavaaOf+fhMZkLwTwCZTH3pz+Yci0y4+M9fzEtI6yo4wT98SedTkreNT
M23phyaLzpWIxBqFZsvNUWhoq6N7Zbz6pGotFrnNVpTlHsDrMQ3hr6VeMNZRIFBt0InKwCm7hytv
C6du+SlyOUTp2jVueeuk5CRJP/wYzhEQubSe9HA1OdCVRDay4M1bc5k1hpYzN6jBnuI6L8nw3kxx
b067m4jwOeXs0mxzQ1PNaL3h1sTFaGUEmJKiOQqJZjgKB+F17Aeo/V0vt00imv5WTUG+tHWTsyI8
io/OyJKccP8td++eLHMp4I+ky/F3opfe17hGoO/y3qfEd8YhbK6V6dtyNFkHsMSs+5Bl/t/WW9+E
cjiOKB05PcQ5ix8iuuwHFgyrpO9NigazH05CfzzamReH1pcOv4BoKKILhPSJUViqnSiEq2kS5/EM
qQm2rUQZtvF0CbrpYU2ITCYMWKUPwkpFnGbSXaH+JldZxK9oG2kl7r7g1ndPAUOw15NW/0lZtU0k
ndzVJfTbBP1KtUXD4wcok+r4s3e19T3dAauGqbW9srwPurqZ2fJDuz/k/sewwgxWQrV7ABrL/Yib
0j7D4yEyPOagFpCPzmYYlYtaRcusU4SeqaBbIalvG1DMCHJuhIAGsa5FMLaHsw8/mbozIUrndN2U
H3H5CsNbIz8keycFhwKGjRVGPKmqupLKCWNwZTEpTahPE9xRqgbDug8J5lA9U1gnkl3wTLsCyzGu
A1hgHHJVhPsn14UvjwDcfwJ7ETJeQYzhkYsQrM+6TUb2TpCfwL7/N9stc7O8kqeTglmYrcaNUbC1
Oj29pVaD3CxXoF7xeLKvpuWZcLfzS38jHGKTWi8VAw2u5LohmJWBADDWWJHSG+gMqQDu54an4PyL
knfgSTQBG8T9y6C+ZeyrYGf0IzA8q6YjFjRCLt6LDHG1CQvXcMvAz2xcQ1GaozP2PBPbElXP254R
jnw4hNlUdZA6DwXO/2YJ1OUV3FKeVpIxIZf7YxbscM/dpZBSoCKlgQbdByjEBfzB+OuoSyEGPxqk
XPjDjerEmiYo7NFPHKoBxy2YUNMS8f6EpnToWsdvSygh1E435D+CT/7sYcONZUs+JEwMw/Ip4q1+
TGV/GpGCUh61jxbKrGBvjsN90sA2zPgrkm/HvbAD2sunItGICU/NCOwM8DX7cD86URvja2wMs9MK
1mHEqmDfyKQtA1+XpqrvU1f7b7heWSw2Yxn6Lf89Myq4m/jZXqmjMGrQDtoNarLXNEkqLkMuL6pu
ZOUTzUqIfQSa8sdh+YqgbMATTdFOiMQcp8p2dpcLMk5fKtSmnKliSQNC0yBgQ1lYQa1AQvaIUicN
aa/6YLUPBPpEmHxviTbf3ZQKs1LK/wcxwVLnPIGjtkbUHsYAHyUkBWFZEFPH/yOJqi77dLFJJbEH
RQaruhRht92wRs3mjumKfghNi+lDpVxMBhTcB9vzmDV4vsKEu7/CmbIL7oOO0ydxf6gI45QSsDag
Hi4CEzRtDqzZovzQk/ou9vZSLnC5+yVr9DsQCKlSabd6ONG4xsd/L6ruNlKvEglS7GZ9omsfD0t3
ovsvMs6DyMt4Zb0EMi0hm1ysmN4zuny092sxeNoDZ4JuO+CSfp3FgWaOf7Yj5STY3tCSWnDlR+mu
oXibOrFzdDtQhXzETKflTWAWOdg/+L2xOm7y0XoqpQ4EiYBUtCQYqBXZttLZZiNNsvYNpAOQVD0m
57YHO6wZD6c07zpw8doTwMy+uMg4pStAePHJilvKlXMJjlSQTdRDBY8jmTCoODz/+J1r1dIQHrpb
mOn/0uKhAoryQPRwPpsEYKPucKv+PkyUoTDCPAuWMF8LnOZqgkLLaozY0XWt+CApHUkehVyXnwrS
SM8kX1TjZhnluqcEKfKUp4Eh+w1ECSctDR/pogRird0CtNn/Q3HATdShSSDfBGbqjRpKlc03AGNk
N7KNu3rBxgHBt0Lrj3FQ/T4sEMtaTPg74LL13k7kga1I4UfdfyHha8T/VpKN4C/NeS6hba9ci4cB
k1oge7KVir2rF9Sq8LIpABMxmR7aLQIp1scVlSwEEm5LmdECFaAZWwfFjhazi1RcSs9bVIkJb+CO
tala+tiB31CiazHVWTO8ilhXfUl9AA4+s2ZSA2WYtGxR8xQ7+hV/cFuaCy34JGgjVoqrDGdRPHt1
/PTaw6b3mHo25ep7Uze/DgcRHV3WD/jr+jTBVXO+Bd0mLmXW7sAaAhEOb2E8wB01JYn3mCazZnAe
IAO2Uzp3xSP/8MmmV8pOH7YfSWzRQquTopmJMuljBRLElROQMdfJtovs4spD0aqPSMeH23XODaHC
HE+2GLUjgfNl2k6SYULEFcP5+7LSAROgQ0BLtxRHoxvx7PROEgKaBE0fwZIzrt4jVPr0cKVjEfYv
ApIvLQZ6kpayZjdikRrR/sBqRfYB9c/KHG2haC4UROvcpdrKOE3PlcQNhtJsM2o2rQf1LOX6xGVV
/i7dj3ZW312pnv011v65jnZoRnDfkSPhGNcdiMC1XV0j1VgOLd2Scc9LXtMFpix6r2jXW5irrRqy
ssKcToTVLrKXhSrlX5qHPbjjOWIIkPi40xFUSQALwPIDqxsiHCcIPrOA2pC+9fw+guixpHmfavn8
3Jc/cH9hE5+UcP+Ix4AgcyNiiVs+J9t1zhgHX4KfLyUqCU6aZWBaTxB9XTvyp0m19IF+AMuojfLS
/hDTmHvbEJ3zxSw4tj4WSeTeBWWw7Xmsb9WPKct/s2peXmAq/vv+j19W61oxLUVmH5WBOtNQg6HF
wdPgsxhbkZniyPoHdUklQ8yRt2kzMZ2V7mk9U4V4SuG3hTZ9ZZOfGiXZcA/Svfw2KAQBgsIlm9lA
Q1d2JoJkNbKo22LL25s0b6l7b59g/gZjfaPjGDG5hxICeinS/cMQn7Qs/Ly0ZDkVGqZd+l4PMtj0
cjZK+Zq2XDJFnjV02vj1GM9emcBUASnKwpVpgNv3AsF6uuRuX7me55kxtGcOC9Dl6TZwWywh4hnD
MbiBtpZyNY5pVssP2rjA2D6REeaI+dduOfRoKLy/sl58tWi58RulAS2gTVQBBrSjPvezfjlHF3wo
ksDDoHlHH28kmNfgLlhc2NY0mazcwcIcy/wVjv8rVQm5vacisbykXETzY6Bh8AFpNFx1HyoilcVU
ZOnEKA4m1nB4a0TMJ3Ftnb9ojGKU/J+7yLpTmG0EzbxJgz5rveJCc7a3nx/xP5v03hrFtpnoESJf
Dqu7UK0/zvNzxVLo/4YuvAtSBXIyTGP+xbnIIMoen3sS3qy8ARBD8gu7n/QcozbJ6bDcZxfJVSMD
IV8n7GdJqTmX4WHoLBQ3dh4BpQsonTAdAxue5B3HSoikUJy2ibKKxIq8KRWyq/r5VyQMfiqezUpx
NL93meTCVkt+ptytBlvD+eYKYSX6RmxZB1o8kBNvTiraW9cQ6HmkX5ciNtaYJnMrdsvU4eQI6tk9
cvqHSz3V3tB8CjDvZ6fyaw3EX53hYAobc79I6SB21TTnk2zjYXXlroMl8qTDctA2f3wwDa/hOYkP
Qav/VMur9A8LMwpL1VZ3dmGw0qThpXYkLFApS3ic/3zyMcp2wkRXm5nXLKU6654ZclCepvF0kWq8
XJX9y9QqB1CdredEedkI4MduGRCs+Gw1Mw2CKcyMmC/VFLX6QITF2BTwGhfRIggIiUL83sYH2V6F
TXdYz8Cvnu7MEjAhpGYhCIYJMzaPphtISD51s7SAKcM30nE24m4weak4Rn9kAlEIA1G1UCiMNGYj
mOMy9JpBAGB1Wq6Qhq8xVsFZPEPeQbMfz2Jec91ngPLOj0RNAFBcXu/3GrS7yRGnQcfPfdB2tOBe
pslf5dZG3LJ+pC8yt3y/uVIR/3yj7Q7bs4RHPUgX7E3i51Us4fUJ1SsvZOl9ZhpcaeQywVcV0eVC
LxQBRRpWJ5/zKR0RAkUGTTD135mUWZg53uewgwwAK4PJHAbhEGadSznLb4jjvygWWxtBPV75n5+G
cb5nxE+nqDIRPOwd6Ggx9L05Pw+D2J0Tu4qP+h9CE7oB4MHuRPvZyJ/WKHz4pHPjQu5IHIZmAbdw
v97hsq4RW+QjRfPA1dakxuPPzXPhhlK/dhwuxSLOYBRJT4KQJMYiOQM/f1fkouJVaJycW2XZ0EGT
Fz8uU3lFjYk+081zofgmyHCxQT2/jDnlNMYeLeZ1S8CnQnxhyHeURCJ31cyBF7wcT8aDeUdnAg3r
4qojZ4tOjmmBNWdGimeBsKhO7/9GoxNji96s8CxtN6wOvN6tmZJA+XkzKxJiTs3NAltFiwByksz9
zSC6CXZxYkxpbkvKKWKiqdg+Ezyn2slf51LaG04fJnB3Y5Do3xXmH1mae9M06t9xywj3rdnZ/y9G
MQmFsBsO+FoAHEhYIDeoDhwmcMFnU4ZgI5ztTQnlUA+069z5BbLyFWc8kwvTjX18cquSUqSX3E8X
BIgau4a6nwpNuHMIS+59X1u/Z1nnECX6U3eCvfbE0SI1lXuqR1F3dLL0uHvIrFNqa+wmykXs06p0
UnX28V2NWBbx8h49qXmj8PgUZrztk3z9K0PQDO8dfSkJNeNeIeDJJVaAgzDEjpAgbFwnQCrxmMXr
tyCytWzdlqczbaZ2VmGgFPHl8DczTfZwfFaxGO1fback6I3FnXRMMyfS8XK0dWm2fIm8Pt7KA52A
Jx0JZCMcRLTkcVeo1eHGVPjs/nkGqfgRcuFmo5IZJ3A1BMkXdGdZO18vieQjI8sX+UT3JEMePJYa
d3v8F1DC+sJbn2IAHifso/cPml/DyAP06nJ5zFGo+qtJNrVnldw+6FDTTMbumzw/audPdHtF2uq9
VFYPJ0i6/qo9Yp0RZ81J/x4k94AE/ktUXOB7SiOu2KYD9qmgn5SZMAEG2XHBiwmOY7yzyzONwftU
B/e7iSUwE8kY4t7zelhvGhkJ2wZ0gF2NPdhrzfnCVCjIyWNA7/uoR+ILK7yEtSITQERMdGXpGTZN
13uUPxxl1m1UEJZsx8xtasillVJ0drSIaEoXS91qt6ei54nQbcpWsBJlQvMmQBbPuJJ4Qa7WRUfP
k9gMkhS36KXWUkf95aUKPSJbQw7jOgtfrvssqnQgzatACm77Q9HxPFn+zakpwGUWWzA/+wUYV+9A
s/TGPk8S8oqXiWHool+FThKhQEImax6llwY3bxyUuU6l8in2i0gOrF01uKmHT0DWsZXXdm37UM78
vpo8iqmJ8iyhdOm02L7CvmrVqMS/lYE1VCbZkFvDmEOsporvtAkZPfFNYDaIbANe1D0GmVYlfmO8
UrNz3jrUkX3wx66g/hD+1izRDJCSUkg8IcF+7mlrJJ0gqP6s/6K9Z/efmg9uzYjhAXy8/A0ZTYml
2uIRB3Mh4ilzJAsnC6V4jmKN1q2PQ9REkEa0KpwE5aEVDDImNT32TSIhdHkJS3ngI0MTgOjJ43jH
SvC1RA87bOpoPRJnoIV7DJbCUaHy9416/Ao5aTsnUNblW/GmTUeQmN6S4StMz9TfQUGxdZdxGf+n
5OyhfuXFgbiwGk84H4oTlDDlATuGqAsSUBiJcczjgJd3scrwkLTNPPMUMgOxkRqWGnyJThgXBoW7
7y5Gi1NTw0TIsh9UVUDuk4kL6DaRoWpuFmZDsKOJ01ScQiBY1v9fvptUsgyjYEjI69Tc1Ak/L+9M
/sYaYhE9F9jRdlxIUFFu6/uBLd3yu6jy/195FdHMt3PpFLhpYeb355IWKG25rqa7/Sp3ai47GZs5
/gdRl47LdU2fVU6xa8ai00dlFs4woy1O+AcqF2Pbu0I20XjLAaqt8/AVV5ggyr5s9qnWZnFytgXj
q2WwFZQyaFjTmZwYykQ/wz6kTydjmTMhVJK/+bwSlqMbz6ks/Gwg4zT6yxZjLbpNZkZvFD2A99v4
ourT/TqxC7Kplb6kW5PvF153inUEZ4FZePv9rwyBVY3YBvkNap4PUppHClnwRwbO/Z0kpv1aeu5U
CMEa1+dkpVZLSqbCyag1Y8KSmkHCbyTNn5eB5/inss3RvE5dZWOSQVjwrvH+4QvXjjMjOS37bx9r
t7MB1pEQTOZ9bEPD6mT9YKzeckCligvOS/eF7MaYQzyN0aro6dJ50sZsDFj8DND950rV/rM0dcc1
WjUE7438QRxOvKiHyHRFgwFAW0YEqR9ywy2Ahlr9STmzONK2wZoqGNgVwgnM5ey1+oPh9B3uAJ3E
8lRJSZuqj+6Kh72MTffAKOKe1d8tm1BSZjaMD1gi7p50BPU2jRFVZToApDRswtVTaXHmFXqt908Z
xN/jV16xtYKut/pj1qhfVlZwY/qzhYkGNW89dC5wqGa4WsGdf1d4uRvu8IspQp+ERf3Ac8QiMUfs
w7Ty9NtaGE7We6tMypct/ysHZDeuGW5/WOgiR4V1k6p5MaQ/OfAH1SrYSfVk1rpnAbNPceqLsdi2
n16ABTjbo9kuM8HNYWyPCa06lpCuUc0KXhyUFtbs5jE8itt3g9mf3QAMlAyCTXCGkoy8evOaIo3Y
cId4vDDcP2DSkSZy9T5wSacB3mGNVFFvGX0++a5JgIS4WKQzzv7vca87c7xTntQRGQhRlCMpU2p3
moXmzOgXEBl+hh9nlH9TEx+d8aHpbWmTUsbkbwAL6XAFLwXCaAyxEZXNL4D60Dy6Q+EvWRfgd0WM
+c/+HrN5bhqP6tKuxpYBBSzsFxZyMgmZrflJOajCyLNTt82NhSD+DIy0q8kNayzakkJHuLtIqnDn
GwRMWY5wmc/vpYdE3Scd76DQomsK4XMhqU9JDkQDJ6wANXe6nXunxtCiR/9DF5wA8Egchmx9shar
y6F3dUru7EYsSoF8S4kq6lBeuk0IRH9vWP9h/FkJMsU86iT7UjeGBBdQROlzkjhTsvXS3NT+D6WM
E9xzKhFuj2G3oDQleZtZWI36WkS0RhwDJeLG/LnTsk96HvRv2CWsHfDR4I1y1cDzHo+NRCcuyNu3
4vNd9lTFC6ECchHahO9e2YA9HEbBIrYRJWhfw/CuRgOn0yySSvfxzXtLjaVViAfDWj+jvquNVLIE
M4bXT3FBK8/mMM2M6wvJp7jrdncaevR7XSbXYTmdqCvuabtv3gs/fYSw1Q1yXHskL2HNI97SjNzL
tAm0Hx7gb+tT30X7a3sMtnj7ok3uavR/SVNDos8L9TU0WS7Qj44hoycZaRoPxjCTrtyvvTYMYH4h
4kiPhfHxW9Lx0GLmLnmDrbyiY+RyJtZGb8fsitPMO8+H7IuW+BCA/E6FW0pdwzoMyLa6Nlc09V1g
Rm3WPxH/UY95l3y3skn7KrOyovCyS+MW1XaSvIBDGVNWd6UyA5FrQX95ExM+qSGsLnuz99Xyc9Nc
ggSjJVbVXjkvAkNgZ2pUJDdjxc+K1wq2k07LAwo3/9XGwDU9rctJqn1danIMumoiWPQOQe273Toc
XeyF7d+i/CA425ffzXdw7rcmcmw9QgHxlKUidounQbKzkINJIsmCRXw89Z16Q81IvTrcovgYySAp
vJhc7XsnQlUQquPFucj3FFtAIgetLjtejzCq9jh0vi4nw05L8tvHgmzPN7+pJhuFXtuwNs02ar+b
KsNXBRDAlNR93E3LzMYtnfC1sINf4x+ph6SCvXql/9Q2Rk8tjuYRgd/rWxBewvGRTJ3wmvv6w4tz
5baLFNkBU3pNcBwqg+9s6/w9Q/i/pqcD8aYiJiYGHFaGNI9G7uiUyyb6QFXDxGobLJ0o/L1z59mC
y8qGMksz9p+XIgokd4kuQTfs0+7k9m5pCO3fHRfeEAdzg7STaIp5tKxZzGwLlFV+WoYIfCnRGFsv
4CJhhZrwyh3ULMrZE3rgazKAFizTbBTpMnjQPc9TrN2lOj5GtGl6O4e51oZs58sq1pSW9B9jx+i6
1kHSx6Fr3uqUxpmjexXW0QJ0NTWOVVzS7NOtwx8qcPx7/0rgT7UlioadH6UP7EyAywos1DVEzMbo
8Y2OYDEpkKjO4ILPoaO3KpqDZVV9rDCq54q5aIEUHqZOp0tP+4EhTqefMXUJbU5KdfWTR6B48FHg
CBhhWqb884fJHfIlnMZ+vjLTtoVCG4MToVaNoNZTILIXofOWFdjuwMTTlZ74+0aDoaStS3w5RcAl
Xx14dae4l/Q7YIL63RH00dkyi6tidwMa0b2pPBxJYlFpShjBDW6Yc+Yknt1+WIISznWIzWFTdXkY
caZ9Nf7+heuO5+ptfKJ4mvHwSNKA6vDl8LP0GycspDXGJMg78lEGpIXv/kAgMBXoCaHqNI8XdPDc
+zuECwkAmoKsVPpNkdzhdkb/6UCLKty0gexZW70FsnAF5Qhf0YPOLyttLTjG0Cchj0ReLpP/kk3l
BTZjH31kOuxmfkVWyc0SgifF5nRA7SS9NCWgNPPukTsCyWFrdh3+MoyVdTMyMDBie5cbbyislBCC
ckUB4CLO4CYQHkcDAf+rT4YymgXzyB2W4btzJ7apDqwR4nEdhmqArycnZA1hkV7aCQkIyzHTJY6X
9SaWsJygDU4JJVKpKD268KQQFA/hjC/R5+GPrli7ZezVUMc0zMv5uiST8gbb2UY3gup+SXUq8gea
2PFcxaHdvFHRBGR5aMY5cXB3kuULsUIV647aYoTNgSBS9yMfpuM46MhRF4xOixPa6mvZCWnlrziz
bSUr/Qwc50as+gpQPEZN1ASHYBcmoNF6a5ykrlARBuh/+Iar6lJbom1wSrfy9hbuQzZJGjKfZwxv
GDX355ZErQvn/o/T897kuU3S/0Gd4CbL0yfTZtusRJz//C85+q/hnNBdbNtIVsV6xrGpknJeF4iv
2oaJIDCp2VchNZ2/GwpYl23McxPi/HypXI29YqydF0OOiQNBebMYJ0dPFREb3m1cQbQnFUM1Hvlf
qxMes/Yt2VA3W2J0rBX6YXij+Mkjq31Xs6hm/BXZa8wETpoYkIqmZg6eWMl/fX1tCGAKq8YkdK26
NB5AZNmoB1+jWvtyqtuDm7H1veh8zFf7lJkBwfiU7/d7/crz60ncPnC0FrCsamyb9igkPw7Pj/O/
KO0ANizG4WBACeb0+djFKgXYjFS9gs6jXAj5lKqmEW9N50y5Whw4jEEspFgAsAXOjhwOFbu5Z0Oa
WMfnBi7OYAPT+WuVuUWdHWteIugT18bOOKXpJIAYqaNgUglE49HSS5asZDsLKGOtXiMFWR4ErIbk
/yW5wFyd3mPyMeJCVxIfQgCKRj3iwxKnZTm3ALwmk2Rtp1KFHTBCuZIlF+OtH8TvROKjAgb4qwhE
X6BCXsNQ+UmCtFHee+L3k4U3ry2HnU+zJCw71qXs8pYQB+py7pmR7qVdPdorfopiWj4P+0K2TbPo
t/HTKO9J7j0wy3jsBzRGuchwEx3HdqXR6XNGmr0bgQUY4ILPYlAv8vIzVt0500MBPp1uVO/MXIIn
j1WK2+E1oCwdvqJG6o3PPsJvuwlwdWKr1zoGhJTjgZqUeI6G3v5qZup+IzGxEEiCG8vXnvM9Z94O
dAbYFiPezquV9OEtqeDyQvK9meqUknKMw2gA7YDBqGSF3nhNc0+JJ1GcHqj2TNnqk3wvP+Osxqbw
knAkXmJn/TY7e1GE+1TWcCYUaN/OQCNKcWZJuCS8HDXZtSnnLcvQ7rRwq3UGpvrogKcVWFfotio4
sARZBZ/g30pgTZQUAYa8TRzVVmQaZrdxM53O8fDi3XBI5kSF9jNA2ntYplXrYMcPRMDjy/goi244
E2uNxqyDzAcfMFRd0xQZ+re7kzB8KF/gPkyPrDVzvf90HdVMVflVXlhE+bG0YmcrzDcLs6mr2MCn
jzwyWOKmjC8Z3A8IZ58+qIPqX5PKgoqxfHBqCYZUIgFONp72PyLjkyDE5auoJKdKNCbhXYjpQbgC
OIMHUEDe/RWL7L4TBtWGt9vMIUafxZzTNYAIhhDL2cjb/EB/c15wKACXLX7UlnSVZVz7ErGWRYKX
QC4wGLcyH+3373dFyhJW1UGtIBZ7zADspclrcHzglOvRpcpiJgRz1RUrj/HWSJb5ujXJ8Te+LwfE
QSGRSLt/gjGzreZBw0Fd7dWRAprtucBKYEbS0B84VZf9DC0U+prBknUCj2DMgv+aYbf6t3hmB6Z8
vaH4+egAjU02JXVkZWuS7Awo/cnI/DvtLQlUUJZTiCuW36UNkne7FeZjdW5e+QeWI2RrN2dpbTgl
vlJ/zFwOztR4lNG/O0Y6mM647C2GRHdo43cR7nTzcK7pXLsrTFdAm4XgxirAyuCcZw4ynDVq5Eey
t0vmS8n3//d5vyivOAOtexOjebcTwlttp07dR2tazbd2TooNkGwjU4jhdX4PXBbdXwnHRSbvc598
KiyXre+VzUQb/YRYbynQTJiZOU+C89lDndah6CYL0ODKSYc0Y5nPhvnAzbPGpwQ0TkNHCjmguzr2
ui5KmxA9RtP8y4SlqYzj/PisTyenQkK1QSz/m+RJACvaBamsGgaf3T3C3fPa4VGfY4qtx98kaQCE
CgYAfdcsHxo6ypLlf9wW1tDYxhNDgXjTFU/H2ydRcFApxz0sxmozCFlWCNf4afu91DFVZszI0t0k
QAnPhj8um0U3HbHmKHJcB6isnLElmRsFeTmo/lyTz11LIRUBq+fIe3GylU+onZn9w3AetQuf+Wko
RTB70mePU1ZLLoyM9uHZN8sUkDGBnjGWZVO7KDE0DUl7+fA0lpNcz0w3cv5WgD18lXs8N777M1Az
kDGWs+I7XX65PYnTPn+45K0LfdWDum8kBEmLMqvptHTTuHM5ORDDIXlvzmh1Y5iiadThqatiyIcb
YrYU3nnz9+opG3q7MFdf1Ir9zvl773oh4S0FaNFEtLvp4D86fNAMPEY3uiEOvrS47NPr3rwa4w8x
oalJb5z77ZOQGzLPBcINPJwF9e55zxoow1hQ1n7Di9uRGL8UdfYI/eVmrphYS1XH7aJyo4aWCK6+
mNvJTICmxkwJFj3ZMNR5w3eSYgDV7v6yw5hLduAZBzahjGvlBkwMmlSDmDDoedpsL8KjqmU6cpyC
JEk0jC0xbQLFjkJO3LjDiD4VlUVoFtblQyYBPOhsJtciQeNRj1SYnyYUl/gPMKM4qhfvF/aeg9Tb
boleMiWYepJnQ4xccY96vPMtDT+cqqP7RJqw752te33e4pfMVvPDmvxLlSbf5pCvwcD0GaWLvHLa
/XPCKwnVq2v1a1/mSYJ01fgN5+1SYlWB4aBlpL3eDYitLQVyrU1DlDiZwzqKOnuCBTnx5mMv44KH
TBY18VXOO7vkpU25hyU2aEN6TNybVkCauTM0anfb6eTKNQTR2Kqw9ZjjxuaEuPDMBSV065avtlrb
rC1TH3Btvyedze+YfTJpZkTKr3tlwqjsN74DQ0CHFkI7DmlBGk+hlHMeBhVq86kWDVjtHQH8OQGb
4ka4WgUkZnI93kYt1O/rpJlTGFwCDezxLDvtWSBV/m328wajUGkq+V6spvXVOMHnAG2pb4o0L19I
RWGx3jhfyL2BL0q7FnaJpP/tfv/sdEa0oQb0sEwDU4I7vQ+s4lpGMDc1/4035NypYWvzFeALucIi
iBSnhEJLflVHNbSRLPCU3Sxg0aRDPMMzk1p10PYB+kONtSaH1E06gDTOcyfoy48IfJR+hW95Ng5S
bal7LXT1Cs8JYkcnSBISnpIf5cGc6QRpDPFhtUywzC1NpzxAM3glvSZbsAwNjquICPrh7VNaoxeP
Zhl16YJ87WkaP5rVxyZN5YAeWXXcudIGgrkzQGuLl7JyEJqJnrXO5HzYHjByRpbRXkW6TPIKKZvE
lvcwZe9/AQ4ycsUiDkdPMEeMeL2AYCE2So//V9zImbs8Om24dy/ozQ4vtBDSMPyzHhLCnJD57Ug1
fhAxR0NrAj++Tv8KgEZh4lVIs1boAjBCzzExDvu2MmemLjgkxOewRXOszfYjzjt4lg4ScmpCI8N+
fX1KPNzvf6n511ccz+hwn8KQk/LbVUufVr0IIx4XKK9fOVfTaWIM0tIdURu8oBwcpaYUpjsTZQ/U
0O81grPZP83VT8H+PtayP3v4nUioBKTRl6m7ppoQOCepfaW0kRi86GQ7k3L1JBkDRk9OGJqiLVsV
m7XILeUp/NidRVagni7KmmvR6F5qtgHwNFnyPyERGFx2BUeD98P4vW26Cz/lbFjMr++WwUmPSZw3
U8/RXSfgy6iUu1KbBnQyyD1/YiWqZJICNEVSpbzh8pndpL+Er/BaICoi8mvT6T29bVgJC9Ug6/go
kFyE1c+tth2uCeYmDI69H457da8X8ua6ygziZGaXWil2ZBQN8J9fZpiWHuPHNFQFVwOXMT+SIJ6G
o0XpvsXEPizYXYgegiOwocF6l64QwyzLvwfmC/Wl7gv5SU9kzGb6RNCoL5to8TOrZOmk9byF5MJO
4W/H3jJcp7NlEthwSc3JKpK81fEgPk3Wfds8nroNuuVs0EjTR82lVtY2Z4r8fiz4WvgsdNr5cGUk
G/A5A6MmY9mtT8byCclRhJ937dhsgOP09ueRHbzLU2Hc9R8y+Ac+QI7ROaPqh/Bb22YCzzK0/6R/
lukqzfPik0dFQGJWcT83+6BeAnFCPbzKkyjUEMTAADeXCjYrRqRefTjZlbG84yL9eJMgAIExxNEE
nwAIbDdiykM8X+B5/IOgYi75MfAsWz1ycFEhbvgDTPGI4gGr6m75FyGYiZsLTyfsXSd+m9hkbDOw
NeRt46QlzSxr+NtQG3gIyAMOCqrFgY1+wZeF6VvufZ8OMzE/dtSR0x7MQDU4TyToG9UvOTAD74p9
fY/dcw2GHsnnZ2MS7RXKEec1ilo4YQCgrchouSRen0ViVFZZoawOcQ6P2ZRSqmcIlS1QeAifgubq
ewzkWS7oHdHM843GAk42euYv2mMsZPtu5PNubcPd67Db7s8bsl65uUVxsBQ8pBHMnFJJXVo09Jzg
uZjT+aN1QVbuVFsAIz4uY4VoIrYS5q0uxW31KCvw921j2MouC2SprvvE9RPBDxhgHQHMUPmKc+ph
Oh9HoEuRYl5l1+Bd4BAfvjjByAjR04PqZ03hNBCuf0IJgP7qe8nd1cm8H603LBD2vil1DiH3WLec
hgehXXpYbZxwCsBFt4gkCTkX1krdefV9++4dTBjgCiChtIdWmFvgZiTbxcyse+VgS3FrkgjF5pit
Yx2OrvDq+51i/aWApc9GmaWMu6QhDYhkrcuq7jDsB6TofsL5Tby+ltr1SzmfNzYYhY5vMtHdyudG
XiF45DWFgUNZ0m8GtLbhlFuqJlyFquKjXeMPY/ZFVHtlrpitgK0eMOpTO2O2t0NMfbBYSwMJwvub
1LtsLa1LoqZIw8FVkIoNz3TfIKNUdd2tSdAfOQ8ocIBNIbTtHQJMJvYvNLWmoVMQ3B9v09rkl+Ge
KVzsiURDSy5fA1bYVeqeyfLw/NFHPnaxJQBGso+qkSaiVIWquYlD/TdFQm4xkUZeUnWnlC38Y6IF
tOqpC4FHS+Kqr1FNeah1tMOx/Hoso0pDiBtc01eUHlira5BwPYT8eEZxBvn9/8pAiZO2zjJiTNkZ
8A4Qgk+NgMF+AT2rsPH8hkyBKdaLELzN/7fYTePdv+e4gdyLmo/qBb38TRrdjIJGEK9QEnhwjK4U
mhqBYauHydQAngmJ0gGedCcF4ZeuJWPEPVutnDv+a2WauhQZCwdGTRLfR+3HEF6Qvs67oECeIdNV
N1q6uX1Xh9hF9NXCjgegaChUVvYA+z4UevB0sb8ZGJWwEoGlceGghhT2gvna3KEVZHPiJa4XhzUJ
SwcpVIabCvWVN8hNqB/gKmtrVgciT/WU4ATyifxcuZuBHNQWGKeBJVnHyDLDAbTd7jZ8fUKPXWZQ
K01rr2eD1hX92K9PB5YSZ1BlETtxlX9Za8PIOKhZyUUzf6fgKCsHoxAjEDVzOY+KAsAL2ahMdK47
R3MAgntMjBMq802401n+8mrFZI1+HwCarsvwESKab1vSkQhZE523t6LApY+yROp7NoNWhcUW5Gya
A0wOyNLkvPYgKU/ekhyNPO0KF0AJ3oMaLdVgmppL0/1k6drJ3SQSgMOrfEmRnh2hgkM4EGSj31C1
f+o3xaG7VqjGEZifRDwFTPHwE3YdksaRXNPqG23xZR80unb6ssQIYrWTYdgXE0MO6cyuP3rBkxBi
evrIX2/prSS12EKb2mZFUAhbRfQYDof20OCFdz735GjMNZ3YqlrO5kI0HMNtF88uQIFm7OYvuIX/
hdjn2BCRQdYqq8kcGve7gWbJx3vVLhJ8Fpic3ypgpNyOB6OgIIgzp60gHHvR75UPjD1atI9WoY8f
G8Vd8KHcJM4W+mfFtlI6kld0p1ntR75FwpvfQa8YiP2SuSt/HLxchjXCYr8/Hs9VV2WUy2wIWX81
X+HVPmTrgFIFWGMf2mEYhTYgVFCWXDTH8y73fhLjBYj6EB8Ea2EzTQvx/cVm+zjCwiPVSWEaMog0
PMx3QEzBlfeLL5h3jSgjiaMjLPgpM9DxsDc0i+wED2fY8UDaAPUmTVDtjuSIsRfA0Cd+mgFE3a+h
vHnyViL7pTH9TUFJjF9U1+JDEzB+2MEyMi2taOzFZDUKUYAQcJWonLpJNb/Kr43L4LD5gU0HJNHL
hj1D/dIkXGK5v9QqzkkXktcHzpI+yguTq3znYjSdVI9h2JBVzNJHPdt1d9xWLvsvNN1n4wT3X5SI
ywsy26rjuwcV+Udk9Jk3CA41qknp9Mi8RsaHUl/OKEiUueYePEtiJQPvYuT+JfDXphjk9YVOE/Sq
ZBtWkZDk8E0XlwuHiIEJwdFLQ3b+1W/72uTQFqDRQcI+etvd2N/GLSQHYE40Pbixj4ioU+wKUZX1
YmZnVJ7b8clSt1okW5IFze4OvXROPiuzCLXQCCzeElrrxGD/J4r2i2LEuSLXVd1KYcpE0mXVjkXq
gtXz4KO72JRqH3qdFAqCt4Zdl/052Zu8z77z72tLRrO99fIwjJ7RG3miSqGetGnXgbQQ3cpT+V0Q
GUKpUp8cPsb2asshxW6pWdAOLyk9PI2BuEO620Nzjd3gmX6Kumn2zwLs+Ao0ou0h/6BIt5+vg5BZ
0qlpN/c4FE5V13kKJ9mn6HTebX0lksormVKVhwPGXHok24018poG7sK1qvfoB+ljvod8TeOj3Yes
RlNaow0Wy5SF7iL/chwjILvfF842lgDytLW3V9nCrRpZSgZRN1al8U7nJagrORYpeMX9ik+YVait
Evsq6VSXjeSNZJBLWADLRWy3LJwjXqsKK0jX8DHL1TR2Jzz58oCIMJ3PM+5NXXrCHVxfJHWpoXS5
um+swk7g8ARE7L+zUtygXGiA7ROLDlj20StbvidglTsB4Uy6dgrkDuRbH8JY+nFBnkFjbOcau4+j
9Dyp/08O4Mu4DlGMT7WY5TX+OBpNZanwTdsEJHCHj59dD3uLydKvqA+fV9K9pp5Xp4+0aytFKtgS
rdb/BnoIhQtgB2c8BLnsxS9NRUk0a4Eip2uRvjzGHFkWiRxMSizeOfQeg97hMcu7/3WPuRj3FiHW
2UdQiSXT7q0g0HF8hWYKoLMER/22cfZpy2nbFIvM3M/qLbYUDUt95pZSmmv2fMNM2epKNGFdtSsN
RYx9B5LD1DqAB9FvBmiCZ33kqUD0L6qPAJOeQfhTnL4TRw3ZCxpBi4+dHJ4B43kG6hbZnaqN1rlK
ZSkhC0HyfxibPzm9KxvbftN5cVGeEtMtZ6dtzjQeHkvK3dynA+XmKlINMrTD2AxFguuTdvQgz/Pd
CYHuANJvWizHzo7VFsunJNi3hsGVOnmBZQdm/cnJCzyueCjVvJOxS7qtR186XMgT7lF+vC3Q6wUI
PNoo0ThyVOPeE0VAuk4OoLtGkDgmZpC66gEd3im8YfaP4ax2QMiXkGQtzDZ6qaGNv+olEi2lGc5Y
L2JkzQ+NqmyeLtxbRsBeNYItQyosLtl8GiBch15KXxaKe7FRJan/usNnaYhuHyuXqoIxmPf4UxO2
DogkW9f3ID02Us42jowtj8pdmBeM7O/zuDx3UeK+U//pd1XjTQTLGHunQiX6V7X6hUOZWx3DUb20
J4QjIRnF2QpCB7mf1JL0fAQ/gBFhOuTs4dmg9xMRCLgwheayZn7b0MWM/OUryHARUGOPNc5pgSyj
qpmQBxvijue5EtiegTG+55XVWPNoLnWAr5jFvMM+mhbhw/8F7HJrpbapCWKnS2K/cu/3VqG+UJX8
R9paqv6IvYwNV9TEqGAdgqWzPvL4cCSWFEIJxkaVHKsr+E1lC64fMdN0UJXh/28egTsh03od6XlV
bRcViAgr/nvdKJk7sYVisg2+KzUvOO1EETJwU0jLVgd60B0cc7h3yn8qgpJqPI5fNxEpvh+rWjxO
UQ82U5RpOpj2psi5KW7dPGDph7zBLPEKvTHL9qdezGBN8wJ2It9TWcca4NrgJWksntr7FtCIUOmJ
GyFptXn1Q85LRjAdpcbmHwsnftvKW6UG0VA5M0s0lkXQUDStJ1StwHdCceGlLcIkFnTLACylOTS/
B77+TOeuZCC7Ssmru7qnWG1QArMx/WR4zjbKdFEcqRpSpaLuqwcbJMVER/ddR3+yEXR49NjOv01L
EhVpQLqWAtqyEUZyZgpabqlsyWQkTevcbuLxUSNTpN0YLbc56ZclHbuJyKlTNpcu9adpKU8J0wb+
edl0mDH6GEUnXYhfccwSOk0Yvol6g3uBp5HABBHPnFSP08GdyIDp3IbBic0TM3jc3iizQsWHUVyB
Lvvw2tWpMeWOdQtM0xuluGfgG31d2rN3iFAQr3ZL22k/PP32uvqJWwdcfu0Qu4vGwtwVt8mPrPS/
T2mWe6B+/MC2hbQUepRRiCI8G1c1ITh17YZidhqurItE1RURJ9sbIGKInkcf+v4CcAQGwYij3Rwc
nsWrHFtKv33aWS0vKAYWXyhWqxysi+HWiOAjDMoqbgLGXRMgsQzAsODrRaKuEzXPVv16PMp+meb8
pa9VPQsULea5oId0HNZ0X61o7SZ2r7tJLOLGQVEk0rdiY5OsBdCURuh44B7WRwHp7lYcm4mnYysj
eJJsRUKZuyq9QuZ3UBDNs6Q4FK0H+Rdg/BopejfYxooM9FJO7JQtkBk7DhGDZLAWmRLYwznrVtvj
g2QpJGjkR2H4L9C3idcyBLoAwPe/7xiGgh0rYTZJ5HMTvIzKZAG6q1EYSEb9SxSyB29qtSGOTf2i
lGKasOSPiBnDdDOMSFnt1pycGuzokcD+JTC9tqCiHFh0YIPHodapnFWAvaF4RcNbxFCUZw+0W88v
kSzsJZsqpezfChCXHEpWmGP4mjfjI1tMiLJos4wqK7S4Z8yM9QiVLPA0EIEvpLGKoekV3MLjsks3
OxzZPK1GketJA3Dki6GU2MXP6ppY19a/ycXMx7ntMWW0/P/WMq9XJ9HsMNRAlci2+orvfVwl+yQG
zXaRapb2PBuaahgU/9c42tE1QqX+vdIbgA+7kjm9OIFHcIgWPKGQ2Y3SuOYmvMhVf4eXaYMG1LyM
2Z4Guk39ywHRy0NbvUWTmPyfZF5KTY+8M8d1z6vBeqUVFppUjijWsGEKtBLlIrkUVg15A4XBSodx
hJxLTSXz6eJWTZ2WTDKMyhEQny+AhjOfNksrcKiZDNtdCuNS0VD0ybO7cHwFaMYMIR6YLzhR467b
eNlGM7WF5d4Q3ES4Tn5B86wurlEEiD3avA4D412Vp0hr0ZsBJYRg5ofQgXtnvzJvpsfLh1YtjcAv
rWQKC6MDJgv+uKnSgmFZsliqI2qgCJEpWb5alyCMVAaByejrlqwsgj8ZosTVQkwP9uueHiJ7IGh2
ivQKzFGjXHBxR3y+IxZoDfjesfQs065Osp+Gs+1q2U/CE4tuukD96MebhqSTo3AAQNdcPlRi/hiO
1h2IUekhPIb64FKT+rBe26cdQr+7rXxetqcflA+4TyqoO8+qkQ5z267Lh64bmZX3WgihCznV3o55
rqHrNSK6sxwB/8MoE0/L3uFKEdRDnDuK8VB2PzKpwjT3MxgGVXi3RE4h6RClq3v34toqIIhS7IuZ
/a2p91roT/pdpauSOkC+Q4v+pH5CZISLlVTS7B444lQdXUoBauvq0OlhJ/3kpwu5r91U2cQnIAxl
EqBo2zQwIKsVi0yNnqaK5dir/NLBI28xyK9x3yCJUsttCrJF/PKdSez/vHLHHiZVLgqJ6ypoFW54
2jteNTbt6u5aHpsr0tH64ppCPcYRHRjWrTx3N1XQwDw2oHZtidqU3bMSmu9vXfXhrzpKU0ZiwwNs
9WujfSNfXuNrMyzmSIiha3cdaHTFIkAHiLXHZH10NKU7ehO6U3y8OrxNjI3LBAtVjnLbDaRvvuNg
bES7w4QxrLsjx9h6btUYF80vJF812zZIUjd7LrP2FtJyN6s9Uxmjz/jNKmBmILs38XOV86HeYwet
o2gp1+pCu2jldSXs+rHDohJKCRG3Hj9PT5v034pUx8TlAP2RMpr7EHox2csvV6l067hecnSmC0EE
GJan9jDd+oP0hpe3DhbZPqa3mrXfMo/YdPQxjNFbjWxQASGxhVzumP2PJiUvM21Z6+pb9A15Jxf0
7sXi2toHjngf/zapYfMo62FyaLcQEEOU/50eLO/CreLiifGkWVdZ4Ng/Qfh4a8BHiq/Zhjx1X3lg
f99VbiMLie0Rs0DSu8bEIBgQ4V2wmynJqe+1EyplQgQikIHNf9bGZPE0f2qH3uHquv7TZ/LDJ2Ui
nKfj8XDfn7oFPwPBncvZ0zB74lw2yf5VwnPuX7EvpB6U3HlC54ZeDNiE1HreP6jvnt0R2KSzYQo6
ulr1BKVBtmlTmPTJrhV+fxnrp2uNgMG+gu8liOkAEYP+Tv5azcxVkxlcXXaMC0WVhL7l3NZOSny6
sjd9Gp6yNPP+zmdlX0i1CfCGC+PlVyKtzQDBd1cIsmnXzolIytmtoRHpcGv8VZvHKJU+ACT3BgiX
Uh1u2IWirn+G0KyTlEhTc5FQtRwFLmUeetslTcQVxkAVgz6InL/1ENzqFLqzqiQqeCzIzsjdLnX6
HgN994VYW+tuFqJ2o2JJ+5QjGGhaiErTs3lb5w/2BOg4ftc/PBAkav1BkfuLq6xDV3P2JSjVqOK0
X6jFHdU2tHXs6ddgN0HxezlJCVzsQEqyuDo9aCFJHGfegcmES1ppyWSxZ7caD7SJmVsDuGfgvCwF
/VlwPgsMjduUZR0mn0eKZhIfIKMLX3uFCguL8Wof7MVGI7xHEmmP+8bMoFmn3X6iX4brGDMhoc4N
duCaihD4SG7Cf6NNnQxWm099RhHgMOpDsVjGgQoK1sdF+Bx3014zC15hOyKExzi3D25fo4f39Kxh
jdF/CpHKUls++fP6jAdB22fvhCaaCRvD7G/9+DLksqTb+5dG34MwlJJAR+qIVykRzGkz1Bxtjk/k
0G4WFcqtpwJEpxb+CyOfvNcmTQyqoNofBVo1THgJdeTmzj2OnO/qP6PwhqNqieIRM9qx7P8YnIaG
73Ds8JB6KL1zZ3BkBB1ow80s3kp1OSczS7/GQKGJmUB+H28s2F/n4PlgQIrU5fiNYyjNYewylwoK
3gRCDz0GHWIgPilgJY7QVyxYR/VWmIVpCUKgS8kcl6kXZxNC+aWEULM1al7aycvykmEVryPvCZ53
3zzG1TjOSwu/mu9OMpHHsx5nbNE66ffndofU8Mki/laotJe4/1nw38JHf/OIh3qfLqoWVenhOnTR
SQIxw19IMdQHJIvrUMQSr25Gv4Rppvb3WEQkexa0nXcLXBvWs7rVgFTZGEZt6d5oFR0GZHDA68YM
0zD2tipsLJnVfvqLK+/ITsOG8K7+X1bDlt5M5lQgfS9BEnf2/ujq+MWO1NwmKx50D4ozLjvfmk0Y
0cM7Tlts8IAihZ7RM4Ui3zOJcq2f8E94Avqs7KuO+Ztqn6p6NVth6SzYKWMwo4g7SCZCQ2NUhhJx
kPnHVxDT/onVHX+xJFGLoa3Rh27/CeXajaJxSAdOu00ToglqTBzpHGGYo19GkhanF4CFUjCpP+Yh
31VA7SZrMOULFpmDMeTZPF9YPJLm1BrkLMjTtEmVGVKCsMWJ+wmG78Gmjy47PiRPyxredc4g1S84
P4eGNTF9yATrINySR1K5HK0uGys/xKc+qzOtHEaTBmqnjNp+ha42ku6mAFHJKWDOvBvcX/maMCxV
gzWWieWDchChtbiPBvVrnayL6EXQu9GvxeBbii89WxhIq4S29uAlYqAqXSUp1RQg+t9WQAbBIMT2
E7F2N1PzC1ynQ7OJap7+wXIEukp+S/VN8bNtZBlkHUbC77KRriodDQtyMr5fVvDyhxWjQPgtqzuP
pPzKr60hkFyXlx0+id0TXynV00AzG9kTlMad3FJxm8g+R2EO4e2SzkEoFenw5WWE3rjOARbGQep7
eCht1asfMZzeL/MLoOWsAczTdbqkPswEzGIq2l8elgogcHgtFMhy418yi3Fh7nTK1suP/HccRAvZ
R84sDL7c2m/WFZybz5YFTyhqw4wZ3Ey7s4em5Z7ky2ul7f22eqzVwyYqcL1tOMrIc1QmZzUBBzn4
544mJ2bkgkbLALz4+5lKtLZqpDJBhoTwDjNlBM4+sK+tOE1BvwaFbRzC2MR+QZNIRWUL4gTBzFyy
D71j0RNoIKu+N0v1+s6vcR35BVZBFs76fwlj4ENCiDu2Xzt6JMXF8Gdm9iohGsh5J5ux6MCo1F30
mobOyWXAR9x/ZyyLxekwytJ/yT/WAQ6XTArHVKOKdJBAnuf3tOoMmOYWCjPNcBYtdqXFl7s9qPbW
Pf0FDZgeTJ8byYSy20dOusdkxhqyNYx6HmLtkriC2evufDGbhiiIoqAe4zHwYZwoVRVGZSuTvtUt
wxkIp1mXSZR+OZjl0vqBwk4UOSOQ2Ye5i3ye1BuOasH9GKmrGJYt5aCwI3No0JgGLllyJvHRB2Rj
1JcdxzanLY+szSX5/wcwYsgy6NRODF2suKa7zrISMUu7noJSONNibXn3/KfMuGHBjUMS14xyaSUB
YpHXBTnWK7QOk6pQ/I2tt7Fr24jvLQAe+sN2mSf7yS4PhPRszMYwvV8pJZLN632VhjOLJrWbTDNO
xd1G9BLIFR8/tkiKW5xjOONDbza2iwEUspRKUsW7jI9JVorm6VOUXQhsSSHaR69gvjwghaxl6uRW
RbSW3QoDv8b7lQRtkrdvbaOryHsPttvjvRjFpxPAzFXWnGUKtAnjV+9A12nlVvsKz83aF8O3qI7U
E/NJY7vevbAnIyGOBcbB8wmbZHrOA8P5JEMs+3Na4eg0M7gc+kopc6BrQYEcI/qhg7ea4iIA0EMN
C7zMmWMF+DsOsG041TkMKjNbeWNlsD7HEqFSDEb7phcP1B8mx22l6/ssoxKgDha9dthbsprKJNr5
CUgqPwP9bYTdj2TUXNW6k6bvrnaFW+XQXEZz+aTkmxkWmXTL+7/GiJuW/4oJs8o07sSiI0MgPVyk
Iorca8fdDClcwX3f2lgZCDRzhbzvkHuR03FOpHa2ZR/opvuYZiZTMgBYSGHYrIomdD7MOnkkA8tV
OTjm0/D9xut4kVPkDCm41B7EGed3uH4biekawujJSFv7NPVos+Ak5Ox+4mf3IdaQCRmzoCnqsdvz
yLG3gOxjOgRJlvBTvxvOsD5LmixIixM2Kn9AQMNhOrHOrh1oOMgYM2qYF28LKlRzi+QwLxG/G8zh
0WNEKp/R790LFvu1MUkQ4tofpajCKqepAls4Zt1D/eEYYwFEDAizPKBx6pO1D4lhk9fLppxdnVJD
CDwaStxr6+LIVjzJOu7+vbHUPmrcnJm2khiOKizSGJ1YiUbutvTWlH/tbn41Oqpc9bA1kA/O9sC3
1xKDaVPD5Y2lHkgRYjOAW+S+BsXqNIEnRWJGycXlua773iKDhkl5haaGEGbCY3nucDYhjH2jDcO1
vEqTwfL1gCFWtuUeAouLHMtt9ysN5IVSC+CcBBUgFbF/u9KW29A96+W/H+SyMqh3XIE1vUi1rMuu
hajR1b8aYEswGPBUNt8ixzzxvtRBFGkBZXvIR181NeVjLyeEJbFiCXC4ZwJivDRvwWEPJkC9kLoZ
3c7dRkDQm18vpmGnWr3KB53NTPgEazA286qATs2IAtCMpzzArvkCNSSiprBys+/OWOHgfXZ7g6nz
kfWuuB5oSpmN8M3bM0TfJFcLerlaoNHwPtCjp2uqCxs2mm3vpDRKAwdrTgdhOiDImQ9PFynvHB8S
+Rn+5hq2dM5S9NzTauvQ/Hdz/FWVJW3B7ElSy2hymoacHJ4ZKe6pVs5opo1pvAZqSPCCAlPZGZ7K
vBt05MEPdrE6IJQ1ZT7iXFn4wHIR55FfVzgFut4DWZRaxtbs6Fl4vg1K/kx9RqiisnuiVP9GK8w1
oxK+HeElajtwVcPD7fKxwIxnZpOS89yLeWhaReAPW1I+eg4uZjeUbSnAvK6DlUlfPc2waOQsmqrV
ZrLhycnIV3mFrMHaxuOJpuLXBf5CFND4j8YyvdMaHrTwFzfBoT7zr3ZqRrDwFtNsbWiYe3RB8vLc
whPvjPLotqloWbVI9WnFAIOgxLon/g5hViIcKF8iYzomrJ9MfaNSURLeYOJHJwFHd8gYoA7Yq3F1
wjxlPb69Da/LLsOPcKfJP1olCjAJuBK+F/BisHFw2QG0pPiFzS1yHqPodS0RlheAy5s9zjCCBqDg
U5u2z+ZJwfyg1yNm/ic2H97DUrMOg2P9Ff6SdQ+4r3OKAD35Qgjw2Cs4UP2v9jVAry6F1Bq17goX
kVtqnhR5nZfHhrWHA4w9QC9Ivrbn0dS3onstogixfQNGteD8FdhVYn9D5CincTuVHlilaXNugDD7
uFQCGp1pEBK97csNmqe1V2VxfQSW6g34xsLCa3TiTOvE2hgla1xR+Rgl82LPpAwZrKnnVocUsWL3
ijaCPpJHP3taHBsRBaWjHHZk9BKRnyOsAp8U0dMwz3vQHhtmD9vK0ckDmqrWV/D2wjJFIo0bRogg
jCwoLPJl+L3FSKPjAm4CwqOuOn632ubnPnHFT2eh4WHJ51nJRTMkHZy73sLEVicsk9locAOQ3zys
Y3maZlKFg9gA9Xgoyt5X5QY8hEjQfGaXoy9eIbCA773jRIr0drRrk8urHvfxJPQfKF/hV003kKIH
QX72nG9zfYJk/bhANJh73JIB0xApvA/zVbcoVid0coySsi8Bkk9iZQv3d+MfDfVSor3SPP+PtTIF
FfsTS1ZMRt4M39c9bE7wjGYj2VyVVq+bXhb3MyDhpb2H6lXMxERS8z0dQDndygcjp0EWE4lWy8X8
Rxs9zfgFZtwUZkrAbFxbvOvSQbEwjl+y03H7FeOriZQrIfFlEBe2xB8ntdsjuUO090o1JX9QCMMC
t9pB+ObUfNPMwVXw0Ct2lsy36VBjLi+QN5dBptiJbAqgW/Wgr+Ohck+hTr3WCnmUEApioAOCTtqm
JK29WshMTKn7Pp7t9ZEMMjguCMZExwRPLthTMH2coXxkeNF21JNy58QyiJPau/Rh1ezZJDvzd+pk
dvaEJlyTMtr4EyUL4UWjlihWKPDCPNfss8Oa9hKahZqb2L0UhLNRTOTOBJA78vrE4Q7MLXuGgMYI
LBHtCIa9ccM1Z5W6uvqDelCmD0OvofiyZSK0/1ZEbyJDY95L+1qau6o6nCSSwKDepG5RZI/8R1sv
Q3eWbqs28zp0118Bid+5O/iSHjgLWyLpr5AUUwNlVs0Hc7xvyDiXDy98jZ9seyjQlDUSH1eAVowC
WqAXJ4/7es1FD3cG7P891a1h1jNAWTZ7JpGacP5KILKgOd8S/HG+XjU2PKGZRGbQQqJkHxDKBGUU
1rnBk8Z9TeXcyIqrkGKYlSQ0LuxA/iyt3U+BsPL/J9rGO0XnIZUZn8OLOWjYNbYJcVYeNvKMbuoj
rpNCX9AY9ZQKg47vOAkVmgVrs0AOthxk0KNHI/4rPL1wuS44i7rnXKqIUrI6DsN38yz5SizpJ5IG
LITQkKFqywwSsvm3l76LHx4COww//52Hl6Hx1Z2fFDeBzw3B+6ZGbCz8n3w3tE5rjEQmagE1+K8U
iLLK0uHVjtjs2n0mChZlUhJfKQVq+8rdJrk5VIwglC0c/C8hn2jKlfwLZArrWWiqyjXjqy0mI+MN
hzom7t4sAHDeU7XEQ4QgQgalT4PwmTLQLIRXV//Exc9nn9FnQX6O8j8KoqOO2IpbHSVpke2T60Cq
A/+rynKsDsPx0uciEHaWZsNpkTKXo1LjzdinQvYPaCB8/hsDrgh4KBXI9gDRFVrNAbzjpPkiVsrt
lfoMyAdT6PP7o3PPcvHDhmBzG4Oi5+E322/KDPN2G+BtiUX106Txvurs5ojFqQe3F2Mt4xEi+X+q
0u4o68+8geel2fFF7REXMiNa5q+uXhmBcHf1HjZwl+9JMsHoaRS8vqp83O3P7U7xbJFnCNljJxHm
jaqTK9yU+ojCSlGJowLXLyvn7oG3wtKIoJxe78unF7wsCbjCOvLd7XDb3qr3cCMuKvJH6E4pFIWO
IozLysMaMBG9T4sOolML+4Sm1t/ganUEOCZcq3fx3UzhgTrE7Fcd6aF+W3OMVzq+h6+hrcP0mFm+
34t59eo9bF5l8Uw1yoB3XTncI5bGmp0n7I3Jt187hebbfcW5dJwOXz0kqKJcb/a19u+0SQNSKZBj
FxDIdfiuPhJwHRhhbjGWigFjD0E6Mb5hCjyfDWuebp49HTU416klqj5IxhlZoTM1GWGzTOBOry9m
JA7BLSSG5EcClKVyWVVdIUzpHCZv8M7Q94XV91kKh89AZqV+IgVP309IpU71ewbLoIcOc3xn0O/B
8NKmAMR4IGed0fKwmNAE6WyzwdfYMj4S9U2VviADVXxFg5fY4WC20X6gas/1G9qCg5Q/L+n2p4V9
1h//gI7VJrQqecVmE6ZaqzdrUJt6ow/NY/G0hDbA1ImW0ZlbTTkJtQAKAtoHX8fpUs2yKj3YUasl
XTlxHa3K28dnwXxJo6u6l66bcix4GtxfFAoc2fVQ9h5Ux+7ty33+0vyCW/TWMWAIfSXeuSUK1XdM
Ti1/ndOzKJojvS5cqdo4Z4epIwSa0HVmsr9cF49hkWMFfrfWhHbB+az5ywEmvcjYEZmN0ed90uXh
oWhlxTAfsnWn/pgBydEtrX+NnDpO5mMwWYNLhY1lLSl0heSSs0xsG4ftJ9dpEAMnluC51kpc4Lip
12IZ+GH1akpzbrG6YJ8J6jeGODA2LtCHkuCATpYqSaebdfYI9+WpJiKCTxbavtcfEiAD0oGbcxBp
4zmedO+IbHw3udwf0E+SXCFUDlXxgsYuKBCjVf5a8GcXvlPJkdKeTwbNr18q26+Gb8fy2bNBpKEa
uEgP2bJUbWN9lZsIyQqfq03d0G5Mb0AN4gDCGDpE1Cb18OewaDf7TecjmsmDqrRZ6JX6tciAeOA/
ASO8+dqcnbYjecrMld5+ygeyIqe141OxPWW1+4F537zmNgPTwl8n09x1+CK5AIuCvIHCg9+Hx7uA
XqNAdMGze/qe+HEv+P7JlZdcrnvCMz6RI5jip/k7CERNKituLZ5nD42wapyu2RTxzcYpUJ2zcy4v
DXRszhqpKv2+YLewKHFkmqK0b/SB1fVKckn1RlgvC3G1fEhq8Q3GChx1hTbKrjdYTNWkjZFUVBX7
bWASXYYclUovBC9OVzdjn2j0ZcA05mTCUWKIAVxSIYaKiYflxijFGE6hYFsZ05oVUWnLoeUQjg5s
3Nz7eitjQoIEKRf/FRu4HVsE5OWteHd+Mp2cCjxRsP6zH3f5S9N0dSlHepvnUyWRforLla45HMJT
SKn1uamES6+fc61cMSWlYWxj6kP0BOo5kUZHUNdYZRbG7GAvGhkjwx7Tp57jArLDQ4MIYykMdMBI
90HIXthGPuvAfbG6TkJxDjwu9ScbiMLS0HRjaitwc/lwuXIocohRYtHDAG9G8+r05ABF/N4yeHGG
5bCmWehrM+XvJQsnNkgvhA7Gi08F2aljOv/Owah3Ni+i5VNof3GX9D8sMlKG8Zfg/138T0HkUgFE
ov/660bgGD/Z2RffbgCe3Puu84IBTnIyBd9YVuS+p/LWnRs9F6cG8Ux8WgIDy77EiSrwdEBVmF2c
ttJMWZFf6SrBkBEn3gpEFcxIW3t10gmiyKrZTtoUY7fowLk9DlIDNGIOTFkcGP5Msi/2BvO7WbxF
vGggWFnsuyBoitq7rjlhgR7TVkEJwxiXujrSzsG6z8mwi8rm8GMFsVi0JnmvSnKEtTpzHWD78E8W
6z5KTsjouohkxcyLiX0syMxPN0bQi+mv7bLCjsgRsoQfqxhRzojuz4DGjjYFZTm08uneEo5kX41s
f3+YoEtSUkZCTUQQx9HH5BelWaMu+lj9SclM9uX/jc8UX2yOntL98myu72IYxBgzC5Q97U84ABhL
PR/HCUgg1ZdVXB+pa0eCUzVTJw6qJfumspUPwSOyh2d2MKSVcaM/wJQuKE1Sk4E+1iHhrC2IW9RF
xxPtzcVAaEAsXrrX88t0FWVBObHNNxtYf7foFnAZn4kXuiRwRU7bO6sw4ZHQvNp5ywhJtBQJtU31
V+axC3TulXGWNFRXogNzzbKRZNeiQ15NggqE3ZbNxmaPv0VmS8D5eaMKis/4ODzm1UdcdwleuqWr
hewQceTjObSQlAq8TEBmFyKwvV7sOvhbT1cX1AQqD+u5GaK9V3uCqLB7nNWYbpvIMap30N1cRzNt
uU/lSAF+u3dU9e5Ff5Bn7iSXGdYSTgTcT4dKRBHqQRJjynNXGEC1SOL0i9px6zkEZvovwMU8gCUr
RQG9mGNlTC2hKZnn4V4WM4OPwWiu4/lQn0yYZuL7Rf7DQhZ71L7LkZvj9yPSmBJ0E/WW2AqnVRjf
Swd1V4Z/++NkJKaQ78oBlIFlj8Fwo8Am+0rfuYES9l7SlP8FzPICOc+KO6N9OIHQemdFtHoJtGj7
R720PNbMh3pOioa28q3xVUGTaQxL10w/sUldrORixR9bAARmoB3rmLHPy8fS7od+zcWrjMnakshu
ro9kWxnRdCvXOOyw18dQS4KNEoid08tiuN3yN5iyHz+Rx0mM1JyDHJ3G+MYKDCYY+IHKb8aAcsjJ
9DmGMlQbaOzx1gwNcCBLQlPPlvCppdKzKRGFb/eelLLeYMHBNKWYt31duV6EBhIEktZ61PN/hHdj
h+dtn7oAlzMvq5UJmicDvddQ1J6DYR439P0nIqnrugjH+sg6x5UezWSUsC69eWwAi0xguNlvTNZz
BRkHVblPvoDoLHxib9ZGoqmEePr0y1yi0qvxAYOyMzP8qHnmFPS4rIy0KNArggzm1sWRLgvDGKe1
tTEd1ygPztBYd3Ka1jSRRPa+Rm+5KZRhDlLyO4C5wCcFOIgT2rL4SNrCCKC4bq7/qEjskg183ZQA
l2A8gBE7cLbSGS8YGBEmNdHssiyUjkMy7PVzoogAkjl1fqSS21GAWu94TqVYxhEKT0y02ygCV+5x
UElcL5AfMscmHhS485rNbxOWQdAyAKr+wmdaUNiCsv0PN9HwlFcFVV6ji0S/6mpl2qIX77+oTlcV
57UrJ4vukn7/sKyp9D6WRN/LP7ZrcVoYWc42+Al/qilWTfrtRp9SoCphIvS7KMMMmmkAcW4YcX1x
jM35lYUQBnQFhOstfvc1qIsyhRBCI16eBCdGIdbWCcFlIAeweOClWRLaM/3d/A4MFjS9H/JyQrVn
bZQss0y4WfCeW9NrRjmSd+cCiiSpkFIhX+W7/75QKB2iknm6PveZfIypmOp7VGwgCsqp2DNVYkDC
ocH0MJan4swqEFbzFiRVv2v/LM2XhyAMny5FQioGNarjT1mPAJ9ghscmrJW4CUsvA3tRBqUTohFZ
kjGA+mJB86X7wpEa4wRzJ8WMxPofdOfKsEe5hJPwmViVabrT1nB2H+2pQ6e7NWbxjvBupPc5OK/8
2wP1OaJKi32zi+2T3phzS7jbcqM9tC5vJY97aM17//oMP77BSI7DacxQqsYxWAcGdiZ/iEmudtaq
IguY+fj+uKD5xrpuUfixhocwkA6+Vz0Sm5EYEkKPshZoTDXZ/utPJftqLie3O2IPuT6oTSPzqCDk
8+DLhE89AAQul0tgBIcGUWx15iDC/WPxmpcHFL/uNmZzbiH6l2jCNKQGuny4vzxQk09F6Cuq1Tk8
aUb8HU/Ae5arBiC9+U9+1Xn1xe+NhRMJYRiFEOZXEUbQb176IISFM72iqC18sYuTU9Io9oyvqt5K
W817Lv6b2M+GH5ks36AT2XQOm9lC/8eFdPJKhE6P/SVDiy5wJ1Qp1j2DklryrQSa2fT/yz3T/xEd
hIwQTbpAaL66+piWilErXOk8uMnAseB4BVZFMohJzfr9bNhIsMTgyyVr9sVSuvTHaaqQkSWSL7KD
/jdqJexINKhXJ+XGM6R4ecrGbkVSX4O3scheZU5moK2cr3IdSmroobg0olnKEF6JdUx6m9uZir/s
Mlk2jcbsbQC1jimRnJYDJiuyS/N2e8CnJ99IPXRZKZGpDEtB6WVK4sabCRYZOrhU8B5fVg+CW7wV
6s6CyaBnQPNgakLLShcPXPVKrymqRHU2hH7wm2kCFKZpAF5bFtgaPDQDmkfelZLmFnHaHtx/Hbgp
74OupR6cuxHrg0y8eiBuxe2sycr2SbPVziLv9AqprbWdKNN3BDav9p3BiLlsh8ZcL//v4nOH2Mz0
zClDCM+0CVVDynaO3GS0hXEXvML6r9g2dxkaMGA2Lqyd00nH45vOo0xfRg4NoVOZofrZCHILVVjQ
l71jrYDr3wPQcruZKunJPVOvlDeQCCQlomnIL1SyfQ7t3hXybev+tg5MjfxM+bWRGGzXATmZQrnA
pjhIb+I0g1qzsVGTON+PaXGDNak1jIUYTSHHPDqhizgL9IZPwSWsWWEtAFLw89SxMxl3FxvJQBkl
tQpP3RmAcck1XH9DJ865tDkibqK/y0V8ntc5f9wYDCrcm9vww4Qod868huLaij9fdtR/D4RRUX7k
kSRq2ASVqnuQVsam/Bmwld+RFBOHpBCQ9ZI9OEYQx2pQbu3HGHXkh42X6P5MM1ysMepPVjzOYtQK
4Xa9g8Xk7yoJjT1Kn/PoZIJ8CQSLtGz2YvPHrn/5WvK9gjdiXO0rES0gSLFCVmIk+OqHiW2F1uut
71UOCj6cpP+U1j7nujMir/gUE6c51ZjplubxgtcO2mQqooiIUfLsZn3Iy2fSMoiSLApIYjiVzDnb
OU2OeoTFmTvMhnq/6rBGKYOu7x3bgt/Xvo3Q5Hq1NR/fRM7KeEE+O/BAmwPihbMlA265rUjIgAvm
mFhsy6e9AeE4Cjp8Rbo/SMgQIKTIgoiAygkej7gJlVM3wLojmFWcbXfqvfvGlwz9GlKqhtxvDl+3
Z8dcMdx2zUO0RZ+5+QX89nZAT39m+b29O4cItqM3NhT+iYv5gqH4pbTCqztis40x1L75nwzmtStY
NF5aAks4IW2UoZvJzyPA3fNWC9sPF0hDbcwfM1h6fEYkP/fWGoKsbBUngf/LB6whfQipcP3PWuxm
uHmCfJs9FMNXSf7PtSz2r7aDCW2vW6Az6BZuj3UyTSNJ11s7YgC8H2/4vSr9B1AZbt6AA13fa+Kx
F5u5snSPjXsnmxxAgOSdPC43aWCY2OEqd5JazNPXaCA6oo/FiaGdjRo6TfEFRsDZX91OjsabXWOf
PMNlsSNqOVKVVCd+MZ+YxgEZmzzs7gaRKypZOiI/ARY2Pt++9kGlgoNfsidLv9cg07vwuFc07aYJ
up9DllZb2bGgigBI3XnW7w6F7iREzeoCAblhm7l8GZkjk8625LfPpNpGujwoTFO7vJLeTJJ2bcUi
5CWdWc1nawsBQuGvAmcLCWOdgAtLKs8Z/tvrlLaWq8aDvQr3vu6ZMmCjGIv/sOOodAjDt1x+Z/L0
6+4pN5vBpGzQqRKuECCyvmO/UAOS3WLBcRFk3dG/885PsUsdgGrJG0WPZKTHXtAfSdQZxNmWtsna
JbCmUwpl5aaKvx/ogCOZdglSacnwuPvyutluZAUtbfrKSt2GBaVvmunZwYcUphCdmeUW7xu8RDGd
ma0fP2brItlpnmot9w3OQATZkcWJDvCjPx1D5wMXfhKfxHAGT+o8T8FRJrzBI71X8OScmB5ExSKo
lwVs9ThmFhbEHJ0IwCoG7GpsV4E1l39uLT4gjW/9Tutl5iXlIljwG3my3LtjJkWz+Dc48p7YbUeX
doM2sW5c1HGxZBf6vEtb+GrCQ6c2BR8err1DV0a5GkDXZDKPv/uTWWWIV2xLzhVynF6iipp7jKIP
sYMzcKIhD0IvkZvQ4fzDtrN4EAm2aWFyNhvpSGXjfV5cMni5ukijRzy/oOeODTrc2EipwqbZQVB3
4l2CwiWmzSEIZL7hw/hyeOtzeAXub9YhC/nbgXOLOqYvtb1Yf9s4uDDnFIHpctegttfqxdZVDhhW
4/eJgL7z1IpicFcBIsFqtV9Z8oEmP8uQyLiD7pd7H9HD2Iw7VzESonGQPf1AwJS4jBS5dEyE5Emi
22l4S+cN4XwwwGljZMmk0Ok+wIDpDc5uaRziLjFsEwexlN4fhdFS9HyjUJGJ89RQgUfOPMNSBV6u
dDPhd7Soci0vOOegQB8PgfkHBknOoMuxm4HWUm/SH6p0+wFeolXcPQ1YIduCTFcXUGS1v48cZYLL
RZ026xlgSD7Pjs32gw/dCpuzsIr3298X9ecWo4n3ticTKKsGH+P8B56BM2+2n/jvVXx5e/0EcEe8
y+4DofsUwMs/GD985iA7LtSNVNHPTQ3TEdbzD9Ws7CYRDewrI1CO1PlFpDE7laRxn9NriBM6FkdD
gEZAMvUX/zjGfWw2tEWrd7uSd2/l9HN4V0vOEPYsHKFGn1LUisSdZqPP9XSWftslTu1BYiG6cyhX
aLJR3V2CKg7S4UK78BcroEEkymoOlU6thA+Yb9M2wzDQH9Ffk7faBt2AWgo5URhXCG9jK6nHdjP6
b+b7dJNSY2oDwZZgTS9+ZWpzGO2MoGNTlcsRGMA0eqhKrnSDuzLmHZV8tM6TiZDnoX2x2+j4vvVi
t3j+6VMOoXXfvHdWVpH+Ty8oLzye0LR0LdUTpYBjZQdlM1ebfwENxch45SQbaSeC5Grj5PrWIjUX
BqgJWxrry8z/67qt9dWbM6eAg3jCDEbI/q9UaZDxBqnRJm565f7VymIWLUMCcp76wLErtLBGMkpd
Pfg0jnafPZT3QzDvuH/Ezk9lbZIEVL6sBs670gJ/lIsHu9amL5cBq4Q4/k+peMwijjtZdb/iLbfJ
+hj5Tj3nlu/J8c402SNEHxVKQnaqnLDHeju2b9yOueAjmmNArvRPzRblzJ/V8ar3yMpzkqnr92bn
kakuIyIue6+V2+xitRXPG5Ik+l43YMNvfPrVtto8ziVsSWGMPYe2eWEOmeoYZ+O2VdJPgv1iiLjI
r+Di2jw9KjFehiV/xUXrwHjNM3H00msNT2jW/o35sjtBUVeOChmZYEMtYXD4XNIbpAlQfXmavljh
R0PaSrfYSF0QhNiY1ejoqE+L4IdIM6R9sgsglS3jBq9AMkv1knBm7fnr3PuZ5Bd7Vb+TDZl3u0EX
95N7N5rn/IquPnQ/e5ZqC6jxRtIX6+a3HwQlVxBDK0Rwn32c/jYtsEJinPJOR6qNHlUO7U4q8vTK
N9F59mgn0Ic5MS8D6AyuRsTPRNZeZRA7JDr/1gFbIQhwwDYH1jJLvsVYq6z4X5Hhiww75k6oh6TI
tcUbwmKV3p8tbPHhOR+SkiUsHt75cJt82AMZbyoM1c0xl677puxG0FRLc1oSoXIePHqJlbC2dALe
VB1i2F8oa/MS89M34+MjFAO/Q+AEShxNlA2RgjiC89ah2BjNTXYRu1Hu4XMoY+flEUN3LMhR5Nab
CwrFvcZqO9LQgcYoQkh3YW1FGqf5bmcsn8eTUtbeg/BMMWp0DuwMTiUuzVRfUm4KZhEzKi+RJq7L
i87gJS9a17Be86Non8v1rxAhOtS407UOqFF4/mw/xVJ+OFJdvHaSjyAPz09kuZS+FZjTq+RoTD8h
xGtqkh0E4vUUM+oDj8Im5hzTojq0uoKrpXOgDsJvTY+6Bwi5D27nzuFyph4XvlPN5TOb8rgJX/IO
WUwXrY3Tgd/gNvF48J4DnoRBx5ba/OO2/8Jch166nsVaSTcGZfaCfnBmD3kRd9NjFqRnjGBeOEDb
CPBIj47SQQVSt3kepWQFIvEbYeIQa5iymi6JBe7T2FTddFoIKLaPvB13enexO0b1hDmX0CCfe1T8
48zfp4CqvNuyZDFnwCKnSWceBkNocBCtAZZvY+2igwc0eUQU4HwYBDNfu991eFAIoYSST3vPGwYc
318ypFJmrx10HGTqGRqffkx913BEYNxgk8gBCdtoDTdsn3IUSQV4lZCdHHialSrNWxMEsyEzYC2/
F/RkQf0PEgcCJKPC+/dgwqPb6WqQvWAL4DK2jt1PbHDPm8HoeCc3uFqGdEc6Iw0id47xdYqSTdXo
UHK0enYiT4aQAAw7jsadEA+bTczTOFuV1RlFaIcdsz5fJ/toWt/+rBr7TcgE9ZBT/zw3lzj1NXk3
xgIq8HGBLhQnoqT54swKBdDUXPVkKTtIjFMHvSeTk9V06EaEXKVb5WxVwv6HkdNmcAIOJLrPP1Tn
1xu8EiMme1kpkgv76UMiAs0t7fKkQxWOwbp0S8uQEVx5dYmnKtjmypXAeZOcRp5GpC6etrbHENYJ
vH/FYz0i7ERnxc7HqAm+dcOo8cJ87FtE6XvcjFfL9aJhI0RFJFwFMDLNGQ2avtW+7kRhGDeH+Vqf
sbJGkKB2TZ/6OnLtJ6dWcMpKS+eH2e2MGDmtuu+MQ8JjzMmER7HTL1AfGv+vRs6k/TQupDGvbPfP
/C/DRYo3YaNOwCvJWbBccw9dRP5LvQOqBLYyFyF4GG8lg6pD3dJCNALwD5baI2R3PPdoUjN2FNdH
Epy+us3Gp0BQsGlyuNShn+afkoKgGvXsFsHSkHw0dam827S/mDZeftZgCh0OqwBI2/S2RTCDV0GS
V2y3lxJuYV1acphdGx0NQ56EFtQRtEHPblDS9jV5CvjQpgFxocAmcAQ3/8FPypSuxW2BSMBpKjpA
Q1OqYykJB+bRWfLvr1qG75hHTy6zYAAmT7bZ1PxKmZPt3cAMzRUJeeD0Q46ypVDoDfA/fseTRciZ
/QfScV0IgUcXxYv/PvYTfaGTYIB2cxeIMHR3y0qomCAm0IKyLQ64NdeG/JoYLfXeXVM2I6VtzSiZ
8UaL/gAcw8wZSahLj0+Y2ri9iHJzy/oEr6wHDY3b1W+IaNK3QI7EHnsx1ecB4DihpyqyoJIaADg7
w/pyNwlKnLdFA2efRHogisl/2M0cFMDzP+B7Bv0uD6yIAcTnAhsAQfWtApxVsoGOXx313oWBkFc4
a++Mp5DDYRDFyxeNz6/Ce417gyRNK2UkeE2xRTZbb3V1KmJopVgOOF4TmGneeSvGjijXdEAVEehT
FR0J5Xpf9+dcXgMXasbsQ/1eoyoPZbCtpuX1j1BWpVz6owlh7GrCscYHUY+IE0ZkWo8Nxp4oCeVX
y2fjmIjUdZyQSkYdDuFKcRPMKvASta5vmwZvmWRdyngsCsbMM4B5xlDRDqwNk7gmgkX3tlxOAwLV
jhUI+kG7ViCycTe0brLLOWGDALhQOOG869F6pcpDXnDoed7Y//yvMX4eh0QkZ5If5fUIkWJnvxo7
/g3ZaHZf4S+wtityArA2FP5sBpHnprXkYbsrIB2cCbxsZDTf9ksn0xuhs/d4XARRsg9Yt5T5yJ4h
7M3kxFXKfYfTCthRxT5iqPWvWHX931ZMt5KNN4K9IqAUrlOxN+plQqQrp8aCqTFBu3zx9m0luMYN
mh4v42qvvmwNFx9L1LGk3pe6nDwOWTQPeYZUPo2pZjl/SgQ0uQRf2f8kodQYDmPbfQ08dkYzUULO
G2U816c3j+egWgXhEKz8feLEnGch/yebD8R/yvO//ilIVbk9egzfpfOiwMoxsdTd474QydFYFKfk
YMbcqJxuYKl7ZoReg8R5MwEoFLUbI95t3ubOYaA+EMqfxs0aACsU06EqHOrqoiyobQYlgwP9qNAm
9Q09D3PdlkvMqaC3cHaqvuWlZEVqEpdE+IJeMoBSVvhRcsrzpRTC+FiBFOFKsRQTgfFnQE/GLy+I
F018+qM6GDmFomB/iZD4i+vfFYQwTsRoZsEy2Vz27phhHtbdkmHMAZTgkLvHhmTZfQGrIGAj837x
lZ3ej/MCgXFJ80LvAGbyb+5whZFAGsXRvcTudymnlBDMGyjRxrFV1vT9czMqYHojQjwRuxox3/EF
ylf6nC9LZ8zPfaq+FHgbSJqIyKK3dntdFcEyNABJi7s4R0qsa9fUW40GRPg0vykYdiKysP34VNOt
Xf0jDd951oAWIVC4g3wnx1Bw++RvGGf1KnsBjB5q841xRtzWu5Gw05itOerfBN3im8wpf9t9j+k6
Z75HLY+ioJUvJFPWgM8Jk8XIfOCyDxj5S5mzquISrLQdLkcHhQZNViNWMWSmwN4cKSRLkIU7PjLV
VRo1IwV1GNENGQ05bHS5ALdfYWJmk4iTxFEJUDvggwQk91GREYNEcvrRHWnMDen56zZGD0Eg1AfT
ZR+elXCprkIJulVIWPHhWXLRwX+DH1AurDXZ5Jb71RkblSxx5ejEunFioFK8UZAV9ZRveBcb1/TQ
D4Axrd6PkqVNGHOF3OUxRVHbTgbLglpgymkGZwxD2nYFNsPVFkc3Vcbagi5ejFa02o/odC42Efei
ASeKz8FCNChHL10LTfcWRI/4TSWXyFESaXsYmucHeMcPT1B3PYJVIlHL+tVjAF1Fgcd/UhfOjHMX
rDv0cZf+DfrZ0rb9TXBRt3CA0Znkt8zCwrWGE/ybBzUMxN6BzfH7cTfcjBVe/fkiTKUovtEEv23I
3GjZ1KZ2JqzEWwGm2Foy/pwtIBDz/xJXrGZwwoDk15NIk/5NC30aBtaXLxDDH8oikIvXMUAOXiOy
qSFxIkGGUp3x/8/29v8yAL+SL9heKj4H8vnilNyKYXMFov1l+DiH6DtAUt/LLKxKJjaqwqzJG+1r
oTjzIeQiaVCPDD9Rmj6n+cKY75oyeD67NL7i5So1DDLpw0Uce8sX9za8HLkJznTivRnvaKRWjX8L
oijJ5sF7sqka78V108J552+CtgW9xB8RGS8dm7+ACRAfLVCPBGLKr4xk8J2dJzhFeNB0QKWcd2rs
E4oUZmQHv1GkvamLQzpimN6enIIVl3L60/+Lzl64HR/2Y0k+NI0vorv8oTgOoKOUQE8Y5vLKV9ON
ZfvgumdFiUTafCAABKAijKtsLJZ7fb8cDcBSF7SnGo8RTInq2ibE/ULJ0mPCMiNwkj8VNPsrzuY7
jmqm8bso4yxj1s3aWE8BugER2T1h+oaA3o+lRU079FBF/ZmPTMcAdrJlOJPMjFcLZAfVFPoulxVn
B9P7LxpH5wnvRfPiUWGRH8PshQHnRTz8oJnaV3A2EoFd/9uz7rri/rEeOcBrv11CDCzq3BWd0136
vliUy3CBnCyeZ4CqRyNzRNvmxu5eXjcpvxjeUehbMyY0yDsS7EY8YgP3lNsVd9B1lSKaq+al0Pob
u5brp9OUR5C4MboIvZRZ+a4sx5qLZQyl/6sPiYGZy9W2HyTS9ZuCU+ObcSZfYGbRBAwc//AFDkIK
fU3bnIJ6rwravUX3oGq8fC7//wdn0VBvXHU+qzgvvjjdjbTFkYAJ0MM0ax6QeCYe+5bq6zkaiCae
RjgDEfoDrM8GbrSbEIOv/DUBuTbn8XGo9EF6mCHbk7PVaQUi4shJ/yvGY9Iehlxq9671uW+2OT1h
BIoZzSdI68jz902nix4+FVRzJeje379QMLgWx6Olx5OyKynxNQmdunwYFf5bGhLwwDq3Zey2y+99
4BS2Fae/N1/CmIwKcMfIYuC/g23o1FTmXiNI7uvR8pVYGnxdmOMdYH67YCZZmvOQRHsRK487hk49
vr99Y6TfAfqPffAMY3RBHHT+GQyefx0BjLDr3wFL8JaGJkxYXU2xf13vtQFWuO+onsbnogqOMd6M
FCgFukDBQeA2UEF70RNbcrPr2O5b7fA8SL4o6JvUH++10F1NzxXy30O57QYi9xiy9UvQOg+GhsIk
f6+u+/bLR8FM6nCRQiA9MEMA5TQwqp66MiSWnO7Z7unwrd4bbFqLD0BholrXrdDTEgMi66Hliyod
xR8k6udBixzerFE0IC5hntmPQxEuB55E/TMSrlOCXswkUVcpb37HX/I5lPQxm1Ft6Mfv0XkxiCSp
lRhwvdpmW3iPFEz8/n5NGtRCNHo08er7jXEwgZKWbkgZOZvlNELWhYyW2yPhp9pgyxmhV2/JUdKD
HUW1pFOR0nKZUxbv0fGa/C7n1J65uV1ev6Xo/EHzwUfcnZSTUCkVEVgazxOzgPoE78mleZaUBWoz
tTYq4dqHipVUgGADwpRjtD4Gm2j1qz1zmgCIwvs6XT0cSiWvvDyc8Zr9sSVM2cW0vLL30t7yscII
9CtwygrAgqsQMBGV9yc7umJVZ3qXVItOKL2ZTyeKXXopoHs8SCUnFDXgFNTrj86un00lR/D15/qV
wU7S8oSa3tBIA+goBpiHhs9w7+SiRuJi4ohdgitqaMC1LUBnj/ZLrGFZopxz+UtntxQe1H9d7m/M
6t+tLFH7fJVxg12ljulpS4ujITaRPekdGDDVsPvkaaC7YnyCzS3fCANV8FjF+TANJ8fDbE/6MwjN
z81wN6LiVXKUxPFV5uXjomhlMC5Pq1ZQMNsn72oCpH1Lv/o6rJydfT7sej4EKzpj8zICgqiBvBtm
aLM9gx9vE/4UxKDc/zV8CwZl/GX28VTOApg9q8LT9r1a5FvJq+rQfnsQCFdmVAW8ANXq1q5hxRQH
FixwgE9YKg9B+20BzeSGFRjhY67g4ODncQBuYnTj0T+7EQziweQMRHLTHYFtncJtd7Q3Em6CxnW+
qg2/Ru6dBpwRxtD5pu2v4skWjE0iAJnq0nAoj6SX9pQxQOFoY5wHmr0j0sgZOhel4flaJVGftMC0
OO4UTxRZ9doKgYbWEAab/yuFYh4UbKXHDrqCK9rhEBJKjeNJ5TSnp66fAsq5lQlZHyG7rudC41eK
lHvhf9XtkJOiZVzd3MpeAL9aBglhv6Hl3HRX7jPZ9X36uVkfuwybowyBAttskjACYp22WQ4N8svO
4x2bBNupsO8D2V/BRGyPPs+g6bqPxZOQDfOeDzINuSt84XgmNFTlJSE9QU/96Aj9+n6LcU9Li4OV
HB8w4tVOgx3rcpXj6dIPaAZmO6xqoyH8Qx3nWWU0L0MQ82D+U3MUKSFK23hHSzH2gwJ0Q+u92SzN
vRuKX9kOrdXeKUvsdp2tM8cT4sRvM3FdH+A0nhXd4B0aqQw9c1yvm8NIjd7eIyjri2g7Vgg2LwS5
syAm8ETHtuR4R47Q4NwXpaKYpCSReTFDwbdDIKfgmZWvN+Us2lHgVueH943cLPRtUN8RLBFeSmwP
8R7vLmhIg+VHTpMKJBkzWiV1UPBYvTMK9vim3AboTYDA04Tch8aX/VRV0wuNL3ezTr9t5xSB32j6
iGpe1G9vkONPmwH7GVpzi4ZSEgAxCRqB3NuzKr5cT8fBLdtA4aDFSqYWAIsghyKV/rkgcmXhjV3Y
lRnV9F1sHmqgnWnpmETWfRdTijoSH0pA89GD3mpibhAzQq2/04+QUX6x4+a8SAsbYpia2Z+jtB04
YtAY8oVM8+tzzRsnslNcZwk84pf7MUcl9NlM/0pYI5oDZn0rVVSOcKxVpVwfFNAlZLZiXpbo9993
MD9JkNmiqnw9BDRYpmNx37jiFxaREtPws7I/JX7hxyKp+jFCGDR/kKYB/HEyxu0USMscCUM173DP
cD/wju7WbByOgPKcMrJ6QSJPdviegT9p3u14qBOK4JJo63yhzMrUomahqH1La582vSA0Kr1vpedO
h6TpVNUyCwQTW0+FO2vsbIPshtm/ATR4TwrTsajiTLuCibydjgPMzq3n7ps6YTXcOVcEUSgvfZN+
VceADEiF02V5bkf+oOZKQcc7iUEypL5BtNzlexyCUbnO+QIOnCWrecf0OPGxfyaGHPX5NfTVhn9J
1kA+gsV4PKTspw7YZhVRlrO9Ua4U0w9YsXQf7r7mHI9QxRSY1pVFMI1ViXb3sNiSQFLP9N+FbPsj
Qa+5JmHtxTYWJ57BBVeQaeDVKnTh4UCJqJTU6bgMrYvM8B4TqFjZrynDXT463uL6VVh+CWw/o1NP
saWnxamPk0HXlm3LWQ0eHbY5rhxM7rDRNoiSB4jwQdYGTPRwzVnhcMuX2WuKYBElgEcxocg4KK4s
Nv8XHzpgMzgFKn+rYbCB/CtYp0hg+FAmP3iP75fcm2mr4uyAH9Wejaesm79n748VrliIOlDAQ/F+
n+ecpW9O3Yw1uNexSWhlHhMMMasacY9iy+xilamOGKLDxo9mGJ6zKL2IeuPUfbB38oFwYHtG654p
0qEOrKHlqu6LO0nYe1aYu/UDk0znDvxM2vp78x/lXs6TMlVhg15jWS++DntvcFD1xFwzm23MtL56
EIOqmFbzO/8LHJxMOSWYI8ZalHBj99UQNH6suxWhi/CS56NRvLNNLpjPsBnnvybUfZTQHA+hKUo3
U9kuRmnSkUE39k2+lZG4lBchmkm3qsxgF1GKgy3GG2u7TGTZePO3WnTMKZi7wW9OlrTBmq2PmMBD
NmLmpsSqpsu+2s6HZqbHqI+ftzvO14kLIf4hRILiUC9eS7/+W0d2RukyzjPwbmkh7d/qxPpDoUFy
YGneh1WKrze5+b6BtxOHdcVSkwZRUQ22JuhRatUjiKcqAFjG8Waiy5kPkCvlTnsV0+rmthwAtzGG
8rqgEZEwtl2znlGtGHOuGocf+6fCzR1FMzUCCFasThaAsS2bt3rUGQo5sZlBm61WtNCohdayoEfs
fTzmtDK2k0w9wdHn8FQkkZlBbvy9ECsPAgS2A5JI4sbM6IV3IWnAw2bsCdczKlbqhLZIFO2IKMDG
XAV0fTptokaIWWqDxbKaf7dVFWNLnYJJYlz5E0qouON4cJF9o4Uup0wf5j4gEvXUHRro+6mY2gDD
NkYSlv89Oc9w3a2sVCjqQsX+ShJVpgpCFjqbq2As6juWsKgoCuURgfozPT7laVg3/hLY6wUZsvym
+VPFXJaCLDV2KeReOXfvNn2OQGsErRuRMz3KIXTqB5LsXs9qWtq2JlbHQslNu+h+jTLiMDpC5Kaw
9GLLkOkjhqHz0f3d1CgicEcJ+ezj9NFlaD33KZ6szbhqMJgg2pAQn8szD6xQqEkU4vgwtuNAjJZ3
7enPZaf+W0Kv7D7wSEyNiDN7zG32SyOj5e0XqYWJiO5wfO7t9FM47wzWfIQa8JMoozOBotC8CaTc
5dVmLxfD7JGJUGzkhjUZOjNVP0+rDdvtv0CXCv55+Ifa2jNfPosDAH+Y1bWOwrc6PRXnd693Jdob
0A5yYFZdiUoEuACNgzSg+pHJ0c1xqItBjEyWr/n31XmPwwhkvSMzHpR8TEo9tNlT7BnBI6CPMhbV
DqOdnZ7Pjj4b3kvsfannp5nh9Uf5ibT7cyhCaMguiWAuHSJa3tcQm9FTq0cc81xpUOyfA5jSy5dl
u8XTkgM2RwmO4FgCNPzMGtmb/5S64n/Sc6VyMxcRcwS37oEpEuMFxKSW6CaPAy6AC6zuz+KNuach
2wdzrPCDcJM0g6Qt/h5RidfHBR3RSH+wiB0o9fw3CVhTYX52qjDfDjEEdT8cEVl4YytQZB7BmLxp
GRnKFSCZ7y3+ymWfXCKMhL00txSBkvojztjdqhDWXfbhAxUAmO4chCSS+yHnnaEyrIGJ5ShDWt68
AhE0DBQLHrTZ5QAdCE9mxZXIRiadPZEZ7+U+z/9yMcwh/llHptiB3hAG0nEto07lmFeGoPqnxNsj
qYwzNHjmSZbK8yx3lhTgX5GjmRQUjzyxiBbvItIDl2SAqw2mrQldO06RKpswFyQCEcvjsz+VT1KW
/1uFQDf4khMqvdhzNj8flJ240NgdMwUlaVjrXb9HIZYxC0ICkc4fV7sfXD7b8AlqTDanuW4LhdLH
d7wsDsxPyTFXE/xGVg5KaaZaoxoN6x7ytg4LBTNaXxy93aQupuj+5TUCqgU1dUe1TmoJHrpNT6XJ
nciF2xyPrQ+lEpwzDA5Tn0Kqhmtqaq5w9mrrsueaZMmF1FfC/8RlLT8xQqfBAP1e+L78PNSVy+PA
Dq+Y/r+BwnRRt+mX7A7s1PclN6LCDwr+Vbbt65yzIdyPYOKtRV+vsHVA2LCG9X3hIEIpzF1G3rVS
1W4AuxFAAh2apQvfN4zu/RCbLoBRQin8DW2SYWM3A25VGxkEXKsteTdBX5PANi5BJeZx/ExEJRt2
qbjezyzHgpA9YFrRHW8LWHopFxdMcTHFepMkxmEyqK2BxFBgliqOpwuZqlXCRAuN3L1HFwegJy30
h2dqEYNQfWxqSk9uojXepI9teWzW0x6hCqphBa1a21qrnYvP6N5/l4EVS0pxXiwDI7xCAAKysdYq
FIemoz5hVV9Hg1MbUE++7WaD3BnsH81mJOLMRuOgaR7n0qcBWzvg5PRE6EhOMkG476kPeUtkogA7
FOMZEdTKNWf1/vWTkp/tK+0CU1chORCWfYeBPq4RDom+FjdNW1jtkvs6LNuYc7Wh6yyf0LNjNHtW
qE3gelWextmW8TLcmpwHOr5GxBP9ZOUEaspwa0bEMO6cJgWHITDdZJFIFe4f9LAXO/l7vCgeGmim
/yqSdfwNu4pxcpTTZ5/Qwpy4SL+1qrBf/L2s6Lj/L1JPk77WOYscIRkkMOLEWq+uZjGH+no84DhS
oVk21rAt3Azcu3+mhA1ntu8d5erNZtbnL+ODduETPOF7UjG6cY27vEpy77PWuEqb8h2xiGbdwnwj
SRDQ8aaExOJvYdm3uyLiKS72O87+pnZmzLEhl/OhGXbANV37J0Vwf+f+eUnFeu9RTkp1w0F/pwo7
UW9cRfQsmjx6yawbUu9lDDRNVeP8C1T1SB0kAQrKBiN8DlPXshcijYtNWhfYSTf0rVF1GGaPNjdP
yMJ7EZBQEfi7HxiyM4iFL0Yti3SSmzaK37WqS8/+o0IcE5UIM7kJsEPu53usmwzAfoTkpmZtHvhQ
g6NpSst1NY0qgFqJk3fxyaGkDHBzxEJ5AEiM/GsQ/1iRueA4CgT+1YmxyY22B6MB66JjZ/n2dYF/
ynWgh7D+gQVQzS7TSlyBQ7fRov5niD6rCWI+We+wKR7uTrPE2uUMyrsp3TthEZV7FsTHMoEDRi2m
xzyoAykg0URnrzrRlX1fs8muJZ1EXUbk3rruDMXERGQBCWvTby4e9MZYB/+a00HtT4puXLzEvcJH
8Zn3iIC+4a79RojdtyfgNZloAYJ6jEsdTYYjARD84J1D/4I3px/22CCbEmedae6UHbjUQlECsxtR
2cEyEWG/WWW090v8FaX9AhpxJ4VKx32e1QJY7m1+6ZPscLBZH0iB/sfxe81LjEox5BmlfV6Cb5is
zaVTnbBETq8u851Bdmpu4QorS19gU1QJgSCuc7YDC/DEdUqKxiikZKJaZ4CfMCxXXooUP8pZnRiR
s9U1tYY3BnkcpZXhGFhbpSuRRCOE9Tfs/jCTaTT95cJIV9aH6i7i/Ge3XfprmzIP8RlQXXDrdBoe
phgNRiT2ChpsHRKNi73R8uhp1j2HC47cBm/GTT4MDad0XTMTPdnipssXlGivEXlXbJG4tmH8i/DP
Jgs4Glx8Ime60y8tSp4mtpJCP9Js3YjKHufPrcxho3IFpm4HSf+CDkDNmxXsE+Ex/2aSr0UPnpc5
s9A9ZhTRRv5gOkTy5EsBZrqIfCpnVHC/olC/p1n3yGHFLUUe79ZVvmSj+ZtL/zsm3uduTxjyVuBu
XP8VPIez9jQOG4FN/QtwZJCz6oxFlbaHs4xz237PmWn+FR2Nw3GkPiT/yeDOxobbRZLada+HDRkl
lNsbwC6lL7+g/Za/MEZ2vawCHJBYPQps/pCa0rYLMka2PbRejAmyNLM4J5B5VMtrPBC2JKGpHrJ8
pEfrqES22H6DKewDSzghLJd74LT+GHmDk9mU2H3m+uy7Ndo2Zge0OhVx50OfnKXIHIEK0cO7FwO9
Sp5WFzvDsNed7FQWRyEeyBeCPBJKNDMdV73FDbBdFGyCvUyPJ4cGoIMCJMTZ6niiDptQm0Ji64dV
0dCSJz+gtWU93ZRaUI7qq08Pj8Ke7+TPfZrbLXMIgurRvZo/XA0xXY/YwMWXYPc+dzmwSBBzvMDD
2vc8+feuZLnRdVYHcQgMWlteM73XlAI22NiWWVsvLp3XVaOAHhRu9qFECJAvU21cLQN8j5GwYaiX
sAjrfl/fA4Vgsn5AWG5CkPlBluGX5XGm4btHkZEbFc58Hq277cO8HLZfmHS09AWB4pXCf6N+H6Y8
dxRVh3EP9hPnCxSBBFQvAoXccn1yT2WCz8cFuX4bKzmE5m0S/tuTwZSw+y9AfwR1yUgGBKpHG4+R
z2S+PWidElPcGe+wmsVO3/WzCd6nL9Sz2/3J0FJa7Us/oAAsWcstB2q6F8EC90774/E97NvrcR4n
yHuBfSzhj8UPuegfMbiEJpKwpbOFXcOVw9RB74HMStHhKmRadf9CnbIdNCzPRtBuzSsVjJEtpAsG
Hb568zI2w5wdvZaMzwOY4xfAJQgEsZsmPGXwp1sq7Mw941AH+uzK2fZcdn+R3C2L5ux/qrjQVkyV
XIWfn7tj4Rbiq3BuGiW9YG0M4sHWMglP4c8Fc3vt+dhZ2flet5FtcZQNF4Ldu1J6oa/PbGjdVA0O
vFgLC7oSbWDXdNzVI+WPbGHm+FkAd8BZfhH74bfts9COtGXd4ejs50xvrKxoQEZRFOOcbT5Eym+2
0zMreePv0M0neh3FdJCQ1pPO1QuRlDIVwTY54WBPXLyi9aMd312mj+TbWAncV/bqsUpMMhy0NAk1
acpWyuZhW9ixljDL+IK5cMdtdPIS1tgHQwME/KgB3AS3xZ73F68iIOCVWGFQHmfm2n3L9kALleDD
ztDbTm6uuEIzBxLf0v7qkdRSrzMb65oeczWYaNnsZMd9Y0ILNwXrHb2TBeBpyWHKki8vvTg/sGa+
cwsevFAdDxYrwJT5UpLb1Wf0u8K3FdCG724Hnlv5WEGeuXAjNIkZp/xlTEXIxudhT4KjXtvvIcjq
UZLv+qnwj2VpPgayAsditkOdoQK89ixaaT7rebh41KWzZWECLbqMuzcBH8s5jFnLFpzy/+p/qRPv
CCmEk+3p3LAqBhgE7HsCMKMxIoVLKO2s9s7APFtQBOVgUO8B0sHpH9qQ5ui67aaFGAz6K5VKOn91
umPC7ettxk/SXTGP7+9lgHhwG5c1McyK79+LgNkxrYdrJuRr3Xly40wKmBJ9Yloisju8kxn6KwLZ
8/AN89GMH5xV8vnMBxi/CvvEv/ENJNLkG6Jrg1YMtBJ3kuqX02tArniHJrr9ptOw1/VHWWeHNlaK
ELjOJFNE4IaGicNVUbTseBso/l4DwAEsh7LcX7N/8B2SXizGmFMm/wigRwmLMfUh2muLZzBt6Tpa
8MUGR9WK8UyLsWFp5G51TrpTvcZa4CUjme6PKu0r8u8yvgQrf0skUbyFcCCdUn3q9RDbCN9bPLUH
et8jyeSbpQTYoZlwAHABtQrxellY6ExpTfsr6UpPxsgeYklcIUdowyqbZ3hOzMndjYs9c1dazcJW
hHPoeGLWXixyjs5ps31njWggQolTFOySct9Npduhxh2zIrDr9/0jIfyBnlI0zGLwz31jDC2EiT6p
tGP9sTAnZQA42FSIZa/JMuorP0apCzgDSJhrNA/+/AoRhbLyaDAuGYFOSzqlTAMTKe9dXLtZ0GC6
lmtvx5+g1OBm0+m7xlK7DVhi1cme+/Dv5dyQRUzNRJtUGsIltNuuBuarAHnJDef3fgudPVYfjHXw
TJyDBl6G3y8BSoU8JI/jsPxtjhcuHDpFrGcYBdyp7xYJzNlQhVVZnE3+uFNag0qI3nn18+iyc2iV
1nejaww15XugZ5vfp0rAAk4tG5vyv9PENF3JkorjHlXFh7K0eJD0rav7ayo+zx4S44IXe8BxG7W5
mlw1wnZus70qFC6xNG6cFxe8pyDiwFJ0kzrohZ11FwHtPnmpDDc3fF/ua8rorUPJJ4QvwZzgtDq+
oomW9S48+/bl8fXZ5fF1YD3Tyb50Wl/fCldwL6lxD9UMn75E5XcMGetYF7uS8oi/zcSa8vDU6qxX
A547zCoEVvl1LYzSlIXkKVsil/H9DYbKNUobMJUVqFGU7HHVUYCE7qVQuoleJjZYluEvdHFovg8y
GxrizvseZWZDyJA6gRgh6SEguax1rr4wIZennwo1sRZzs/W+PYvXJ7XDcR7YYplNvYkrXjxGs23k
nG9SlRuWI01iVyuUyCwrfUrQxyV52wZN3TM24HJyARBMbdFYv4h08D34o0Uu00UnHaJ54tobsoRQ
kDnlONZT3B4mc81eYnA3VgYzZWV8b8+RN22kSGJep04vcbzsClvtBh2Q/MFvU0eumSCOq+Tnq653
jWro7NQJNazUaCyhjdu3mFT7ZIvpYhJXTo5mQ0OV384xvlcpXbzeXnMUNTqu1rlPvVfhfSz0T3FY
vXkEuqWYvPEUqI1HpeK/qxc7UURLilKlNmagUL+i6/+gCCZiQBDDmIODlyJDrN8qA1rSZiLBP+a7
BrKvwj7zQB3zCgpL2gtNG3c1taVG4CKqoYagBKwyyvLHjevH4vxcAwOm9InT9AFdO9q7N9fj6jx7
jcQD8siTbDcc7sZMuKwSi0dFxvr5sgYEqXlLQGPxuLqzKTl0ksvtw8Qx1POejC1htVSR/bS2X940
+OylYq/RTGkCfp1P5hkMlPZc93aD1U0l3LyArS3mKuOp9q8GeH1lEyMk9g3MKhXqxzwpaEW6+PVy
+mfc0JuHQINv7Ww8e71k1B2e3dgfQ5rLjgr0LqSjCS18+BdfD/ZBUbpKIGpgZN79QBg98Cg4eG++
FOwfw+IGFRC0DRqzkypMS0yN0o2fVI7uEcmGuOCDqY50CXm3fCcltyYY5CS6gJDIi8eL5CAFOcsx
zW1w+2jt8vRK9csUuYvwzmonfCOZ6TL/zQ/fh3ee8CdvU4HtdHuo/mYSnd2gPJYWezrgGVn6VDsW
0lVeXdZAF/6apkp4DlLaXAg6VOF8ZzVck+ZMPcN7O3LmkXHi9VFEv+nuzUWrughi72ennJ6QyO3W
3WNL68gkWizv5SmNfC30PB7DsAUoZo+a16Z3Jkwn9wqHWTkecQzgjUbboUJaR3oXatFdBPNn9Z82
TIUJHpkwTA7hdD6z9pv4BRIHjHwaCEWi+wxrTy1rF6giVB+zInGt1p57M/xsdQVbLy7wN3l+PCL5
KQlVCScLKVVmeae4Y96RWA+2uSuq4F67nA8dVpp2dORtDqi4rW/w9iEWBmwc1hOpEzBRvvED9Z2l
juqjkyfiP/HgpGsbOpjXMLmOy9xdgTgmlQlWDxp+CIIuRgky1l4D9LlW6qnK10qlBzwya2bhshhv
a5vs2RXvK81/YtRdRaapsQnB44FumTETcej/J72I9YhZwVagJhpoeN8KUL2OaKnTWdQSNPP5ur1u
PJwCZT6EiYdEK9EtzCqFigcktKPi0rcVYBA9u662vAuHMgRSLc2ZUrbSMUQ1Q1FI5o7rIlYmVnNY
ep7tcys+CIZOXf/24QrX7MW8gppEhBYA9BGNiQgQar8MXd5Cea6qXnpU11vAe7yS53dpbcutw8jV
SUu/TzzFFZDcT44xdx5RBv/x3nKJ3tRg2EqdGqxrIe/7KFkp5f0bg94E+CAtaAdhZ4w04EbtFfD+
azOZSVffJYPDbT2kh+oxY+6OI31r5jQmniHVb7ZlxHrOLS91M9cZr5L4iv1G3SolMqEurEItjQWc
jdZuY4uFqMTHFLkqVfY1amUpKmgHYNRWrFUPI9dKllfgHBuxj+7bAc6z8ECaOQtyroa+zuLw7/5u
QbpF/UMKnor3A40jZq8EFrfGTTX+p/FYK0OAYd8ZO50gh4QISBV3WD/JFx/nguGtW/EMgOt08x3P
WvBo6DFpFoYDBt2Aggb4MB5qDQ5ICuUj7G5g640fZYaK5h9G6cWWsV0Uy65dCKkRdy+nTwp02gDh
sTucb6/e0taqvqxgxz+koPyamCkjKWi7OvXN7q7PB8WbDA3YsqqXOTR8X7fB+SrASW5ty8FscchF
cASGDLgALJuleRjz2kPLmtypaPLB6x3AkyWxYTcHZJYUb8hCVAATps6cTA6W0+julVKRGhtdzLgJ
JRXnEZxjsKRdtksskfQydnzPAKXV8skur2cGv/UQhGoylTYBzrBpG4X2vxIHH3kEDSVuyXpqVip3
MSAedkTOXoFEemrJn+K4bF8gYYxCJJ0OmPotnG9asi/PskDGXRBaGVvtymD8x3OPqvaa6winTTqH
Zz4iqWgEGA6xTrzES8ARz6Sp3BoSx18BOO089s89kbuPShckqxEY+wHQD17A152X/BMMfWtm82Xu
nm5oJIolYSNLysGEYQq2nr+btsU40nLCeLTkAgZvZBI6zuaHZtKmgw0vK10x0du2vUddMOo2NaLY
+/3rFnsv1PXOFqkfdM+YnY5mzXAnGw7Uo1zEQ7HLPnVRue8LjYevxU8ghEzzQVNDmHsFB+HtVqeW
TfooTEXIkM3OeqWjKfM3kWpVlruhthmxNGIQk2twz6E9OT/e6isXsQKBlZydoGMTkIzKIXbyruuv
1YUM3eu+h+mNm3ivau3KaucXHCr80Sw23EMDrmqBWsLexreP1jcIA0j3uIizgGBRR+QTFnG74CMm
5jRDpE82HwBTZLA+kX/3OgCnL55X936QXWvU42Xs0255gKD8T/94HfT+ziKsN0OWRVItNSgOkY9U
KfLl7S9EM33tTVgwSCZogHLGPgqCE+tBBuNiBK6f6GcJZG2WCQjEV/Rin7seZ+4VEg6pSEJKy4x9
gI3YV9IGmbGeH7PchvTFkA42Wl3Nmui8TVuYnYKQCnVBZyIqqClgKX2rXAWPGBwy2pBtIsogZZu1
ybeBtcNNI9N4BgiKAo9EdP7y2ZEvAr4nCsBesYyy7dl6PE0/A8yBTp8Msn04YSrFaV4yIAFmFteI
DR70JN2497UOaCQgCtsl/STapFiI+Y+squISMw9FpYFIRuWRufaXRg1Vt8Gwk/bYT/C95/Cu2GE5
hqsP14+jrUWxeIsOfch1v7I8/3IuHuct56I3VakMJ5q0ZuvuBcpn9OXHPi8JY0xXpDUJRpNBCdKS
HO/jJMGlcuNsTXcaL4+vFfB/YQLfU4GJbBQFZxRGdWhDxLE7MckxfkFwHs1iL440Ehimj3mk9vGn
jxdNl98c8FCldXYzlSodc551MF9MmtJ04tPaH9CfMTEXmSai/JWtS5QBv+n5d8X4qa6VaNRZilYB
UBSAzOYSd1MdeG6SyO45KaUl3yFqtI2nUb7PtTrGAipXawhPoqzbjY7+VpcajH8Lq0yH93gmJz6V
CHz87puJALXouRp9XMeU2l6vDSyShT1R6x6xZ8Y1eA//uPARlyxjnSAhoCsi3Ejg4bzu+QdXlFtB
211+LjyWZ5liu8/yMpPChtVWMTQE3l0Si3IBdgfumApH+sV6DHKCjSWrDa+iGvsriG7O1UzcgDkT
y6otN4OsuV+mF+MUsUEq+7T2EdcR04gQSsZgr6mSXG4Hi3PlFaF+QryW4JUYFzJ86XC3ekKGqmcd
Tb+oxRCAJsMsmJAVwg6xQ8R5n23ntnw5BZAH1kLeDaH/nK3h7OraCFVfPOUC3iiIYsr1cEiyLNUR
wI6z2cWMVC226xxsvSfZkSI+c5vnG99mGbfMt6Nye4MjPCCmL1sMY9Xhy7Ps2R/WmrzYGrp+i/GY
htxaVI27NsNryR7dlctoD4kT2w3sSSYX/9vsvYW82qLE8h8ART8PL0PHWJIC7Lz6UIJNjCLaQJOu
hv/2wVyz18xUIF0AO0XL9E4YlksNXstxAUa9UliVnXqL75nTdE2ZbkxtVCTGBIjdQZYA22silabl
Gp/sT5+oebNPACDd42jVwEyPg/oqxu8IdmAhwJauDwzILuuuQYOTKM4bqiquMa6uJlL5xRJbeWWV
ErMgH1VnSh4ge4OY21b5JH/imEIqbY5sOb1pDQs7BdgPS1dYbxcgSs3koOWzKnbRQ4diJug8GBPg
uvR6JenIuFKl0U6+I7XvanePygqfwnAhqrsV1NLzCCRFtBAzf08upyQi11QWI+HQcoZJzw1FSXHU
36V/pEqqC+AvjntIi31QUdSOh1ztPFMBeXugx6yua1wQiy0M9HYF6uWiRgCfFA9e1ba2OYXh3wco
Ndz4LjA2sCZtzQzklZ/IUMhif2RAsf0t/1616ZE9HPes1vH1eFsbkLF8cooNW9Env7mfLBmmV7jN
oAkWt4+rIivNETrxBzLnvDuOGGAtSFCLnaWeWiNmnYXTF4qgmWHVyK2z1V70PKwfgjlyoPf3JzW/
TadwXsdu1164zL+qR4ZkUq004blTHQS6Ywc15Nnr2126XOHs3U6njqlmxCwi9nVeuKrpHxxsMxaI
kmvJvkGtGNwb3LEh1utDuedejORQ10mAlC7FQ0pCpIy512OSy1fJDkqqL9m0acN0ZteRVDMXfFul
ToStB3w+sXBCUnUiAmYZaEo8UUMip374/bF56jDimI0t/ErLyhyGwpyB1O4n5hH2XX+Twq+fy1O0
/hRMFz4v6t3LoP2iOjFAaLgTvsva5dgwr58C0JDLRajyjbfXqKDnG6+rxHPsMI7PTdFsYftVqTcn
NOmLJjCARCy2NJX//GxM88uEWr9eLWNknC9s6Kwk2LKP1EWnQEaRRD/dTajJncZgLgkG4p4kWtoA
N3uf1YcRb0Ez77kED+HinnHN4Fq0pPSc200TgdUAwGn97ZjETlcXTk/RElyQRa3DQRuYuiwSd/Fy
H5bSCZ6odQBmdCRP7TjzHxOLQDLJMLuOpcU1PjXj2iQXy0MZKocpaxA6lDZBq22RZijDghClHCta
IVZ59st+RKB4j8Er45ao6n8gnLD0FUuxcSu828Wh01Dolc6gPhhivjZbhR/qsjx3glVycads5KII
8xMouhXvxpnClZcpJ6PrKiu2nm4Lhqmk8rda+3SJ5ZDNhzRb9mLDMNV2EfB/L21bAIt8Bxosucb7
pH34yUyfMDjZfIgkjiOaixg3n6clZfMY5ckbIA62DjfAs0ak8m04lMPFFExA0US8pTAeUIL6vrgL
EWObKYI1kR/YweXaQ0ram7i9zEIQtJQmoBtuxmSR4GYWFKCPtTMVTmX3karkd3oD1kEvPpTTl+D3
AFqM90lP+bVqHLi5lK2cYpe3F2vzSNfg0mIewbwAw5+bLa++lRg5+W/B04k/cLkRoDbTAx58kRAB
Nn4xbtcS1CSXIEqdwk3vULIIUqQ9vjuyyUjzUkPR6OwD9dslK9oDA1ltuxR3RgSeW6R5LEQtvuzY
ATxW7Sb7HSlxmqU0hzEkxQtqYptoJl3+RRxZW0k9XNX6UgLPAJT0f8FYNSeaymOr+Wa8O3PvL7mp
nWU1ftqDJZgHF3CwCM3nXTwRTHK0GiFKxXsiOP5NAPpfh4er9Z1Y8kHXrt5jCPYMvlk8TwJn9nnu
ALmaPai596XfkS+BQuz6Xmaua6AiKLHsG6CYtbL5OqL1PJvH67jDdWGdA+J6AIhyP2K7BtyQF46r
43vqnblXdVnYtbC2YPYLp/4Khqwhy6gpm6DUKFq9ZnuOr9md0Re3ncnqaNjhUaHpsZwZUky2RSMR
VlyQ1/FCtVUzqinwpf5qKxMEWVBUA3by+7ZG2LtFWn8U3A3dKIK+0xgv0uf2P5/mR04qH6aFvKz+
t7iRmBiIurHId8//aiiymjD43SUX0GjnQXD/yioLoL0Du8JNwj91TADZd0dS8l/QLd3fZKU3cZZX
hVC4w/gjXlPcS8FIBeFCpJRl06r6Ah1tlGgclBONdjymJ+u2FYlQfisEYkrPsFFsjWKYs1Kt3EaA
f0Naeco8P9TWGKFIZuODu2iOauZh26HNWOrkMMQCl2tQtVrVuiYtY45FACDf8EUXUiSHVDci2oQa
3P1FzxkIj4hFnbWJXo9ksmzRoDg9UOy0nKLzi1GbKD3viYiva81aryWyUOuqLWG9BCmaO2w7hF8s
MAWLToajuFPFeXUJdWamjFga4oYP0vXg3o7KTs+4FORmJIpCdTo0/R8wsyYvtBZZOcL24j7JO3xs
oDuUnIrqbniIS4gVCno4GQlj56c97B/CLw7mNTPPKAGCmMOYuXzigSkSycYaY4yjHeqC1XkgkU8z
vD7A5E3357B89J0gEyo4eKuoSfdZ5YY4PeBjvZA6CYRzsvvvPbQwh6+QWnnQjvBFtfATKVKpD0ZG
FPkhOyduwOE9eUiMGX4h1VQDQ/OLO6P+3zdCOSOA6MQo8ISf1X8LL48EYIbOnTtS8CeYKKRQG9io
vMw774eOK7LVVJ5qGOK+5Em1h+pkroGgJWIc9sezFoyLL8TRBRPI/4Izhuxm+ZnMqlKM0UQ7/m4S
/oOuHEC/HuONOOFWRvRzZ9w9Sm2SaYH9yLfLWwBTA0tDSxUJYYqMStc0HG9V4e4oXVf35xmGZFhK
ow0wHdS69vSES4ofHyTt0EuAN0TL+ijuRomTIGdw0HfLmv36W6P6ToDRRxK8W903eKIT6j/gmeu5
ouCOavs7hXaYvGvEf2ekbKyAsg+Um2IprtZYEqQGBka7wzXWMEG6IyvmSzJ4nD3M0s1AnL2KCENf
hBLuOeOdalUMf+fCJWRKVuejkHfeENWDkVQSzJjLs23zkMg9P/u/HNiZn0xyvP/RzWMgLvJYyc9H
5yum5oBK3cDAzVP6idkEtPx0LE54XSto4pPzYIiiqDijTsI/oDqaihZb+k3kWqpnC1+q4NOxRp/q
rg971sxoEoABtaniRY+6wkiWYjtLmFHhYzXWvLFP9z+fOc2ABa9sToxCyWgbjR6H27/uNrlnqsXV
i9V94wv+yCKMt3cA+DvYTRqYIux20ShijeOYOdNTKPAnWvRxMiAmnr84Bhi2disuKIzbquD8I9qL
wU8fusM3j1ujB/lD3gtjQsFnVqIPCtKRPHe8SKGQwHuQvG0QcNCCyuIJTEBkPRZYYfeOWt9IaNuk
86pV75zhjqHLtdohqQYGg9SwFltRcozqv7HlCEfCIGX4S6I8rbWUq+kCB459kRlYoszf40t+xpP+
QY41ppSlQTcyq1YM4Z9ajQimU1iV+RAFHbYBkPb1zJ/flCMwnCNg6Kbo7GddoPwCTDLkhiN53RS+
2GqrF+rySwpG1JYrdjMrku3eix3d65wKSrgCIC71cC4aPmTX3fOjKFoEGwTwMhAYmSpBBFMg7WBs
ADBNGuSXrx/FZ0tg/626B1RDstxMh3Z1QOM1GECJZIRZxo/Fpmhb/7yY9TDc/b+NYvC+QLbhiFop
9gOp5838bB4taztg1tZbF2JXi7RAkFH1yb6T/GQrAvY8qeF8u79y52CGtvi8WfgLb8O+taIj4L40
0WXhcpp+WhD+Xn/n9LljToVQ4eplVHm/TLiYc9Y9TorhO8bz9mbmlW80ckiLcuTj9hKhFD+ZsWjI
nOpTXTGhOXOaEQGtTthzeVhowFtFofVCyMcOsG7rfxeMBYH6ZSUL0WLlB0P0uMTbIK+HolyLoBBv
lG7JrSkYGkaqwNEDNHjXNwxKRPfXr6LwCN5T1/bmlc7j1KBp9bQVznp2rRAy5DWJjuFC8HPbQ2xs
kwdVJovxpiA3feCc9dF44nam2uj08Ish6EB/IPuc2+am6T2Juo9W9hBRRG0iRq3GKVYy+I/udwFl
2q8mL00HzfVYZ/9O0AEyJ6J6WeNRa/bE1wnFZwpO5PI5sXiMqBFl9DMu1SnotxrcUFvivAAhebcQ
hpErrdIJp7kbkyZiOyCGTQ8Fipu6TOhkoqHBGPo4yOQSAvE6dNIaxajYTd1cPxi6Mloll82BS5El
saAiZ2EXgzXX0+M83XnkW/OqHrDi4MaVwuIqI9fJrOUgmqegznilN1QLXXwYCapcMHghDF1WgpKn
OIqWFZW2wV7qddTlvLR1VzU7RJ1WVWUhWhp2KddctbuoOgpuRzRTWmQoh7T/WQzH6lYQPjcK2yrm
Atk9B/xoLhNRUPKaIkhfLWGTwCoXdcOYfp4FY58gI9lCFZisI/zsYtdhHtuyueNtwlUQVaQfBcYg
rlvihhgmF3Sm3W2uUAADTL5zY/Yk0TrJP7NV7EZllzvDk3w+IPzEsXEelhS5UnYgbzTpHRoR+z8v
Wc0mprYZ1DHde9dhRmnaxkf0U2yG2YmyJF7lNzeosmN6Eml7mOAvS/LDBGQb/PKRhfSfScG3aDcX
x6R+e+IJa3aCFKEg/CX8/FoGUAwMHYaADH6MEGNTttx/6XJMeViwcvZzKG5e+h+70fH2Gyb/d9Xl
qDCXswnUcs8sGI8h+kvXIEyhPmS3SWbTzW9sPyIXOeL3/dUGw+m74ZfvSXrhOMa0kRCIgvbIrzA/
beS3gAJ3X4vJTd8FZlnhpARAjSmsFldWRstpLD0ZERbnM2NmGQGwgBwjvqPAkn3HEWAXoIa1/HtC
6igo/jkYQWbiqLE/h0SvfHuQ3PDqx2lYcS+hwbbsziFl+tLUW0CrRtjMBg+jZknRG/D90QkrrXrT
K4Fz+bqoY7/XXoZMM+RfVXeXKVyMOlKDpDCvHQ6aCx1e2JmAgEdZGp818fA+eBwgXVulypwXAUu3
97mEGgEqRX4WHLwwuBWBuelYhy8Jg7ZFFhKA0TmMMznXtV6whVIcD4wG7qq7L1ofXyhRsbr69mnr
NKu0CIqOwMXIssIfosfFlNgpKz8YqfBlCcdcPm3doGHSEwwuwIqBlfVFisxElHt5sEalbK4F3OH6
aTp6r6vr1ENLOCCd+z9FOKkfNdFt6AyIEVa1MRlyYAxuaFFsWld2vFbqCzgrKVn7jRs7FolEr6UG
vc/hRM0l3NjGovF8ULBOkAe7R/G14j5BZe6F0mJz0kz/1d2xU1E3F4TgxB88Fv9fpOEAcpvqeBis
ecTfnXoJJh9UIeGmQxYphN74sM86MazmPc7VKQTCD8qePwtWPTmSDYKl/8jor1eY1zWB2VMnIqMO
SIPHT6UKGqbG3gj4ON9VRSkA3Qv1+goera/pz0Kexx+3ijiKAfvw0SJkPg7ycu4QDqgErYpeaZsr
mGt33Vxe4x6YBVRRvvD4NGHGjq4ah89tF31y9do8wML6r5ffEjGFlMej0O878SSfay3PXUOyAfKl
Sl/ndnvLwlSYizl6kH7dG5Q20ecTznSnx23oQwsg3jTVXEHNP58eqdDC5WXkrKZMYDD3oAFtdmT/
9JzRQmF/n9ldxHBTG7XYSdVGzkpBYyBwTn3t4aEXCMZbFAS3s/l3Q8JvMD7B4PymBNW17W2QwDRD
0CN/YEternDzxEbn3B3INpcMAYUL2qBcyoodC1r5baiz4ucwASz5TZOJBeG7hlbq5SkpdIioVNt7
rhfAIjRwKsiiiTMq1/1U26riXVuMHt7fxpkq8L9UvMiHjMLeKp3MrSzU8Mih1yFWwqHr0f8IXAPW
Ys2d7OwdH5rOj9ypnl/lrzocqP2MwGg1QRHbgIPCFfCbtLCNcgaOlg8XH9rgtgI329UbRwp2HODe
IgzbX12DAg1NzjOtRIBBTlfVyWVUH9QMvmRfRGfnoN1vdVINqBw3IBBZhOqdlf1DZjqTzSF2mhRr
ijxLeN/tESR12seqbh+RwAu8WnOOLSgV/95HBOFtECA1B+mnYNIF/PrdfXnvIYQBw8NM+801ts1Q
SoAmJZsFulyGPDW/Dg6CtWG4wh3At779rcbR/YpSCA/IQX3KP4d/4U/LQ4/Wx47NM+LFa68JLOXN
SJG2KY/jpD4TMr7yswl3K1JURS4STKgA8TMIumf/LwVKxRLRRIBx6NLNDmZS/16zsVUhLfQDTqnm
hX2HhBMASZSjnCtOfub+FtehquA6G5/pd/pCLZXaa1A2kcExQfGM+d6mqx/85wCiE/swXZnpm971
V45UrxXCpxRboivIkTZZ6Kw/MX+ofJsqC+KvBycWcDAnEGVh9SbCcQHj7fNMPTCGHRobGYZzrtiD
c9d0dXvOCZic6U/zT9UdW/8+MC1th2zkFoMV9hLRN3/uPVAaWnlSd2q0vGIyVOS66mg0KdiiUlIZ
RMHl94EoxJDEYcOBniVD7l23VsK5fJeRQOtouQnRELZYr3LN8iN9qA9cvTunjh/FEUZaWXMD93mR
QS6dCgH/p/SVBqRvzCzPOS/akEczPri8cj7KfzF/32yIX66W00O7/NNi+SBFAA3J85RGkgA/krN5
urwHHByidkQBdNoDJsRp+oYMPYMRA1jk5LcQI9bXEoVVyp+Fwe+41umsERO1K1oB5Eird0lPcfJy
YAm/0550FIXzsaJk6FOOwVb60U1Pcq75CQN2uRT0C7ZDr7oS1TjLGQH0HuY4s4yFvv+HmnMfVTAu
e60hE/PTvO/y7lCQKUhfnr+TYubKX7SMZxeFfDmNvm2Pu+Y9cL4/jDjGplHiAyqYzCMXt7fwCKbS
CX1Q7M1Fp117ype67p1YgjxiXFoGrieFsstP/hy1yYyDQ/WZmwOeLEHVAM6g9N2PxVgKz7HaosnR
j3eQGc9blJ5hmf/Y+cgrt6eQh+nSC/HD5pYfqU3maDnfGEvL1rEr1AvERhgk8XS1iBuivRoXonmV
Kk11QVgrtyZSEfQ5Ct2vWBRYBm4/2Lm5cfPG3iyoXGbRBRRMSkJEKKQUdF+dbTpDau5l2dNStuTS
dHcqxouoMfoC3I5ONne9MmcQnT3l4NU35aOCB1UQCVY7IUrdZf7YcOd7xfjq9MKDJ8tCcKHbzH5N
yZzwBilKWTMz8GrG3e5WoroBj9rJ6UGwz842mlbOcLEkXBTlyK1aS0TfpVopwo4UhvcCtPkJ3QoN
xL5aGciQHvi2KmXhMzZBbyKPAKydrwBeafRkSrN19gbr5oYQyAf5aZVJ1Tih0A4tbTdimLM/YiGR
O6ahgEJtqkPdC0e7LDWceWerHl7eVM3xKUfKdf0qxtZ5XZjHB0/xvcFN6u/XjYwNMa1sa89MUd6c
DfRmte1bLeHx6+8AsC4duuAkUVbv3Ga8UJVFBPT9oaKIdjizpmZlrlxtkA+XJVkDvQl+Hs7vMj0i
mVQIaSGs2Z3dxSRVoH28qbPOwj49tGJbOMPlQld/Ehbe6WKiMVt3ZafpzNuSO4cs5QZ0rCl2sJUa
wZw5g8nYJZipcp5L+fm9LVsI3wIB3/AeGjSQN2/jcNweuKMlnzekgPqpLrLRq5Plb+v9gUrZVpHu
RRY49hfgwDSoCGGOI+W6a0t9VnzfzXMYC8GM41GBr9Xwth7Ds8ctu1qeCzfP9etz3lT+KeDNVrgG
V/xoMFUlvOZL446U2j66teWZJWd26xYDlQNezbMMgPUyKUuQfJa8sg+kAKGCPn/geLlXD+BSiyBb
N8O2i/bY2JFTu/xwfhLYPe1epZcph3/ysCCiTuFPfPZYWM87lFNbRhZUlexJ83bwuFhUSpwsPXe+
lSlclWhGk8iytwWzrUWSZfIpkbRw6jDulMMqBonnLgliKrSeJGrYMCnHmXEeKvHkGYl2N49GxgUP
JUoIakMwPmdcJCMgj49mCf5MgHWag709USNjZRflA3VuKHxd58Pimk2PkvFeW8Xryq/ua440fhGi
1Enl/rpGbiMr7EpRNjdQqhXi/GZyuwfkXo6w8QZGNc7PrqFnqNedjSUaX+iTj7RGZti2sj9fNvuW
hzvw6REzGcR+kSW7ZbaPEkEV1G25IfqKr+rQfp5X9CHP3esVlaFPuSl66hbkZmDGtV2eGkSKN5z4
dgvgc2uSfLV+4+Tmo5REKG7R3EzXNp9+JYd8MKZsm3IjMcN0it6sNJCMDsW3sslsrJl3fOAB9nAV
A/PgzOmZcDqaWe6CvMWEXaJ90P5tzlxg30CDb091QdxZyv5YHwI+jYz9TofBXdmX2cWPqIIO/svC
HBglfvYxt6kzS9Sy7/MW5lAqwQ2LbloR47IXnml69xZBryiVygvTA1boA7t40BTzS7rRREi7N+4H
2TiEHHtWKWm418/TVViJBYT6okm0Xsri/pKpQYWso8vxgDMIOkDmwrPIl2hfQ98HkSwgu5+k6EHP
SpiWVtmRNeNwijsH72P24zOgGDfPvBjwWESFLbqOXSA5gzaR+5b1eSsSXOdpcEPL/ZgBPo+t5aBk
q+ZnGUyyaUUI9LBssjXCB4QG5omZmAUAVSgXRFmAqgf7XMaJGlmdQNq0lhX6z63RChrzMfNXSTKR
B5JE4ibW5KZ0fhfGnlTEIPB088TA9LxOioZaAcVBOIF5fQCkFwg0WM5/bsiPdCUgfQDdjvA5EeGX
1oyJstsTJI3RNNkY2nWKeVXx+vkCyb2RTcMozfCzqwgfWbcXrPnJTESrRIge6oJZq0cAey8tsWCn
BA4dK1Gj+HF80cPJr1cGvp7shJfc8eUY3b+svOZ9152YdMroJLwZhXuKlX0bb1XKI4HuV7BJAkzZ
kc/nz1t+3eqXff0MypPtDD/3J/HAz6+0uGpI3PRSYXN1JyvOO8e76ntpHU4nhK7tDcVEnuue3kXB
Nd8YcRFASpk2Uj3gA0VQzCsSBE35faLGXEWYWHnEUMe4KDSsZFAgQ9aQJD9I4BR1DRqbZphZCgRR
UPLc3M/qoJ+Y/49GFHJ3IId+6Ngcg5H+vcfYdKECRME9W83/y8Fm+pZ1juvo6h9MwIddIf95P+KY
B74Eu9MPntcKlmc0a9NgO6oNFfdajioet3cHS0hn+OVeqLGf2wYQYsYkcC0gUd60Y2gTY+XDaZyG
uox/tqddPJzDYJGZwhYTg/E2j/3zTE5doDoHlSdRjTNuvpa/Wo8DxYXUqQ0AWWAmMDp8t4jwQJxG
z5dPW9t07CSngHjKL1uZ4hbuIE7tcW/kPuTzLmOXAlgHKa/+PXWkRNE1/GXTsoEr9ocX7vYQjNYE
qocJPTykhvzt7hKffX261qlH8dubFVqH1Z976rMTu0pcJNWkSCUmDp/IyQ6tqioRDSsc4YL9csc7
7loIPWsbCBr87Tk7FO1ipTLeYvpzjvWUfrJxlq7khc5XOv8A/i49iXenwqPV9aZi1CjZAB5FOiox
vlNTUpAi4BfEVh/U+3cSZAlXbuUnlzgbZ+XsvduJMHDNQaZWoBdj7ruiM7AXG7pW/8DFzQCKsb/2
TULrqGU3vJnwULcawjOOJm+it11pngX7/xmbejecJc5Sa5jE7JHZAKGWnQpEb1uEdqWX+MaLQUBt
XeLVKUhi4vWfjPAa+fnReQBlxRyY3RrqYrM8vCwmulHHFjBbMgNXove/1pb8nYIZfd2ROULTTaOO
RbGZ84BGreKYzdJJXFZh7hLq01f+fAv3VqnUnk6s1g1aRA6X7XdBR2Gb44YnNL4GEG/ESHFBN1r0
qvbqh3MVg7Ub96bidqqNrYOEhw/2d+Vo7cCSXlwrwRyiN020QaoQftH/pOEqAO8ZDRS6JwoMEHoY
PDHiI8mgnsN0v7GxK13mS+7B0vT1sYn5snFUGxVwtbS+X4wpVDS786zPkXhL2VO5cZEyjJrSapgm
feD+pIY+j6jQlyjZEhjqkMOVXBMvujcVNAQPvwJloWLKAoNWGxjvqdcVF8QXRrkntTxQXfnn+xml
+Z0PS8CSKPMKRrWMvj5VPzYZmsIVQbhOM8gV3kvKZpLt34Jr5B7MM7RWIlazvFIxbRejW/CG0588
sTTgJAod/KALhmlzy/IaIjeYY9OGPCm7I7hpvXgvSI6CgmGhW4wtcl2bVjUSQn75avJWy3K249Gr
ymtaRvUvli/XT4OEK71EHSuKNmkl+IEics76H3KNx8tjCwANZJctOYjEpQvUi2TzW06rR/K3BD1q
FK+5tLDjGSZo3ww7NBvspM0MOjfrQD9smAXbNYqFFfu71ErnWlHUOQ14tM0/MurXdB9vP8f9K75t
FDXUlPxN7l5sx6JmIGn3YWnXZ3HyEVXCFxEQTGARhbWjrzeRLoSdUL7VasDFafWyN/tlpeZwdmD6
KdmN1h3Vx/zPbxelk4egArbSBT2EmeGTfmiFzHEmL5MYmf2Qqep1WvY5tEglA3OIpO3VMtClGGNP
YywUI214AEv5ryiu33DdblTtCPZa3j7gDWuGdXzJw5RAlInqpD6lC6/8HFEGJW84OjzysS1Cq8DT
EHC/TPOIzafeU7Njl+6CWLbuyW4TNhlLtITnnqGoAv58NncudYdVSJUSAhvP+Ma2vEA6H1IJfuH7
181pm7sEXaTe1OIDYCZ6864fMcx0AowvxKV4wQ2a2AvGI438UrS4ikL5TDTpj1Dztbo4uG/rKpJ2
iX7Q4jmJ/9lIfbfdjITQ73aQhKIA3dC+Vry5Gp6WEK8BTEk2mhHAxS6J8QGi65N4zmRqG7FzRUNC
L8flrXaqRxixVWgnIPuSV+7yH2ACuVK9n+B/faR138W7DrzdKbb7ggYdjLmwQih9QpxT8Fb2XHd1
Wd/S3uV/dg7fmow4aT+H/0MKf96R9zNneoSH/9nO1lI7LkzGJsHdnUaob74712B0pUnTOUoJua7K
0/0KkjVWpuk3jkMZfAUTzoWCFG+PmzwxLW14EF/+BjRsl3xo1tbyFEr0zCBVerTF4PGaD+4yMaJg
Uvi3OGAytFeSgG76JSWSZ866OqcePgxO/6OCh6/s31NE0CjySl+402mnqMb5Z/4TGyBTwe3MurYh
mS+FowlI94oIs+QckEOCB7R/ZgEsrhZJTpD5uQXTSUgn1JeZmi/4T7qxcKFr4K7K5kEkbgP9Qtyq
2MApwJtaK24dmm+rOaP1RN6yM6i7uanRHZiB/JSylSIwfMvlngDHe9tCvQinGGW7+G0Qsh6uJybF
NZJ7U9x0b6selEdR3m2YEOKtjp7Yb5sKY9Ozd2hVMW6cmlxj2sKPvFbf/sB9Q6vh17CniPYRTugB
iU+tK7MGYU5HgKnpDa4YKvF4+8/xSByB18muWu0XRDdFjt7eh7YlQZMMypTfDYKP27qhwuO3Lyck
LaABcOphxwOMAjfvBn7Qp42qilJcP+nrV0peEw44vlS0sgXPTwpyZmDZmbFE1wo98786RkF2T/cU
pTGgKfPk3tzs7Wp9DBKHGA+qYmZ91wxQUHoigvgYhShDraPmVmUZV5l5+yJqau0QMyn0emzhwhkQ
kQExwRZJJoNkFiA7WEPF5nPHgoUYQ9tjV9K4uLaRKGtDdF9WUCT/uFndVQNEYDjVOQ/bBytU89Tw
hkRfURbhcejy1B6N6xc/xER/4UvsQZhxkDlGZ2uN80VK1Jw1QooB4YtgXnX8yK+949zViw+V37kJ
mvmLYd4z+Lrn5EnO/M7JJiAfNFeY+7Ph3fSSwmlarQttnZGMqkLB0sfdnT7r4yWGZ4GeKZzJm+JE
04ftA7T+1dTLbIX0BKE6k5KhMOdQHWq0aYK9auSaxm0TY+JrVqquRPGwTAK0LymPeCgjyrfKzmjC
5Ib2t7LMumMDtLi2XxveKrMVa4AZ9WnlgtJR35vlZQCUSg9L7voIVtxymwCMZAWJy1XXCC7WcOuD
uSpvhaDzAbxwg7BnizsGtEdDG9Xg3mTFOUrOTn6Hjjqe97Fqtgb2phJYs+emkD80gcQbeQtvywR1
/KdYARNpQ8E9kwHVwEuNkUGHImroRr0l4cvv8/evCtSwXgz8NNplmJ897czKfBXvrozMk/duBxd+
VLWA12XNZq8H7tcnWml5l8FGdrYZ66+zgyB06QcUXZG8SKLocfLhYnC4oGDhyIX95DU9ZA3Nh+V4
0n1qnujaszeGoesZLGe22BinI3iAoVjQKiXq6cAGFHUiRGIqS9AbTHEK/fdEbOn0/Tjyk4HX7bDY
8RGjT6rgDetxlvtL3ENVFSlXmPBaFLg43ijQTigaDGQZLraxG1yfdsYW1x6ZLJXZ0gtOOL0dvIgM
HkqMV//h+4J0iF3u1NYy/kkFsZ4ICGVYJYErmWx3ZCNM9QIxdakldaUlSzW/+ZbdEsH13slRbVmW
U5ABahZ/dhAApJGBk+Lpya7mNlIv51c66n/3Rr1zuhrIUn5bdeLNVlfSu1/wrdvj+obQgsdopwsS
IB46vg0+JUNecMp7/iFEvei0MLZ/SYM9gcoRsWvndJr0bkPb+FfIURWIPlb8dgiZJzs0BGNakjp6
gHc89tQ5JWAlmbzrtmys8N8eit9D9cmuNAaNjoOQXJbcDUGpZKsmaYo4nEa2eIhzTSPPIxbdMFM4
qxb2O5Y/491rsAqLOMz5mUocrhtREL0akwrvxwYaxJYFhk7vUW9S6cm3mSlnaZ012k8SNLsdK6QH
3s3BBmwu0xR1pKJZPWgBMvXIGysoVW8KCQTt+PD6GuuSJjvUMG8zNeZJd67hEd9aytoQ1dOwwtHl
wRYG0lUBJeug2jQuwk+k04HbmlUNtF+VrTfwq8r1YTbalkAFEudvvG8gBBYVAmUAZqWB1vqe+s4M
6zBms2HF+qv8OIISeqMB+61V3e4LHIuotLPrFrg3H5Zp5/meAzer3f45Q5hmpR/386TFSfrLFtOZ
wc8AJ9in+mmbveKzk9DLn/8b5fnKoWILrYgdLYMPSE5+YeeIiIFJbxaPkLp15prWWh2lZ+fNO2QV
vGm2FQg7tpdUaF8iaY8f/W+l9wOCkj00YPOJTi4uAkxTDTQltzD30NPhoXibp4ldAe1uHpj9+mAj
1XQ5HxJqmPOcA9Qjr4l/Q5eWbAh870MaOhxv+Wf7g14WLsk5CdNd9tXkqZoeKFAkWPM4CKUlEBTG
MIKAE5tA988GD0MiX32RHQWww4pGXYj3z9ApP+Y2xMYcHCAJblIOx+J2pFb76g6sNawGyrfO2TYj
X235VLK62jeTZitsWgNjBvqOXWCTaj8CjrDqAr2dE1BQTdEz9AqgQGxWHSyfdubZ8UwHCpyz6PQA
bMKHRI18jAnFPlCmzF/fUYPdF9IBq18OoWkPka9dTPBlAUQTldwpLjpOBg8vYKF0h2PqWjBwNIWW
LLUXjACKAg79Z62XZltE8XA4wtbt94sinoD9MyxqIlyAEYbM3HCuv1E0FnM0oO7FsEE4V1viU9TQ
81tt7H8cjkuMyexSE1dpIfjAXHUpuCDF2pVVzsQ1hueLgVWC7wgvVXXLB4c/43+OvMPbHS8wYSsX
boWSOWN3rvXIpRMEx+WE4e3TrjXZOLDn1SI2xztc3f3gbaUwDW6k+6l0JLTfSn2YySH22WLD9dqz
tVevLmjSVAucUHsT+JQHo9AR0kqC82V3bb1L9cgSZMtW26h7CYBY0I3gaatj38c6EBj788ZedRxW
Fgt9CBEnoOCm0tzHvj5amE0ldUjjugGGCUhBRI/bv7jWUdt0XnQP3LcGKjwUfWUminxLmAts8tN4
eBzT+s8Niuqc0MHBrlfbZDvE3daePhdThQoghCc81Zi/SLnzuyaXom7aQ5QGYY5KDVTR5HURCqoV
dfEOoQFaPKzZORvtvXhs2ad+rViz0chND+GzW6tbsYvPCXH9zjhnsxkYCt/11IKJXgS7HQ/+NwoS
2mPOkKJpfD+L44yAFEmE8OBPBDDYNLJBjKSef1i5Cd4sHquYtH+b/gmhlsZ/DU0d9rDm96Ldu+O4
0nzwDM/hHmgS+wNeU7f975bzYKMd/zCHMDwto6ztrE802camfqI/V19Zvfk48KjfzGa9fQRMzZHP
q4at3FTY6IOi/z0bkTmGHOmf4h5ce+aWZVQb+04fpMcrfm7e1GgzxINrtqmJv6cs3rZfZsu+ovNw
VvemTi7a/pr9NmpiUUKAFjoVWLBcxvTdzRHvcD7TfFNaF2y9jkAq9oYYlsNmTjE7Iqv6v6hreN64
xANyKoSql1oP0D/2qEg13fTc1IaRRGNYTR3xNwCqzQZa4ur55iIICyX+wS4kfOwnRxwNX4xpu+yl
yJDPwld5PpJ+vc6eD9EodbS6celHFFjtyAYEaTvOvUuqscLV9iXInNBWSkeFICPMXc/yQ+7zTgLe
XeZjNaBfpv0VsFGE8FFXe+/FbSAOYv51eACVcqWn0K3+NsOuvUDIFBzPLCBpHyyImQIOS/9QBeND
KxHIAImZXKDJYLr7thaIyg03Wq1XokOAGf3IGztowDsIYtOCEu9C2XR7uADmnwYgYTGqC6lh5cbL
+r5R31Kogwishjtn0ZiVPBuXkMGABgBQEc1PnjOLKHQ9oUhj3OkDZwHWdj7nBWlq3J/x0qBw9M+W
KOHzkNHdMMH43x7od6tsO9xYAue6Gac5fQeoMLHl+YHDXiJ9oQDqwjJdeM2Dvd3u1eJfrywzQq1X
av/4RLA8d3K3YKQJLexhYPLwoS5tYYUzHkHIjTj64qAChNbpai2W4UG1CsLnTjm1Xdtge60Pkh/e
4NTha/htF1bGrz4oeY4xIJolx3kPrp4PP2yRN4XWdR/zMPQKGgLOi9MCOyd0aid88L9TXqfyNOI3
6W8t1sGbIquU7kAB4xsSek7bGu/+i0V7qZqaPNO+k/Dp+4ikmk5F0Tx5rbPo1N/1uyl21fOw7+Ro
EkjJF0gUx2+C5bFVnyUakxyiNVCTZDOtrh5H60P7RD80qjNxuwe1S7jFEegUde9P/IrNkEr1p98/
5VkoM/A857ZAB9v1xg1rm+e9oeZdMJUg/X+KSsS8WrWd6Fly1njFj7h/UUaurRejX/zuCAUjgVxR
Ou5Ck+QHsTvWd52VUUJNRovyZ3/xKzE4ffc/0dZWS4uHt1n++zxt6o9buN6Y0znaYFxNYopUeU2j
a0NPElzC+Ob3oc7OS3o0CVtMzXC+Mb3IV5rmazANcyKQuwCZGz2CGs/J6pZvvnMzRTtSPTAgotJR
KPSicUybI5hZzYANOhMS8xbU8qI6ExWItm8+ivCbJ9kNOYGTfrCW0qeVohj2UE/5SKoyymeRJtZX
vJ5MCyLuwJLh4c9hPaqkrSjEb44ZGmz9Ao00eX3tcKr/DErsq6ikdOZBHp49CflD8i1qibCMmxEN
UKE+K3qaa+ckZ69cPbJJdr6mjnZP5Q4psSVE1qzT+MXLKzlUfyV7NmXbpb1iVX7CGDwMOp/qs58Q
TjNfWzFTIqNvi3SFYqSX/FoHeC+BuwH7Naa/JER8qLqOHFmQF++SO4boSi2l/lNTF7T/ikVU7a5z
hi7X0G+SfCxsPnAhLAtchPKfFSGL54a0c5ui0fLx++OROP/kAzqrNrZzENRjKY/Seww2Qd4+FyXa
Jz2OLtPTLfFryn2H3zf7BMt1wnrRZRRTLGr6KdoJX/WyDjHJlNNSfhSWpE6Q+96zltGbTvatoJ84
lj0LvhBzmTUqx7LlvoSh53L+pZual8ZTUcegZOVIrTpW6/4dRvhEKevA+wyE8Gl+CJI3nIwThcPh
y006yAIO1/EcejGpD0J0b3e3JTQniZFJXJ77ZPfkXWY1uiEgJYwIH0eCiP/OeBULbLmC2Z0EAFah
D6ouivTCKVo1+8t+TtE7Km8IhAW9oPgfIT90FDwbj3mGTNdBM+fXzv6/40I5G97T0bkFTbnaGaNp
l7TvdyosD5PObSY/ft/VkLw+oAZRispbFWS/dGtu5HqMOywKj4nguDB0JXcz8udt9rBJOKBWkc6a
fU3TN0OTM09XFbPecbh/ZXTMn/Onnb+VfySnzkbq6l4RWfkIyh5H1O0fVzFUKNe9P7QjpNDqSmzy
1RMDgjaJ0nUjKiiheMmSVdJccwYiYzhFiBnrQNa1sR/A9dzEU99SkpNYyAcvtzlsb54NO/mFsGkJ
lCkqIAzVXXDlBk/1F8K5ApTVHRdeSAZZdZ7T+G5YdDWoldAXw8r8RDLgtZQqfPuskTk2XiVo0dB9
6I60MZl4lMiROJwTyGpADfMOjbRPZrd4OPcOAnn9pCfxwzm9pf3D3BS5z5WKBhGecZy2Ua8JBfa+
Tv7s6s0CnIqpqZDUDN1jM+5ub2HlcPh20Syh70IjjWsslpp04/rxGOrhb7wLMHYdTtxFEGogk50e
ndj2gfmX+kc8SohyYcxf9dGjvu4qupGJDxtpDK1z2UMV9JaGs5uavEDLLajJY6q2Pd0J6Fn8nGfD
Ki+KCVks6E4zD/jw5ack5iggVO6QJF34cfKx7/fN9/ipKciIs8hMvS15YgGA5x+LNlQaKgyWK9Jk
pt0QRKLYBWBIsFATvj0G2EzO1tXNr5FEw6IN2dQ0Q5fu4Tpyzs27k9AXW+gNIu+PixITp3X+Sjk3
3XHBgQOIFMbxJL89hb14hogsivcCdG1iqA/3r4cayhGdM2K5qdV92+8GQl+w6CwpuIfc/k5j2ijK
H60sTU1snCqDxNc9coLX2sKQ9kEfPuMGZnOmXmI7I/llUh2xHb1Av6KnhDYqla4DeHpbjLSSx9z3
XVatfBJX2dss2WApOi1MocCLE727aG3UZstx7ZSPQ++XBVxHWl3N4xHHnu2ktS84qLl0n8+gqkfi
Ra3BgA2ASnNT9DRTYEQAzb+Sfl3s3eEeu3hbZhb6ceD3xus8bbex2SiWOr+6ILJdu7avbcmsrGzb
3iRMgyHQocageH23svevjzsPe0/lh6hIYv1SHAcxgcXEooC+yCoWY6PI58eEAIWY4+Fx5BhscbqU
4vcYFTp7yr9iRuRyMhvY/XrlRVWH0kcvhAdf6rCisFniJABJk99i3A3M2g+5xCyDOWHvi4boUspB
vBWF64sykwUczbjRe/kumUrwxnCwUCdR92ChCENHNaHnaCBuw55Y6MZHOG1tBnyzwnKSxMJTgSU1
Bvh/W8tl/7vrJhtIpK7yohI1FBZH2Oqih5wCULrGxnQOX/0ifEd/M0fzorA449DV66HVZ/LjIgIM
TsyPSqaD+BWbufZgyOc0/FM5YOP0CZxe26xYXzdDo0esrdeAzo9WZMCDxNvZJjdOlNEsvIIz1SY3
98prjkOU5LqPc7Pp0hJDUdsFKS30RtIWTauG3Qs1AO4s9O8q8xv1BR6A2k77LgUp7VZJ1Aja11CJ
KrmwmkNlHEXeI47moY5cDDvVT/A0HyjQ94V+iu183qSq1vxKiq36ivo0PAFAmaCfBU5wBY+bU/30
cgWaZ3AhKsje+QlONtY7xQU3I+pGDr6/SILosz7w5My11zYm495SCAM412SbxDiF8SO4fhgWWh8L
jQYJGQlur0JwxLeI3X8DHgGG/BPO7c4FsO8q+It+53iLsSCSoPKI+mAh0LuxQsr/QNcz+CJ1YyQ6
62xuzgs3RCWb0OL0+G6fcIYGu0AieNkYE7KwNwM1LQ1x21AEkVIb99R421+lUcTQPvTp2o8Sj8JQ
fXe6seET6sUWYxLUcgr01p5H+RSuIFAyQQWk8TGKf5EMS8drXbsRa2qzzXX/yWh0zjf1jxF/pNxx
22T8+Vz0/ds4urfdOf/y7+3LExzn+KT/Lh25VmIj3oDCa2oAc57f3HdK6Xt5P9fLxE+8r7lEO9tF
pPR055pBTgxUKNlPNXuBeYfGSz6IOXxAi5wbahKGROb4ukosEAHrEFUJfhn+O6/5cqvYt4iNTeBH
nQIj9RkjMzqpv/ZvUQ5MtDlgK10gPUWdN4pLt4VKz96EHFlV3fHGun4Lh4DCjliCcybH6c/s6nxk
zQhrXXcntD+83msueSsG/PuAAzo6aBvyAvuNYQIRkoghRBMq3CdOTwFbOGRjRqPYX71lL4Yf7NJk
1I85YLUfpxBx7qA0Lpo/Yz6NiTR4QHIXWQkNI3YpQEoli4X2T3cB02zaJmLlql7qjnLT6aeXtnZm
JtvvB3rC3Hmlp+bjLfYWamcvkXPGG6J/iRo/p3CZxMxVHvl6uGG7GsjVODnrCePSho+60lv1uGXk
vjJxD/psA1KpwWv6d4r8XnFdpt34AP/o2s0r00PgbmSdTelKdKG9VyuEsQHiHaUXQQiGDe880Gy7
qSBMrbVbXFLwd68w3ayKm2J3oDIDWOVaYG7TCOeRzvOaGKnJj8tHpDPSD8zMkrlYlrjoblsViS7g
MALdvpLshZSOGS8+ZdnNFdTGQOlHlNc9/Iog2xM0zaYJACUROi9qw3zlF1gpZpK6I1zYCKaqiWuR
Wh3/8aGNSEG46AgetFJDYX/1QSF/Heq5DAHZFbJZqV8b3oBb7zYk7oYB86iJReALKotdYy2MTMWC
KvQ7evqJzrkf9GS+1J3xvlmJuigSiemg1GJJhG0cnofIMHSHlEXZslJ80A4FoS7/ffl20KyAw6y2
Af9k0gq0Q0/gEiupnpooLJRVZTttAR1RD30ZmE7qc/ZYKnB+igCD1MCazjHSzlYHz0aCxGiX/b8E
iwpyEsgqdjhli8C1Xo5yFeR/uVoeaJFyv66vDdmHNDfn1TNBM3piUUz2LDhPaZ3ZX4lk17YlomcJ
lTppnQy5kd8mOXsFcYlCOqButONzP6I0n/FcWXK3Lklghjr6uSlWVZ51DDZvtgcbnSA5D9FgEil9
RsTUedWQv5Hs3AbYk9/LwsDB09Tzsrm4mW4FVwCpwb4/YITQWzUruHi1aTFZY4WLwBUnLnzguv8k
3+/3IdQr+TzmtnnjpLqbHeZwcb60a5TRbV4rs92X/U0DP4jOZAfWDY7lSK1m9FQSqTNwUhNPM0aJ
DvIjSopzWgvgMS5IG9eucf20jILqIzJCfyJXbBjCdfvFju8OApe/FSaiZ9txkPNht+kOluVAGLNm
Bc1hN81LC26CehnJHIpFqhS4PEdWDQkh8ADAeeUgM24MHK9tupgyqiHp2tEAtsOSlFv7F8t+Syjh
y91eXJl9jeqFmh6SrgLaDlhvOfV4/QWPZW2lWN6s+0l3H3nPFgrRCpeQUaQnc1PVaQhXFeFQk+oR
50ggfOQPDv0rYXxfQ8jKOsfwFdjt9cvPbAQUYDFIvfAiMZLQnlASdY2eZEmqfSaLsfjPohNKmxuS
0AI12lpJcqbX/XhVi0zRQy8CzP7K9baAPxT7cco5OLvyBa2RE30sjO3jn0Gry/ai8mfnbSpDCrPk
sQrGWM7eAKAFFajk2cpDS733kc3PxBZywsyAkEaJJtqb4dJpHYs6S6ovj3q4gU/5THkT/m8IwI/L
Br+KXb2iOKC64TtyTTedr1RDfszfD7kb1HDCZuEh7sTVxOdiYzPeDoxVnYO3MbuKhbY3gVB/pjwd
VeLoIf42tZttMrk64WEsi5YvXfqQj9mZtVSKulfHPx3XfDunHrm1a3KluAVRlFnSvZ8nw3VQp7Fz
nMoUiTiIEi9WaZvescZT1sm9HWo+TGXlTX7Zk+hrPHL8XxDHq9Sixf1OVApJjKYALECnOvqc3U16
J3cuU4yMFA7+94ZXu/GhuOwDx7d4x6yuKwmvepxzzPOqIbHEFOh0rXXezg5PkF67KpsBOhHyOaou
uCGy1iXnxLjalukFgSwqFnL6BQxTYQZ3JalpxHF308C1NfXP6ZnNOrsUDykXGsIAVGToUIrZKCSI
U4DUsO2rUmaFPw1CEPO3YYBc8iGqIdQjPMl5c4TpVB+rc+YuCLX3ffrbzaRdtTBD+2QjaZIHOxYi
dukbZb+EjIdQv1ByYrykTojfRRjtg6cuEFPhWLC85JYgC1wFqr+GmLaB/yO2c/jsOBVV0bXzDKBp
01IfYgFopYBfX/sI6W3VGlBYB9CknOURCAF5F1f3EHXZABkP21PAH60C6QHK565Tgrc0l5lZKylp
JI17R4JaZ0J3Dc7xCmmCDBY4qPddkP7pNt0YvlnMozbqlMeBLIKteJchBgX2BSF8X0Zu+JLo6Xy3
r9ND6UfN6sZoYH4GLfiW2TX7fV7dKykPDksShYuIE7d2cOYFAabQefgATV83c0PVa6VTcPcuEqf6
irYpA2LUwxSGMWIyVC969fsxim8avXaflF9kN7fFZxvZ72ncG3A+jiGdlk75UPA/4BHePZ7NxVGi
vY55TqqtCnxWvXZhiSqPRT/0sjt29fqvRc2gX34aN84iyHj3RnUe5sPBaxrJWYxKuSEd2GP54N0H
mjI3ZjcFh+r7qU3DxVHT6rcvqotvet8HnMHfIM19+fxVva/JMwLCp2P+SgrIDgHoJKBZFB1RraN/
ToDYGZsId84XcfV/hSDY/U8OMaKzhZdZNbcTcTzqfOkcIMvV5grWKX8wDYrDi+LxCuGETCWA9OWE
gYAPB8VU9ocbyADjgBAbbYAaldClWGtzMc2ITPYlKlksCrrXUkf0+dxOg+b8UW0QaiE9JJIgCE4y
2oZYyMdKgJik6ZLny2oJiHwvzwd8hP6CKsYniLWEcFrT0euont293spFGuyCt1qDjKRh+QAskuOJ
2avSD1avkhh5ptpi+Pk6KEuKWaqcY+/KSB59MSc+HA+T5rJI3h3Lm8Oefgxi4BqZcpr6q7WNZSch
U0K02ZGua8TnTNEwgq8LVfWh6qH3AcceAsCI+p5fY0STcATYyvEjDnUi11XT4pHIVPe8+U/XGavZ
3amfl9oPWqP+10IBf3eyhbGoG/PKyQGwPw4FuVUpjUOG4K5Vmhxd8FK0dVpj3I+JO4csrPCeJfvf
av5SZrkxBrObkeriivj3qvrh2WS/uakAY9eKKg9ZXYnJlvXEoOvwmHUoaGxI0e1vrT/1YWXyRXjF
5kWkY/aawyVBB3ZmZdd3TLDWK72vLW9/94sghjpw4zfFewcrwfs1i3+yK6nonSzm1YaaR749C3cP
7gqJfjj+0GbS3kIcU/pxJLyYVmwCKrZGZf8+FZAQBLFQFQCvwy1lj6nI1l2agKl+Mw8MBPUtLmL+
DILMG21Z2TeHrpCNaaR7+xvWogzj//qLgdaTAlJUgH4IDO+ymLNpfBQkw9yb9J6WID4FiF5339sp
vztOCHgc2flRAjhTNahSZ+OD3AhuYOAuR8h8ByVdzD1VOIG0DGZpg7sksUZAMH6FNjwcl+nlTIcG
Xt8HScb1VtnA6M2TGuhDDnyN8t4AugacSQwNXrFPw3Em16FWRMXyaUt8FtYcLqkoSbMAE2LUTvhe
BUtTiAxhpNg6RX68sf0qyi/9EwZN8Rr7XE75aGOCxwszhze/3LQPqKxZVQZTBpA2EDpI+NC9rf0k
IyZgtaexrv+YUcS1RfF16mg3Rx5adtGRJAfJZkzPTDxY+WCaqmzi5/+2IQYLuHRKYZc8FAW1kNlU
jMgBfagfesFK2jMpAqFKiAzg8T4zgHOFC1Gs4hCSLeRU2AGzsuoe1AGGuluPJhb+3L0gUbyxNrLB
gnbi4Z2zTp+sMJqVUeZaepjhEaT0dG1NjZSpqdSQgisAkqBnaoMd+DA4Gx20is6tYlXDCXCtwEXs
kj08uOrFPukn2oeufY+dpcTsYcyBhRffwcZCOfMo+rASusnRwHd5Hnh2Ar+13O1Dx//at4Lj0xjn
2NQMrtFuU5sLEyPouUAX0zwGDwCXevAlXwbbLTFwPo236V/jx1uiEIH8nuF678Wu93BpWuNCniP5
MrtV/bxA8waO3WFaDlOcyMQd1ptbpX83r5NTSaCO7amUpHOSwY4puT+NNTDl6z8Qbm1dfEXxIz/Y
RmR2CTO7xEGdu8MQQEpUkgpGyZjxFxjeN+W3l0Zu+N/eZxSzrIRk4cgrJAg6QGXc4H7iP9gRJ8U1
QWqAp/FGqplVxynta/Wcuo72nnYa70ydLPIZAvY9CBoMBz+Bl5I6awxkCjM0T5QMhOxuh8dHHPFx
d7hnW4NpB7jEACmLJ/SVs0JcXGtsBCdO9r20Q4dGtvClsEBNjUcrpghmSvUFQY+pMyQ9Dnx1L5Ez
iRFLJlzXblMoKQwCIh9/LbqFlNRf21FeJNX1jCVm5gxNXamQRkCT9OwN4aRhSfpZ7p+Ha682Mdr8
iA+/z/d9nv0LAXtMFE9b+8E+xgLTclP1RxBpfZ4lGDSj2NBVpkoQzwB0/z31ms+tPMYetmEdVB9d
V30I8dHm3rsegu5KVziV4uh5d3Bc7bOFezcmFTjBTgE93ThnatPYmnl0DL+sbMkJutF2qRiWL/Kh
f0+cvg1RkwwXWeopoGhCoMlpEKKyikEENfROPtm2GCXz9Smx6VLyUzC8o51A7OqOlVTj8WkP7ZcB
03Q14AiRoBqxS60CGv2nuBFMUOSFrFeyhkWyDvMS+rvBOKt6Jn7+UICHRaIj41H69pwKcPdVa8Lc
rQ97OHbXA7ts1tT7jHF4mJknEVI2iRDD7RIx6vDHWZibG1+31cVXROvN15NZ4o4uyTRsUuj6mCri
liuqqajhUT3kD8EMxzZ8NwIm4AHHY9Gk6g0i+mpTzxyMyaUSeE4MHQPlWwB4t0GEzki0yt/kLV9M
Tjy6GMMY1xwHHtArNbJJ6De0Prc5QYUpnGKxVbMerCZfjqLlIUR0DP3O6atARhNcC4dKjQedsHD8
TQqY/TDp8cc5sv74rx1Ibe8UsQs53tIBNi8dHZ98dNoizFTvIhvmpTxY6pVTlSIdS/NCUjUgeIDo
2PjjE+sax3ea/ZKV2WIdFyzMT1zehZokJUfQIxlXWdrB3JkINnnNfjTajJblyZuvXjH8jngQP+FR
cyhJAtBa1EbbjtY9EZEaSrZ8Fxe9nfXbPLgGWjlUy4oFlym/jTF+XyHmL5UQd278YxiCrVGKydFz
HjOYJKFw0k9UTp0WxzUtJl93VXIfUyFUpmpTZ2JiAe25XNOteWoVkt6zkUWrEBeZYuaryu0vZYV5
r6u6mCVv8ihfoxCVfk2u4reiu3/smy8PYW3IdYE5C8nwtAf1q4/393ZSQzjkGF4n2o1ATXGuZie/
ioA/BZzFbAUN96oAMep/u8v+qEtltG1uabF+kJy825jbXEdtlLunEugTehocN6VDrHzoBGltDRaN
p+UsnW3vo8+0eE6yKTrKKZWmQCPI5jptKo8ioyIUN8LuR4fNAzy6k0SxG2JEAxxpn6QDoFvtWwsd
AZ9affn+Oir/+jZxpPHWQziV+ID7PL9TCBbNUde9QkB445RNGwwNAokvd7LdNCnLD29yniGsx24m
h9ceRg7pN/qIRbuVPOTb4/uoQnP1FVvPaWiyCQiI8+jjuaX4RkjP2f4SAjHssabuT1GVhaQ2Qey8
75HqmtGt3MqaCm+uQzqiSeTlIqFhs49DA+jK3iDBUgWe+ClyTOCbHPJvJvuPC6i0OeSHpn42SI+r
d8zhjkcHElTJltCTmTNE8cWABB11j1CZ8LRLeSSKzdYE5qDed9LuPf3/ld+fdINud5yHwUBaQ6Ae
JiWk6c/4ewJwOhoW6ndGhVEAPh//NZo48L0B03+smAGzef/b9n+vsVM6Q+ceFqIdy9wDeRNcmyEA
qfqBOIClutstL0QXeyNncMC3DF/4vAe2mlwGKF1jVxUCT9/AmWNDCkBtRRGPd5pZnBRz8SWtwh9A
NPTIWlbMTHq4O3F0jJFTjoATrKxuk/RA7QNIFJvPw2qFP0eGTTyessMOZydlUfquTApzKY34GLs4
qVPgBxiIoCEo7bYU8HMxIAsHOymZ33tmFf94vvpvKIyc+KPl8q54YUFc3irARz26NOrBdczEwoBd
0NsXCNrZGUK7PGezyFKUT4jefjItcnQHLgqoOrsUP17z2jMcpdjdhUstgjGP02Xde5zMYOC34YIq
CqpacrDiapy3/G67KYI0lFHBiSW6LwlpgW30sFsJ/Bs0Wf5qvpODBzm1tUMdH7rBRnf/HFjGYIlM
4hwbvLuh0+MyHL593oiPiPZ66zTJBcowLG4psODEdv71DewYPG+hUXvsebvLse+JHHe0ErFHoe9q
h59E/XSOr2RgSbshzacQSB2DhcMHrblg1p6J7Mjd4jlRpIaotZebdT2boQ60zFDggo7KAo0FKzSq
PgGTjj+FLfRJd61WtMPh4fq6Lf1bRRtDto67cwaQjWuZcErlRXY5DRIn0qY+EdCKG5TT18st1XOt
0zCCE+Nlvg4gjPleAHCGR4iALiXmQhmrGz98i47yY+m4PVbq/gUgEOFhqO3Kc8WLhnTnRhLWS254
bXIqHE8yfvu2BiKLYz2o0/VrwLH8VHFmIikViSwMKvOLlebfp2YutOJOB4xf7gpflpxqozsQQ34x
sT0X7dw1x1GehTolraZjs/2JhiCfdn6RpWSUhHHB78kHvMAZdZVTsrAIj/LBaRFqCSS6z21UIdkQ
1KNIElswRFdXd6Y3kFqwxy9VkMGkEO9sltJunXp9fqLPvQjBy/JOGRyhzW4bAFJNHR7X1gIPTmsI
u4KDiyoCK1KdyejVWuKX7CePpCr8sF+c3QYmrDeLe7y+mxCMXkJjfs77cwAtlvrYJlH7QNvibR0P
WvFMoNnv7eJOtXx1jK7BuiJiFSWN8fwA8CwVsWIfYgVnDhjgWW2D0c0KuaQaDYz7+FZs5SWAPDEx
TsHl040oDVn0dhGRHXxa0j0YnMOS9xwCspOU55DAJ75AsXaAZPfyFQr0+IP8JG/iHG0lKp6DpSwM
3A5zd3Pwr0RqKlfwslt4Z/F/QuWdo+Dltp3GTOcYqtHEplPPB/DWDim2Gxalr+CrpIBiVAqihE9g
B2trQyIyhO4fF8uo+RiYsCQ6LYz7/t5SqJrTLogbzyvZXiOfQZWqXfKzWRxlDWZm6qPMxZzGi7cH
U5JbUfab8bXdGoCmGHw9AlvGlXce9g9moG+yLdZIQnliFgdlX3SRQMDYipfrNERW0xR5LFq8eAvO
OT8K/j1ZEtwvv0c8TXSES8L6MBk47kNfhkADeKjXRiWyBNP4BVT5xyoNY+mGTdLulsTV26v6xt+X
rMJdNoAAhwHoe9jln7XQ85FZ4EpdH/CihuABgR1PtMweD6PFGvLeJyjGeiAX9h3yzW3J1wDf2WhC
DACvDx1i9/O79qkU/qNW7Ar7/qHDj+Bave0gTVdazLPND9oPn4uOk+qya1ZORKTtxtKzxzz1v9rr
0g05LpGUK1swfAiqmIs6l/9BcXvZe64QrlYKiCDSC8l9yQ5fPlfLKji4lPPCxqks5tSrDzCBah/i
ox9zwqe0lbD1n7ETsM6oPVltoOEcqdY/2FO1OTb54p+DgcOHeZa/Efxk1cyF+TpUbDcU7QV3cy7F
VwXK/OayeqBano+eegMVe99m3iQwC7vApJf04yxMRFguPNV9tP1oiikCU7EQhrfvEbGAWl+9DEVR
WPLlNVjapOc0tBnYLcJ3uv1X6akk7UQQ+SjYZdmza1SQfDxkwACsT+IsoH6uPHoUn4+oaR4sjoyo
dPTc1qxtPqsx9QBREJ7/km9kqNrGza0/mAFQjAJ2ARb9yWY+PVYWozhY6GSchA+bi5Rsu6HlRp+M
9bw3E2ooi3ijjgxucO7n9TFHHmj5mdG0aqiBMapRIlQ/tDpJzBoE29UGKueXKfI7CuR6UyIlo8a8
d95l/UEf63jnO1tKXCNs9RxovEOBlv0dy/HnYyByBRequA9RrxI7s4mJnmxNngdnuKptUkDLIsre
eWpBte4bs/u2QOJDBRekNvwJcGeMF+luBnzcmkho/4apQZGt8Z4a+f3h9YJH5XyEvHtzmJX6nkLh
yVUIpEZqcyebO7B1qOQH3RxzeaTRNjyd2UYykvJxDVsL+1xnGZ6XrVrOuUkJMpcBNf1p/1QjEsqq
CPrucXz7m8DkqyR+lvwqBekCg0IRnOYkbXbqiXPUNwwEbm5KFEfNdpkcnHr/WB4YnWSUjjl//I0C
/Cu4IneNcwR4pTpPJnBHK6v/rdDxvXBZwcwpGsUGSgpdpCCTGsd9bJiCGke78HYb4yMmUXCN7TZb
1gvU5U5WtEpTk0LUkPjtd5KiNx8A/MngnNPhlvh2+Rx46RRtrM9k9ezERn5MR/y6gSi90c02MNpM
EmY17TT6Jxh2AADyG/V7PJYTsV/vrMqY54R9susAwFGoXRxkaowoFfb5JZRT8cOlZcl4RYfiZ0Yq
38d7yUQ8Eh2gcbifhFzuQUPLhVokCZBDiL8yRvM5wU+/6mxfr43kC0V60rFkUisdC1dQB2fL+gs4
L9w5yXTF+DSIts1Ilr/JCTxGUiE0PXFtBnZE110GOTYauhWTEZezUUJp8aiFAJ9S8CGIfcc3pY6M
ZVIznUfH+ISsdrEPTrcnXnWalxAHPN9CDfo5RiSq53jHku6Nij0Df4dSb0W4+6xhUx7iw94Eurl9
HuJ5OcoRWnFHBjeSndlHxQQy7/WrmOv7+BynwZ7xBKUjGWyg3V3SBhsaDylP+rTtyitV0SMpNH+x
OOJvQ3OJOcSDJ2XOn7gy0Y93p55r1Ijv1jaMJTIwRdBssypLO15VuoUFmHt/79aSecz8xVdTYO2i
DnfxXbtMumcVnWVVf4hBhlhs2V4WU+bGdZTT2Ss6T6ZneIVbHbY8GMv+fYVYLsnjQGZ325h/mixk
zJF9/r47czQiIJ50qrRGwvzE92wW4sfdj6v1xUA+pOWjgTmRTypFy4v3sHNbBv8vQ6Ws1J8F0BQR
7VFzM6oo+lLDttOfltrS7W4ynmiQA8Y0De+VmWjQJ9fSIpDF1iS7oqLVXaRYVCRLlNhrWssL24uU
Iv6DO2437iY0gOAtO5XXEcesxFDhIxwyY/L79toZ0Vzc3/EFA/maGtDZZYdprpnxQHyv9WGlgu2r
o3m10Lckv1dnqd1rKat0XyB+RCRIpFAXrOx1SghDPv61cjTwzL7cfiz55O4i5c/E69uds9pdXfI5
xazNc4spkl4Ls2gbkw8EqrUl41QApgGVzvLrngydWCQ2lC0skEFJTPyVLaUpGjUmWU4FHLez+YyV
+cvtFQ3xw/Y+WRW28Ne/7RBMQGlSXcgCuSF7QsfU7KEWxFa9nebX9vATzQWuvmLIIQmTQL3v5Stb
5kOfk9d/YN5BQyesdEKk0Kx/aPyBIrztsUCEEIZNQ22H9znKG0y46Ao7sm6BUUwW4rX5TWeyX/AT
2Nj44b+9r6giwovtIyclDM1dzotmMbhywQitUpxFr4axmzH2KbPSORnTeBlFjRo6Y/3i1+SdmuoW
vpJvr4mkEBnyM28ojkrD7qIPzSDx4Exp8msTm/aGEXykuN9oi+cUXoa1JkHPkjUQHGuUl3w2RmRX
7PaZ0rPtyPaMARpX2FfWm+FGwCCl24+HAkygsF9okGttSABseTeafNfce/YqML918XJxqOY+5BLW
TIC9R5MA9EF7OGcBE22j4E3Wgl8baglSEv0HUmetrmnUJPUSrbRLC1qWYEuqgYUu37NQRbdw26lN
fyd2CZNiBCIHS+9gOrpRzjY4vSQMhT9pO5ARfB8tSZJF0GPGmNPn1ewJTylSziY+iOE40ezIOpQl
g8OjJ4j4zB22bRbO4KvESDXTdcTFDFYDWvpTXiyCCCcX3Xlk2wiK3V+PPE1K5UzTDFLIeZ/j4riE
QFzWZdzv7dW17PemGZcUmjoMJZUSQKbRBoTDKbAYloc4qx1Ubzj6IIH78dqScmHPvuCUBsP6CD6p
hS4Bay5txlSDoRtJ/UetzpFl5AA0ImyEsSn7vN5/aVxbcA9++uYUVNcT0/EOiXHxMOL5AZ5VImx/
S3vs1+mMj4xVcw8n/VeBHknAyBt4NUaBxPCihRnqnzxAq6h5xe//+6mhXyHMdOKevTS4IbzqUDQa
GPcoPoSfdxOokQIlhhGYFuXQIs66XdmQzquPe3TxbWc5hNaO3yelzK8WDaHRJcbivVcYrG6s/BIA
9GeCVSOhx1taBfQjgQBW8NGRiPxDEkTWWlQBGPy4sEufZPTWtoBgwltTq9fZWiguZ4ptjeWk5E7d
Ysq7iqpOKj/dAdYQFbKXXnkn7nzZ8bUsX5UZwleJPyswqg40pZENUhzgKx9Wtgy0g7cA9eAD3Suq
rMKH+kuM5u5Id1cbYZN0JiN0VvqcahskXw/arkC9kzCLYY5YN9X8CrxWoDrNzsgYjVx/rpm3QTY5
MspQ22TYk7RYZp5g6g03qGP1h803JoY0KQo4C/1BwCV5gzDYVixkOH6BevYdRhjrTw+8LzjPRiDi
Y+1+xaZZVgmjtlaOMP0uXe6yaq2S2WuSQNazefAUzuLz7lzADME3gZGkpAlVJm1CfLfTBQtdHVaf
9jEVd0N+yMeBXk7QcXwvbX29duOMH6jWDDuKD8+2i0Xt3tqvq0ajYhyZbusVRtY8Hp8cwhR4A2GG
aPnNNIKfATUA3Is6m1c1VeMibnUnvL8Y1sIYwDC6gRpg4zq6YwzFZKCh/AIVRU14bhTeZIfwIhbK
IM+MxznrLFb2SgYTpG4fjKVryG8QZU8AlxKE/elFB3jezLnZz73Vfgrb4WXRYEP+uHRlZcqf/OC1
ugeWUH9Havfcftst8ODqut9vLNw2U04IHaSNGv/uAWPBBFdQCo93vxHqAVQdWdlbJH0w7FbvCm3p
F/SQbRDa8o4A2MSjSAI1fXJKHDxE4MMUjingM+A9VE5T/DQsNR4LK+RVFcZjvw54uVnpQQM9XV4o
NIg+v3Vk/Ainzf1IjlILF4AkR+27eO832A5zNqMTYNXnjbYuBjZ8KBLtJdwtOhP2W6kA9+3PMwRT
clI0494TOytjTyq6eqQ6l55Ybfhwm3KFkTlcY20IsTTvyOPdSNe5wrxFu1GtV+TdMViEZWLSgeWC
AuUV+0dAWBq/hF7L1hj4/mqEVGXllwxf/DGOU+ZrSYnJA3kQjQPf6JUeJgVGd4DCH9TVDJ3klxrX
tFEKPU+du3WoGDKUcT6wOFyfobbjpGC/PxbSyLAz+wTwVcfIIl3z5vHPq5A9qFvJ/5GxKO9JUNoP
TMKDm8mdR77FCq92qSW9bagBmo4FpJU+yqD1GKi8zyDW6oSD9Q/rVy7H+98RIx1d0b3odYzBbNHQ
xoDJPWNctPz1QvDApdm2CX75eSP+h/j75jkElSIUlt0HwZm1Mx8PQ7VWGNHqw40h80r0f7P8YsgL
jW/jZ1AlehecDxdRQM7eyxEtYfBlH8fG/Aw06Dgr8P1WNo43YYKuHXwSW9Wh42dNYg9SEXP3YwUy
4yObIBybBBsA6IQSoVydLkpN1FV2XAcGu8w4ePU8ZRC9SnEkky7RR6/yGAsz2jlgcDQAc8mtLzvh
+qtUJOju2Ikp8itYtG0ZxA4l9TAELTEryElVyXsiNf50wf6HFL2jNdv/EyyBbpGPP/ew4J4fxtM7
CIlhIoZyvIp+ZEdOcqhUw/yuvCZ5qGh5LyyGd56IMEA/c0IsEuIFn6/v1jj+LSRreuX/CKau/t+i
XtDRHzk0ixn/1gh844/ZkV31t26kHu8wxIdkPxvn91t1RMOLkxHc/IQ43MBlUzpr1ueFOiC2WIyk
LUQRqKNFOpWqoCpChqNr/khETg6viayDrtvr70aEMRI+BH60DAw4zMLpA1/xd3kjAJaWwXAmOkob
+3AcnSeaLK34OC0uuFXewQt3UxQXPUHoyo+8RpFYy8CY9l1/GSje0e8NJdiaqL/8oWB7BqqEuB9m
MiIH6J9RPoS1shjR2Rjeu+8zx1QehEKIvTO+HgDP1XR+wHUVR1AAcxCDIOa6Ftc5RmHyMlYBtGLu
XNTS8gMQG9hHjgvSAdKmZJPbfV0HJ4eaC41maY9KDFTHYA8GIsVG2Fask7YJkJc1NYD1+Kjs7hwG
7ry9nD5SOPe4rel8pcNh+NmWH58fVcF0qijpobW3E4bQTr8pxNQs741G1G+3o+8UMZEEFqfcU582
uSBY/MzmniBBDjYT4BR8tu6a13/PLQD2Jd8ZGtfZJ6ByyE4BlQBeryoPV0hFLyune3VROdiqsBTu
fMCPRi4gCvtdlG9wj9vcgFLI067GLbCZ3sYXBhm2/sP3pxLHbkr5PzBNmjiGD4ZvuMwC0KGAAGO8
FjHyqnfFo2cyxCMvUb4Nqum1AjttBO7i1JxUb+u9UlXAnI9K4JIhzAUOBRW8tfWduAfr75jhPVsZ
GUimzksu0Pv7b2f+eCaULBrIZOzKA0kipVMN45PTUBIZ8voNKejz5PVKn4bsDEKdjkZDsZpq8RB0
NuIFPIR7jR+inYtyyiuMp9nVVCoQDDOczfXrzDCPHcAPQnceukGrXr/BrRtVz0I0w/erpN+ddzAt
PQF7ruIrpJ3oaKiKcy7/TBfD8JUeqp8ljZFQ70dGKNFwrNI+ArSslr65XH/pmszZgrhqPslJtXa9
8rxeFYZtV/GCY7APOD8cRe0uNnLcvuz663rIOJtGYP1fAeeFVLmgfoRhYdwHCvITiHE47lo9MYzR
yFkT6NWxq7iyw/epvu16Rft2BFab4DwhIrEGa5qrP/am9vwwbZg8RDbRXFXl92iF6gz1FYk3wI9I
NWyDhxqVsR8JCzm9dalaKdT7/L8x+aKU5EAk8RCuSDcj99u1dRxo0/3GAXZSI6G61e67CB6uRxRf
yx/f8h2WqzCoOCaAKYOgGS7P0wO5EL0HJHEaFGykXVzEj98+UkqhT6g9dYS3gbtaQx5JaMxdHbzM
L/n7uf51LIK9/Dk1DmdzfbgwfUJhejjs69/4WsD/E5O6WwXOkxUpe2LdkCq9O+UCqZk9x+ihTdp3
ndjmU0szLHabwIRGgU/bWcQo5nuoDXG60VWRR3snzdzlcckhe7DBj3X8e7SZaALwNi7DiHSaB5vr
Uf/kkjDcGLPSU2cI1892zVp4+ypDxlOdMmoOVZqSG5UN4JhxUcmGlVqcLk+Zdc0FNyCzThzqiRKN
GPSL8pw38GdBW4oJDHVC2Cz64Iqm3hzjFnRxoSjMDMmqWsf/8gYc7c5cGDicH8g1ffUIrBdeGa8f
W+xIQaGTqzzYWucrTYAQMS4MY1u6OgQRPrA+YuPjQJIQUPTvwuLtpF8y0v9uggKSw0lOwzWpY0lf
HmtSP3Q1Pjn9WbQzso1PJJB1tWYgurWIWeEyiVlOHsLYvyd0hpzUm3Tj1jkKfOGbBPLj3cxVdUFa
wi8Lfw5dLt8gJcc3tHnWoatVZqpYdMAkhVXVi0eVk3+bFs+i+CG6oCNrA5a2fpjEBPy0+2W31Pa2
OwbSgQFwAICQX/nP6q0yaUWAu43UYLeOwT344a8W6LRAK/BMlIawNGIGq14OCGfmfcgGF4AhIBMU
QNYneLR0Mc54jBsQs4oQQxmQOCQ+/+wKPW/8oFwbOMgIbP5Qyqa4Tzg+bXfKK4IBcXzQGap0DfMG
/OHHEaTRb0ehsmdK4fFBvNNMz8rE9PjRtGqppHo5418G9Zg+PFbPu0TkKKlUgo7QKQYSisev7eIA
tlDe2gF4wr3dFuugZEz450RCMXtDG3y6CZ2z4zsscddogszZ2DveLoUyVzwBCXwCLBCobJPl9tvm
CZG8tBUE24Ql/vRmmoQzfUY8pizUkICMxWUrRNi8RFV84e6YuTuGDZ8cZbwLsBzYw8ss9xKVCoii
vaqTLn8imjhHnLCe+f4YtluTZRITfvBlmQEaynWTRdTwvLgX7kpOaPjPuw3Y3ktLV6NZB7grDsC5
eMKwWG1/Oaxio2WcKx+MGi5sPoFilBdA559aTlokuL90G1GptfofyYMbo5XVO/PHG5kX96C/xXWE
6x+2AGSAtf8j5zKS3NMzjaEmEkrnayTicfTIYQfDxmc+GW6fD5gXUoItKJhec6knDladrgoPi4d/
wbVo13v/fdgb9QME5zLz2FK33yyOPUlJ73Pqb63/wYnOKfhighNBVy5y6SJbp9VtPeZiPhBYgV3E
DbAhzy1ENBS12vcYp/pC6KPvxhK4k93mvdnLc0Bk7FqoWbELxO04+Avih26CQgiwzZoJG3FLMNJs
wyQohqP7DWkxAt0smz79cnbh1oyCwb8O4OclYymW9T/YVKdj88fFotFRK0sjnQ33YtFoCCY4+0Db
OmGMa+PcDbRXt9e2KTPxuxi3aRED8hFvURIwa8QQTH7Tp5Mo/9MXXGHKzJcBK2MvPW9FYhSMVUgG
UaNqeCkq15EaitS8vZnPUZjmZNu4c2ZXcWj4Dty1ShkT78qyIB0EyXJSbGt/XI64FDFdfctHaEgf
IgT0KjCCr8dDmX3BvLXD/yD0MLdeMCi1Nejq8Nqqn3xFt8+EQeFc/C+rkdcXrvmKMyRV3p/dvekL
/ue8aljhgnuLLdxG+xN60YBFeDs1QqjRkzTT3heTnycSD+4hkSaVsj/5amUcycUfU8lBIjf72rBd
qOPJ9t6E9Az/qXOWIktjINhtLr/48tLg+o/63EqzNxCUMC3iK4nh5PTMHNXFmO6OxMNJ0M/7+1K7
aegfEQ65HC/mS0uIt/tBdW3YQAOyS8IxKcY/tNPqKNb9iSvzpy5qdm+vcWbTQ2Jwbc1C+QzJ3Jpd
Nh55aRwtGyTxN//vKmqBWborcLiETXEKeE9oQnJiIqFNZfZ1wiYRo/IkKnv9Lh/gfz6FN0X9JbF9
tAQW8nyB8YwNgJdsOGG8vBKWinBDYJKuXZC5O508Sd0hJaQYvQ1hwbUJNkWbyJ7DJy04PxRWgyJY
pEUd5zzQRRng/lajyIoOeVoI/s+QfyX6Duh5GAXK84vk4GXbWlDN7ecmOnmXz+FHsAVjUGn1vS0w
GBH62ttOztdbRwFhlyQOplfqQ1au9yvcRhD9cbhIvu8agbzejKyS7MmRGDUi9PgYTmrWWnQB8ylO
+dKqbAJN5PfkAFPkH7+B8Qo+YMtqCEGlXyfncBYOz55ayXF/b5stRtkXKQEMmjB3BXHSQzpcK6O8
WxoXPTyw0qEei6V48JKFjbRMnMyLK9leeEm0l2qTvn/cx9SQXCSKn8tow0Nf5q5Tq/8tIuwSlHJo
WoNDf0YNoVcveT9b2GQeU2bzH935g8ChDTp97xGziTm209ZJN2oWPb3NNibw3To1nmi3zDVAfmZx
phbfQXN479BrOIVAN4Ze/C1QoV+42kY+ixw0XDvffDaTAY5UVfSV9tgNI1Mqk1pizC+PfX97miAZ
NecWFKtbKNrpAPeYfG0Ou8JEHkrB8kB6a5uG4RQrFrGLHHayFrP4nSDgoPJhQQekmN/SwBSwGhhx
INweWruwb8FB4XjNGEbpuWf8agf/BlKz526kPj8XD/1qxuhW4v7qpZEmQa9GbVd/PbeSaFWyrsbp
2t3A8gL8Bwj4PcFTXq9zXEdLKIP/0+cohvNdm58c8o4JYi0Jq+wym6eYKpj2uz0STqnG/1dAE7m0
XDPADOr3W9UrYl6GBY008SvALWx1JKSjK1DapbM2GgFzQa1OTf1LNFq0cn6giHHiHMEIFLA8Eylj
vt6kCEsm0PWPdRmleC4Td9qQf2CwtIgafH9hL0KuKFW35QUVlxyXuZ2njoleaq19OiE9w57tYJ5W
RA/EIH7NTb3rLYWDZqNdEDZ66x0DawpL0vDaSmWMifTh3uTiz2MODplYRIMp8ySRdu3zwQPnKbjY
qmE1PasP0k+7VXuyeJXCDMUjZ16/DiMkfSNbF9X73rqgwuLzgedFmWoqne7BdfSrs8+bS5AeMrXK
6UJWbbeidMpKONLQdASjVG42Yaf6A74CEkjYCg/Fqf9TACsMBJvJAy0ep7sIb/NtoQIGlcqyq+Eb
l4CweYPbncN/uE6q4VlxOzJfz4DSqWlHJkQoGT0Zm9F4uwi7YIlSrjJNV9VZ+mEGiut94dzvKCe1
QRrl9kdidnH7unO7HB+iu8JVSx7zpCrF24c2hrE4zI7EFMvG4aDJkdSdpNz5sn/1GLObs3/UQ1/K
zhWcj8WNg4QJ216KhkKTbT8HqqRLsludO5vaE5clzlXtOswa16urzuyeaY5hsjxv8yB10MxK/jFN
GvgTMZQabxV5qCDH0UvcCHmNSCowoi8tZx1/fxfkYmRFo0Z0yS4TMf0t5tfXQSIizy6JdTw17GM/
/dLwViK4vapwqIUAHUZ92UJdAvmqcgxq94UYf/VC0R/JmU/oNXLmEqM4Yj3PmN5drCnbFfegJMUU
9rb5Yh/ooetGXBt3vmOyrVXjaPCXVPYz483/bETZCz5sAJvRk6C6g+WYlmkWkun/ecBDUGIS+FU6
pEwRSHhgaUsgz6A3pSGp3Hn0z17pl5hYIleqybZqY2UzvFbteVZh4/XSytwgNtrT10EklPsPLf1o
29yRiqgT+rJcQc3Q2HuHQfgxPgXgyC5XJ5Qsrks4rmH5KoitlDDueAv7GmJejJeEyGQHOigVlgsL
IuD1XddSOGHfQqo8cwuXwFfbEEeSGlc2xFFLrUGJjHtbuWLpqMaxVi2a33wB/tHVA3X7g0pIMpt+
AsI6Q3lzcjBID9nQhbqUxjz3iCA1u+nVy5z5PWpIngPuwwUnAY+CIP90SX4smE40mb8NfMDxgJQF
R1wlsPrPydsHjdEoeSGyjXd8BPZhEhEL3Fp4F7UBqtmVLLyKQC4HTANXOgHUmDo3MvIkNeB9d/Tz
FIhZXIR8Uxns8bMy3X9QkIs5+wXJGt093DkwSwjFRYmlwUt7HoX5eN2bn+hMveXDnJNyQs0y6HZX
wmMpEz4Bwyn8/W0ixEWpEbOFcqHTckSGjW4aK/jJTyw+aYaw0ZABxCYHjvWgLIKirzfrf8hZOk0e
d45/5Yr9Qi4MlJKTv4vWV6YsAprtk/C1MUyAg7ME5KUltr5BbsiELOY1BYQ4kw9Y4ISTOcYU6MTg
Vas0EtMkt1c/XoNAwWy6Yw6FAxdT9yOFEJjtXQIXfiNpxqyNtlof7VgBOKg+T5MpIex0H4Axklbj
akx3zAoW8TKA7x4vJhu1nk8Lbe6sZ4egPm6GK0sHNBiB2qOpBmTURxtYiAdGv41Tuyh3c0Lk8Szl
e3U4UkPObVIDwW8OvNfFvA0Wx3vm2k3LKv1wIzuB0u5tZFZubZvNU34Nm9JxqwTEJPFWVjsUhXSN
pE6BbeArupl5yPr6WpF4XsTzlIvXEdkly95uVoDLldLLFV45htwHS5qkCp0acOBmVQ8EEtDxysiZ
ilHDRb9UvlCOs8gl/T1X31U1okWNhw+YpVVPbF3a5m6gxvO0HaXyZEU3tswXc8Uc9iGNa8N54ZE6
g5TkBMTih0TqMld8OzfqRks0ckOL59YfmsAFDE9SMzK60jqAwXgb9zszOGidEmT0sTNN/CEqxWAJ
dSQB2n7RzWrqRtsxWl1tLic7UNTIkELxrCw7Bjb7SUrljhAcqJpBHoz6pqFr//j5WIsjLgvxWeEr
cMoer33Rers7H9mTe9H8thGMo0idigx4IvBmpfwnGBbrNX+K2BLBmdX1IVrMnC95bHSJLdUq+2tv
SDhM+61PtNDt0s78+laxTlvsv7ocR8JY0hYxemH78zfjrso/ID9puGl8CPgbOU2Wo1UHNidjjqP/
zuSkj/xsSVrDsNB6HFkEfu621DxxtiJPsbLPDtK/ZaEmjQ74nru5L9TDQeCc8EkwSrgijXVn/A/a
FAMNTO9GysNqxDUe6iLesxD9b1IoSdaCMMz44Y+m3c3BCN+xPXoonVlmyApXmqBXRwYpcGkevAuy
V0b4CSbdu8fQiJmKS6e+kx/xurmZOpUyBc3sU9Gq/FKVCgVEGexGX1lU2kzdgclLb/hgDfE9jw0R
UshkrWd4UMdTkK48QqinUbJ9+/aG7eX7FM8dYeWEypGLUP5rNmQv9w7uxVIRqg8rJAOPg0P9Ak+F
kIV3p/TlB6vGJg9tQyAhvd3/7mIq/AiaI0KwuWW+kv79c19yISIyUm/aVA8CbLDDuYTTX/CjcuIB
oRRzpB4XfNNiduTpufgev3tXAxRyVA9pENGe3pT5kqjlaqTtEjIotDJoAyId8s8anGc8OFsHgBF+
trQ2UzgZ5/bxk+zPfOwYVdrOS4AvcAc/XdnfNd8xrKbBoD+VvztbYS+BQOGcdavJlEvcGO4KaOWZ
+byJj4WRkJKdg3NNmSA+XduGoKaa5+1vc2IAs4R20LqzjcUBj5dIoQdhOfTbzrWgxq9Oc33yrnqU
rd1SviRJ4TT6cThBsp5z+f6315VbJjxUzG9+cNSZkQoCPfkOIPq68+/FLjN8LKEIAzzVQoaQgMFd
BpMjAnruLzfavoFVhm8BysSr0XBe/gr5sBOVtNwmNfBDIOokdgyXb1aL5SQsrq0I0ybpzW2uCQnG
joR6+HRRp1/JUBDYCRfvok5ghU+jGUQq8g4TdCFLeirMBBJXLQMP4xIwoK0xQ4r7ffETnKNs71eu
NYRBN+YUWClVRUdj95Sccno9skVOrf82gVddwaZ2wqkb3zJezti5U9wwQzLKqmd1luB/DO0ODBZ1
Fg1f1APC0I7f18JNw4q/PtrVjzVqf9hO6SJkGH2MVutOhHjsIuY+zUIpyjP+HF33GhTPb+0uYtmw
mYlPkXO5+bmENCbZxKtXN3PM11MUw6Bdt6N4EW6JXkfbI3RtYz7Y6dZ1uxK6h+oWTF/hKGR8MZ2s
AtAfpwGADmJwpHaif6UbqzuvMGEJ872SpMXBb35EaEVqwNSt44psZ7qgt8J6BTtFw0BnzqK2qML4
8GI1zjDvdxTOP6n/ItNCOXsGujFKYteEvrQL2OIFLsO0r/68jbV/e0ws4eOYI0KykiYIL+gYNOll
SsYUU3GjG59RBOGEVKDqtq5tKreNDjiA+puDyiB60cGXlRmtbJMMwakoUwHe8NuorArBmBfQjl0L
Ypq5kXoKpNEuSVJVLeoBT28pevFwp0iz05ANPoXmwLMQGsMhigVF943O0UC9Om6NJdfcIIPSxXHz
mMQp7uD/IW6cfkBX3gYwJ3nXaHXFZuHYZZ4x874KNFjNhS0QtMUgU6tHR3bT7hW4hKbX6fOxKTXK
PN8AMNvXwSpAhDM9mxIaRVHqzL0X7CXuZaB1V6Q0MMAsXfxVl1BfTG0rsQfWjWTvE2FQWgAu4ow2
Bobdr4K34HiBoKMl5c5DUiF20wQrWJn7EeEJby91ev/oIjgcdC+M0FFQViyXTpYqwFhFLQX6FFpT
nBx1JwBgUTORp9tP7YR6wE8evvxxwG0uOMI994iN7P25wKB9Y/7LzTBXwytGIi++key5jgkQxj8w
ASUI5VtIyWClpSdDWi8Zo+5DxsakQHzdAZKGYgILSBnVa7wZyNTDdqBukwEaVBM0iHjCDbQfOac9
f7DrdeSn0H/ZGKcyz2bH/30Yn5RiJfNXwG/MDDBzkJjyG+eDePtlrY81Tan3IBKZ1bI4qo+2i9v/
j7BkT4XPFyLDOjLsraa6J9uPYPbSOzLwIl8SsmTd3fVdO+i1/qsMXfrNdsPTzHyvet4hdLcKySL3
welMxH3lNnImqusgShCSlD+WGCDq2Gdr2LRylJgmP1K89nCtgmx39/pSEGYWocMJkHrh8BkecdE6
o13ymp4VE4kEKOkQbhutc+HHGcNqI7tIyN6PGYpbcEU23yzK5GX4IJGA3Y3pHcaLpnlsK3FCl8Fh
ecjsO0l3yiANUdivJGQavWQvBcUhriSvplJl+shPGhB4Rr1qz6dUx51WiI9NMb6Bt16d3jyj4Hrw
8hyDizV6LxzL0efKWZqDDf4jQS4GZb7IsZ4Cnxhf13/vbU/D7HIH/5oxObEHfqvBx0G4IO+N43ip
jyXvZ+Bvxr8uxA7vjFlDYOt48koP4EZeVHi/749lvauqnTP2HVYWO9q5WK+sBCExbQWtxqjyvU86
d1wU+tlVGvHnmazU+iV/IeMHx87as/8/vypD+PH5sDi/jT6Sa95p2bPq5ddALIZeiy+sySd96sif
jthidAoADGdcVODFkyfxXeFje3wfcfU/CP9jRtdfV2YoXtFqqxuvGupmQ+CN3vhchkZOX053/rJ8
B5ThXU91l0lltnL42dlRQjbxgydISM4qcnAtLXxKNEGrZYgnn+LKTXMNLKrpsRsq/rlupNtQERBj
E1UK8JIlVGdFHjMInMxVzAsVAoYoec0ICjhFIYtE4rPGR0h2qXgbJUaYjK2brxJNs28XIcgvXFVC
AUjMpmCw62KurJO1TUlAlsYcMZfF0+XlzHb/QjA5pXfyFOQefe8Cq6jcJro4Udgs35h4/LTpOIRf
Xs1WMxqKek/aI57F6anD4I3vB8Rh5+wL0uNtYMmwrV0jeg+il6N0moxWiVnuaUqpNgIP5dDiRTTe
nEjkIH/+gVdm2rowROrpf5ICq0K9o3s1jaCB6zXWFmWncZsfgHF42ngtHf7FG7MjoJBdiF6g7H9+
O6Tv+4lj7QzCecCb25sV9VnZwZ6yVKwYmJoWHLAoupflKDYB3DeTTZDNaOZnkNRqEbDo7rfqPNUy
MGQzTN+C5npYUEUEe70+8M/kmDR5qAnxL+rNm+a+njAS+K+11yHxm/w8IjB6HyM7D42tfo1oUyX4
LzurYsr0Xsp7Iv9mgOp9pxAzRKzuldh93gcpeoVFO3QyRgZQ9zHUjhO4A5PX8WKrmza9sccEpSyN
2Ezut73VnRIniLS38m0eszCSJyEi762X2Pk6bMmtIqwPwfOlKyPCcVklb6E/Pp9FGkmr5w8eRdud
UmRAcAk3SaB+R8qmXViOLndXCyceiWoX5ZIqEPBn6uVttdrK+JY9zi0UX+N4ZPSnHSQtGe3vWWD0
lHWG15ZYVQ+b25L2e3Bghfq8N1SmEkr1JA4A2MgzHBgr63h03yNH1FqPCPtcGgY0ikmuFpkprKOf
RIw7LsptYa60o6z9NGcX1gr44VWhvbJQCKsdQ0Tgq57ySIajuJ6o8me24E+prN66e/55st2mm01z
7s3D2tpAkwKbHcUi1xknkNC/n5Hpgx3kCeqflnz+Uj5XwH9VJrfB7SqozGxhbRwQEv8jqmuRw35/
HAduLJrcTEcXwpIUcgUBkK5YPnQcNBpCI7YjRG22oM8qW2vu+XVAwvykVzFHRTjCJwnRvVhq0VqQ
OEhTS9dWdqt91gHWz+7Xm2ek6NWY+haWc5wML1SSojBGtz93FehhGT5OcpQVgwlP+x7MLRfxYpiM
8iyP86kF+jXR+TPszM+3cd6kB05BDNH1G1ikMgz/jXrxglpEIQHuUZHTy1KnURf8h/LvBESt/B+d
qrYJGnGhRso1ZqHQjE9ohe7xPGLqPUK81nzlp2Vj7JO5TF+ZOTb83LoOZ07UMuJA134Jn9mucEem
+6vuIoa8hS+NCa4op7qN7YJQ4N7kXwLT3meOxi6mA02ZAYBlbN2uln2Ctnh/ty+pCGvaeMEnyDO8
KRPgmpg6B4haeKHLNPLf8rp+RdNXMx2zOFeXeX45Mi49VrmqbHQ6uhvIMWX3ZsH72F8/YHMbS36j
qg3FFc036xD8GGxbMynICglkP126/e0k5p80mYAbgfzrq8NDOnfGlSYa+xn59I2VZ8l7B8rR9nMF
rhqxY0459LWn5BLpMkFyBkUXZ09lt2kA5pvoX/xrk5QYFx7JJaay2VoVuvbN/rs0oa1cO8WXTVIE
3Vj9cinjoIfgLRwYpsMn/99KmXdoH7W/QJjyq5HvjOhFeaX2JXWr0DtRCqrLu6Ka0uooEXtivGP5
/+ms4wPr7BDfjaeDjSv/GDV6Ac5/aoYQIyDH7qLs92EPt3opCe0fm0hOtXLw3dTLG21+lLDiCXsN
GA1+XUrwrStUoi/+xEFYR9Ae5sC8SBc0zJE3d8+mrOo72KX199L1HyA0+jeELmEc8U7p96JY76n4
+m8tAvvfswpiUJjWYBCWmSkCf4yxW6Oju1SXMithqcpNt94ZIHqXfOWeIzQd9pDseZQMpDA+N8d7
y/U0JaKAEYEbaAlmeJAG/wTgDBMLfR5C2eo8S1EgSK2o1bE4fbaF0eTqGlwSir1K01+D3FVjWW7v
NiF3LH8oY7C1GBZ4PgNdGLhCCIVAS5BElByVQoGCBuvJ3qGyptWcxAe93Y/wkKNqlhlKf5UGpc18
GDZO2+1LMuaxZAU5dqN1rOVi7H+pl/Ocj4BnCmVeeSoBtarXitD5if3OGXekfRAgLTCHoaCXNpmG
vwviFsYD0iJNHDtC12M4qmw7HiCq5u6KGzvKS+FxZEgecd9JzFH1mnARUyW+Fe4TzE8YkA88dy6c
Zaz69GDF8U/ULEmOgnoHhaoGrhEukgOMC6LP0EcqiJyDg5jqLV5bma1spqHwoiuVB1v+ioUMu0vk
+kk35ltN+Ty/yRZlyjbpTLviDVk8DEr/vRv08Ebn6bSD10yWn7gPQdGPlL54l4ZYI7UhLz2FO5Jo
KnXjbpJjRFVV9cnqEtrq8SI4UxAIphZvjPGXeurIU9yzp78P3lE5fjzxyeh81L+zsTJp8dll/OGc
oQmTkthuEIaCzgEkCwZ5Qb8RIieyBlXy4+tkq6LoQxTauAb/aRuIxc/0mdElJjTPvQPrMWZlkX0v
Xz7ZGaEtcq3oJiUVo3M7nW2kFuCoKZ+KubQWF3N6Jw9oM17ppu7LOBaCUZjRP9DjDU7Yqknghn8w
VVVbl8kgR1E/oSQ6vORxVGFwpQ3+xFSawDTvkCprpXzUDw5FEOgnUvMTXDpAqww5U47NVf2UiniP
ceeBL2+19RxKCRzhz27PnS7KnE0HyFfW5A1n65+MpOxBipd167nw7sf74VY5+bB/5lJQXXoeo2mV
aup1LyLWzO2dauU0ps1wMTgfLbp8ucTeO46vE0F7wOapuowDItAloUwZbDt4vvlVtrv26HW0TU0v
yyWb1qJDFFrrXMdJxYAuGaYFQC3MvjsIElN+zLDqgSCBZ5kiOimpVCeyxdOC2KkVPLSChsFM8PjM
tERSuge/6Ty8Jv1BcKaszPP+4tSkrHHQU5p9/Z6zORW4GQtMcuuur0cfD/RKRym/CkI9l7BBEXNr
4mo2EKRbBsqEw2Z3YGu7FAdlUZty7VKwEHL8BgYORB3w/WezdZg1Wm+v4KL7AT+LtEkvWiP1g2PC
eh3JDTgb+/2UJeyJpe/6drnSMEEcwh0pnJxzjrWdW1WBbnKBrcp83esRb6c9menHgoi60fvq6pWL
svL0xageMgPm3OSSBXRzI4QOHn1VrUFPKlfdEKENkIA5pOA/luryYRnIb9ZS4nYTdJioOc2LtwZr
264433+lc8xKhuz5ldsL7+MWSabXSFC+3LFV+ph7uR59Z2s/qq5mULg8YsmEIJbP22syX2tq5h8l
qgb/1ctOQgqRxnRRveiPGkm4gK3Idha4PTm6qzNaQFoPGuW0Za7jEuSdkgoKs1KCuQjFx1w/EMVu
UTHY8uJqLe5+jRY9iTl/xgszf1nZj6M9lDTo7YQ89jAmzAkOqWxXPW6LF2fY+wQ6hJy/X6hCOSx0
TVD+0sVLqxAwYYnoNY2ZRcdvt+w2u4S4Ebxix+DRDDN1RL2s0Q+rUXV+E5EPw/dVq6fCySKpSe0R
2iWdz8kvQ+WbXCiDlCMZpEXYRLzKmTQVtKtmWjW0n51H8IeWHTAuCBnCdYrHx9gwNp7FwhDyt6ln
hB31pJILA1bunP+/vqqW+sUmULtAUOnRii/DGE0JFEg9iDRiMAydgFTvaw2DaKGRnlrm4DueizSi
zCtpYlD34VfdMehQ5jb07N/hymMHbM+dWAJv8P9/fnjg1Z3E1ndiUGACBqOFbiYS5dcb1lF6q40C
xnyzxuiqU12Gs9YE0MN8mBKzyPbBMj7h/t1bRmQ5e2LbC79lQ0q003uEWCSfGhUhyPjBZTaKaZFJ
TngfnBjdOG+rHZNMS3EVMC/YRVNicI441lS+gSneVknKL5YMdTn0okeFTXdhNotGYzyhFird4H97
rYC2MVRXN/15gMTzg8bWMXTeK630nbdRVF9jI1n95d7kxzSGjLuK91pe+705XqAkqPkTpBehpQ74
EJktEKzpOyLk/G3zjM/RsBGIO/6CCkTFyojuMW2lP/rq4w/6Z7nvWPiDleNkdXajFgZ1QFDG2ql6
oS+pB2wtGwCXTlZdHmbjLZ46jZeqUfMfsDHX0g7qVfJ9F+3DW6Be7fARDCv1CfzrievVuNm/uS4L
mwoZc0f6o/wbbCPlbodnsJQ6mhzxiRIeKiCu5HSesucJDodC/E9nVzbU5JtIRm90QnmXvWkpuLL5
SBRwq7xbMWCK9Rn8217NBMDJSA3H28zMsFBM75nhMjpi7clzh8l8V2qlbBaYdL6ex+6Nh9Zf/s1L
8NCJPQLcZ8oxF1ef1XF1fLP+mlaYW55Y9uh5vILn5r3dBJjVPlFHCMoGPRO6jvL5ILigyVp3Ugyr
NDDjzMnUAiv5zHX3wyKMrfehLCH0MXWuCD5YkUdaOROIbNoKvH5ZnsmuA9LHa2ZzhhOd5rGTqNIG
pYAZKi6fQQyk8gxkhnIlZcb0WXcP3NebWXHlA7uZ8njxM0AzVzHe76zIXEQbKp9nH6LuxPZBMZWr
KNiF6mHO2WSLRseC2RhILtmr3YIyiz7DwQsbyKPfzGVj/3BCuGqnnZHozfY/QtBUZkA5Cmd0U42y
tTj+Zbgkji4rG9amUZKpF6OP4Sq2UB4mIYtU9n7uO44zFFqYYJXhAeDBwdbHdsMpTfHo127UC0MU
TjoF7q6rBapmyzusYd3Xg99G2bpP4slJJVw8nMkR5uN2FAVZtBOrhOGbpZqrjE7RNuROsDyUkOQO
AO6Tdk1yw/uJ6hgKqAJHzxIUtiPqFu72/mYpcWLaPYdHfP5B2pszT8mBack4r/+RKzRKW2Mr91db
7Wg2n53cwcrdYVOtAd/XfzT9EBJed8sxRlcCqj68GCzjgP4h2M4WIbpejB3xCPYkxu5X3E+n5b8T
CCgS+t462rqY7RV85UYf+4zHz2JU9ybK9r9PupQ9fzT63imOi1iOV0dx69upSPaHEeTeAPdnLJN5
d3Sm9nWfP0O+EcpIDti+nFXz81AKcmUtyfYqG7ZrnNO7py79S4FYPGILjbLnbmFY71573MO4z6zS
8Ct4QSD2TZREKPZt+qefc/JiYM7TcyOJW/LZFUU1wV2byn3D6w1JXxV78+whq41kDrCJz6VsQ8YR
JsCY7J89UO5LnsTu8kdPnio8kdT9WyA0RBYoxOV/MaLE7ZOmmAN4ApwDk/Ja1o5kPGSXIDoYt/aT
w/3lTXFfRnHDm8DkpGzoM3EKZ3Gq1VuqW9oxmczF577QgrzPzoJqpo4tE6kh3qDvnOrL2RdO73EG
+mHLvWeE0RmhA9JdSZHCrS2fSLaY+bVOrd6J4p+C2DqI8JAqlqaQAovSrdyRBUIPUPSDIakwuvmT
cp0IL6RLMQxWE8Hz5AmWbKqOBuRipVymzWgCLKUQ9P5chlkeT47Tc1YN/+ZQ6+EyA4kY8IYmnX5h
RXofnP1VqSvpK1xD6PGprUc0grcDkY/2G8SycGaUyZ7jgGSntMF8wExqWI+3mrBFkUYqL/MocoQ+
l3EEf4npA/fAz57qpXVLQHIPNxOS5BQD4e2OCht8oQhTt6gz/uNzMMbo8QDn1clmlK9geLLKlGIJ
TpKIbloHnsBRvnD1E+aBcc35d9ZK/8tlZ8amfv/5XDQUptsiws9j86B/03keSNXdBIdLDxPu+WG3
UKX1KxrVVb5rvrF8rlRhfXwCYzfKPLsqNeCbbFYxt7vdihVZTYFcZtvo4As6a/m45X/ewWHh4Pkc
Bjk7SwSUVCjHOdRA7xvnN6A7hjtMo6rtuMvm46T07tvIhmzNTWaF4TyjV4L2BtSdvj4ALFVi3jWU
4WQhlGYWSgGp/zQRYHzFlL1l5FRbXdL0vNy++fdKlsdE5/qNO2IqYpdjBoquIkOnBv4Uu1lRaLwI
eISq+vbkJ+teLn/R74aoUEjqeW9lgCotbbTfRMRYAD0t7WdeF3crvie0wgbNFATzu00C4NPn3SKV
wGkryCu/w1tBMC076fNN+A4mllVmN75MAGBk6J2R+WNNlNsIbi8kUP7lmfDTeu7QhtretXyF1Lsm
IH7Z/Hdt7YtkIYK8rqfPGa6KxhmpYZSTi0uOGaqRFZQYbiYZ0i+2pt8JPBumqqZMkIcqFTpguhU/
YxLlyQagpNIr3KAfWBUCAs+I4bFN7QL16ulWwCSR63hPXfbTc/GuGYu3vbawUBtAkKcREezCyeOh
K7CAkpykSrL4V1XbG89flsuOn06yfjAJa36w2gZcnsEDgl3Em4W0hrsUdBsuwOheVpD3vpEoavGH
26bypghlvxWFylHxFWKdyvnYI3CR4mMfRCpCSUXHmy9gnAhFLuGPFQWLXZI7PErdvCktyKW7+2r0
OSuFRIr8pTm1ETpzNt88CSwPBOssQjTYQw2/8LRLjHTBtoyHOqDCtZoHIxA7Hb1Z48NWI0iFdFHw
XP22Ir/mxxXcy8SbCL5zkKal7QH8F++tX+TILFfxp2eMfOASU3Q/QJ0sW2vB7OimXjTBhj6rW33f
vbUaIWAv0MV0yehlOVJgT1VKkNXLAEqMBvCqnSKmY6weOVorPjm38iuudAZf07PFE7TMQUXVt5aj
YT5tIAxM4+xtdEzY+au6n2J/FHBUfsC5FlBDAw/64Wgvk0Py2G87lpmOzk/YQUp2RFyY1tDMBafI
Z8t+BfHJMvVS5TmofMhn7g3Xr2klP2dyp82WvJzKSvu8vsu0tjsEyXA1LCKcOVM79tV9UeirgLQE
GmVa4E8yDwbeuWSZIWOczNC2Ig2tLq8F5xLjhJ5K6M31fNWzI7EDS7/O8zI15/LF2wncMlYJDsvg
hNtL37E1boWl0l5amb7gijo8nVRd3qKWTa7zLLyq+J71ux76pLoz13f4GS2f7rT9cY776ZmoJWkj
UrFvdhJUilJeZ22MKENIy4fuPheK8v24sUnAK/ghz1OqvdW1vlnwcMcAD3F18c9AsTF+sOBPiXx5
nWy4d0/Do4YcTxiV5wsSs2B8V05ZNt/l+FQ3Vh8P2CvkssT4kssMBQfajuEuQC5y29xd/T0lDavK
5h/FxwpMQYO+RFh6kh5b9B5qA8UNs80ljPH4EriEdh1xqPyGKN/SzC27F+D10pvQQ2ViRP6f9M8j
bMsLV/VEEnL5UVR/2txkIB5K75NqQzOCpvFKyXKGWFDPuPpLlFPoje4UftObjuJUeUrslSd89c4q
bujCpGpS0nSx+S6+wmmHZ/+Qo6YTtrDkvnPZlkDylB4atvgStGkzPdnPG0LmYNgDz8Jfenz/tIIk
NdabzGO3AAt8djmt+p2Cf1JQrM4wcBiDFI6fYtFi2yj/SRbGxiEIk1RVB6G99BbcVdbZGlh5J+CC
txj00d177pPkF6C8HpTERHmzOT7InHKy2zqERShgktZ/M/Aw4ipTncxyiDFm/YZsOW1NECSLPtuR
rbPOGwVq/15+y502fRnMMIS6we1FscObLTSBDbNRYAAx9gJ9wTehDsgw4atOTmNVYkDAfAnumZK1
RwarjpPgImtL3+kO9K/qI3V0pMXIoABW0wCg/IMks4mH1cyyAPrph0EkxfQ966W6+SlK5eIPbc2e
4iI+XkwCsEIe8Y3qD1HvKW2/F013g9r0QjSuOr3qrzBKErsHXRy420bkAospJ1o9mO/lJ4mpqxSJ
sAAkXUYldtAbbDwcxYpzNpShy3TYMlsCrLW3Fq3FtVFGjlpeczCmhZgGetTF86C0rBOwRWWmHGPf
AQcfNsyH9SyEe0hCp4N4lUVit9Omp74Mr9rDNDZ4f9C2T1KTZ9pSqj782KKGTMQfEnT6Pk2nej3S
fjNBTe4hoJ7xdSrgiy7MjJobKLuPI9ffuERa9hVKvtc6Nyu3/v7hxUDMgN1yCXNxTnNH9z7YVWpu
qwGg2CMz4w07ejHTZwTdvZLsZkrY+E5Qh/mVTnymj8FcqYEAo7/2y6mC5JPtdkHmSK/0XFGqjZgi
F1D0LD0EqLUanRDplIGTG7CoNR4ELYXTJovqXG2hHNDtT2HsMRz39ZGoZh0kaKbVdRuLsz5eL6PK
E7UGB6V4K/7XGkoU/GP5V/fgrG9TSKQSECkkpKEnletIu5TAUN752eHY/giSRNfv35rkR1NwH1Sh
g146xvXN8StV9/k5yIdJB+2tf2abrsHYOPymQSKb3+kT+GqPui45Rnr5X/oN8b//ySs5nM8QXi4K
lQjUbgBW7oAgWn+wiYK62jyzMDJyr7CXsmCUq7bUWUpmkBYw/UaFN+94SsEGvLEeY+SK3HVKdjB6
xYFTyzUsxLWUHm0O2Ub3gEncq1MEX0nvTWboj0WWyhiUyq6TNHIChB4b428edtGl7GDVTLWyQuvn
tfQfYCnieU9v28GoXgCKkb9o67RFIW1GfGJEkZTb3TmgepY+wGSq/65z75IZf59PtBtb85+0yXYc
r1TozBjglYI3YQZV6nQPq6kKjhtNCZu/GqHEPUn4Eq9PK5UKayEsbT+gHGUK8d06u4Mpnv/xA+yY
YybwJTzDanUX488DYd+sq2JR6apC3fXtewxQPkX0hzmbVq0PD3PDWmPtK46ue/zZNhtIbGGLv2ib
FffdJoTnwZJ071Eg2cyXQ9HQBLE21i7iDUrlHbKNsCCv3JjRfPmWlnsGrXXWoaqfhKQPe8y4Cp5I
ZoPt/p69eshanHvSYGymL9M+ZHwNW40BQ4yKHnyestBzxEeoaQcy5tuoompOMW+6IgIrF32WP0Bu
1SSTdPD/1wHfdon7plhATw/E7SlKZxGSlq/Dzw/UcaANXkFr4ACCoOu61exKNu6OotEfvc77Rmen
a20KLFfkRVSwmFoUdKegRSBsBYN3djYebTO9GZuqlEe1fHVqVNtiZSzxAwwXbNOfMSZISa/kR5np
K6iRKGlxChNF/BFtIFZCtwXDuk8mVExdoqrJXQqbYYjujcAr9dF8hz8pUUeOePD5KVmhWEIX6+P4
O1CWI8c0LFF79irFyQV7o7hWXm3S9BqMX9aXIeBdbcfUQHdSaMYIy3LXRgBHCYyOQYEqh+EiYf5o
avBwN3VvXWdrGgTnJtgJhcWowvCkaQj7mddyvahNSD410Nor9589ufSsO2j6qYD+0FPNhAnE8VhC
DsFXhjlPz1Hq06Ish9SqQsFMk3wAS6Sg82jtgdKMPC3GKuHs1m2AiZSVgZsAOZ+MM7RUyXA7T1xS
kktU2Oho23AL3bL1pVmqqr+KxMV3tLnBTEC+9vaLcdYThvWpv7PTlxGAr1bVt/bzOEGUSAhslxja
jOJy6WFJzIEZfeQ1CEcZpHzbafLFFd/SQAlXwaIlmDKAFPQQryZ399y8VYCyh5gssVQL37xJlrfP
4DV27BuuI+Hzaya1g6Iy9N6lzNWsJ6fqWWbo9tHv/zAyeiWGujU7SxMgvIiL3TyvsSUOoYs261cK
qO810lczWHQG693stNTHAqyfpRjVUJGeQcEcUE0xNnX/qqI/XAnxTOeQrUjapDlegCdjIHad2TNG
yzg5gkqVmTy+cizkmqhlzk49mvg3giPUOalXzqsfYy3T/XsL2SGo86ebiE9/f7lF9azuW4UTu9GI
bJLAIS5whIvh4nDKF7J4JQ6fxP5sMXBgVP8Bme5YjgQpJdUbEkWb9RW21yfWpds1pCpd+iKUqdV+
zxPquZCdlqGY3xBvuuKgd+Ob1UJG5iUFqkgEJ08fFuJB5JxllNelbpTKXB4c2RJ+CuVhv0H0a3tl
X4bLw6XURQpiEFPytVYg/+NN+iZiHM0RZa+6c4eR1PyZKeqZMzzDxBZ1J+0tsDIITQj/qgSkf3Wg
/mGBn1VgbbrTZ+ELM4IN5aO3YQo1L9WuyJd26CoH1wxuyr/46UMXpNkzNGKbulW4AVMqNqRO1mGV
wQ4l2tG9UtCaV9GvvJ5KfnGJ0Rowa2cJ37+zQqAfYb8Wl9xhClWbSzRuwZvMweeSz3uf/M/SquHD
LJ95WhjVKUUEJmXliC8OfhFxl2DIQlYYziGMKeLI64MoVY8JifFXypahIImKu2LPihPQ5hMqIwgR
uCFG1t5HGdaAdq73LZpwlDNA/vMyi6vukzdDG/2TOfuxsc28N5McDqeuCnks+Dw6L03yo5wsj0en
gpoOA0cEptapRtkDC3LGWSQOo/eCAsXnKVFM8zzNGDMSG4b2Crv8y78i85OiIHqr1f0D2uoKEHXy
u6VbgL9YiHZ2LU+s/YMbRWVfvGjAnfOibNjIh8rtLipqCEKFbm+LvESTyf64nDOgRdNOdbuWUu3K
L74cQI5XHl0hwEKohtpnqw3h0ycRX+neBVrU1f3xi85z/Pinfms89jNhy+SUCqzPniC3f0+N2NUO
aEmdT+WL6ScLETVEIiKl5SUYn4il8c5jkN6pxEwZ5Tx3y47w0WA4D7yyBWGZVIXAxsVBUANsJLQy
tqJdpkOKz69TJA+J/0LcaiKgL2ohOFKrLMH1xZG/1i79MaiIuAhIcsA4wP/7zev0TkTSFX1G/NwQ
jHlLJ/etHhaV1OvB/1z+skSh0H79JCrFDPs1Rykx2J0OXCg2UKlk3/pHQ+t+OdBUxqvwERg0KsjW
rbq2k30Y/BHKk7ResEMXxLgRMi1BE0zuy19ep1p/GGG/tDgfj7u0BR0U/p2gbZ9+h+vOgPo6QGX8
++0k/LYwfJ0a6BkluSdL4eTt5RAdz6LGHF+J5MuvrV/xMHaEajyfnTfoGeZtSOpUF4YTjTqYtgY8
Koc2afZeyT/RwFgziJgYLVmILrRj8mPZjxFmHm2Ee0+WwKuG1p6v0YDhvmPFXygm3qwT0uDFNalK
QTrtsknyVaE80w+snnK5PQgtGww93iDVyzjUkoMCUXcjhsD/87z9VYtrZVzItpHjqV47MoVOfKsr
U2HH/zR70Ms3VB6uH1+3IAjP0Aa36rX/rVZUxr7FEThX+GUEzdKXfvNDPxMXSjGF+VUC1OljDe2x
1i6eaQ2I8T8ekq693q7NkozqmF8EZRn5p74EQ/wpxTFPzQs34cN8SQTyyQFQvrRDEq+mVCz2dwg7
nQQJnsB15MQllUErbFWazRzO5BbUnWMPOH+Vyz582DSVRMuiciABSgMBE8RVtFa2GykKv4JvusFS
Iu5lm0TV8IJ2O7zSwwBNxQ7VsKeJcBZuHTC12m3C6oKJ3vSdayx3R6bNKcvP7bVtOzp83m7jMa1l
5n5EntOeEMYeW13yK0Gy/LDiYjJgnUInYLCA5pxKkYolz77Vzk6a3MrMAVCUm7ln+CPhGCjpKLwb
HfwPOJxollZimZZkung8YkIZ7qq1rqyVLhB9dYdc/lHx2rH4wgykyCnSCst0h1E98ThfVwPbpWJS
+doGRNjsMOZXK4UP4+Ai68wT/IZyi70j7gTRM15DSCPiHTU/R9D6yv563wnpURA0HkuDnVphK3SQ
Z27AJojpZGHPvous5hCD1AZFhKlSRwAD3ePqI2OFURiouU4zJmCxJIBohwwkcjY1NqVkm1avUwpP
CGgbFekt4DdvLYJkMogn276n9nTUXCmRDm+DDk7IO5+bWrvbgUAsB5xyz32y0YZfmCImfEEEAw7C
OhSVQcIHGImv0AyeaR6pgZcB8mq2RiY9Qzcmyx9hWkoKy0kCNb9frgcNFUx1ksvGRQmgGXzy80B9
6m8WHy9P6JcLe0xvvnAJV4Hu0oX6HuSjvsj1acTPYB6AYXhQuFKCuyDcW5iEElYnD8Wdk9uPAmkt
3QIrRso0/T5o9aKHsxmMZokgtgX+zzbPHV9/FAgDisLVeRcWHgPoVZ2oiXlBX10GjYRkKt3hLkVz
cXm5vcmLGhF+smZPAKGz7tbW+Yx6trBeuzqLy8JE2+WzCat7nEtyh1pEkC3c0qpVN/NgwJ62eN3s
Wr26wE0zXx06U4Gd5TndQXk/5ZDWE32JDpwE0ivXwm7rgOexFkxd6GDbHbYty50mJ46PanfeOlZU
p5Z5OwrCkh9XAvM9xUjuZR5xFnzOydegQ/3Ss4HRwi0H0ZCxSC5A2LRAFY38JlJ8Vqy8NMV0JxrP
UPWGoHJM/90AJyyzqjTnuiQeH9idkq8KBB0c0aiHTqYyKTKD8pda5Sdb8bLoMH8ejodcvjHaiUBs
w8j/rz9AeOfP7v+UClZkqOlQFRwlZS6n7L4zD1iy7noCUsxiLOY8LRywOjVdLye+Af+fIuahR28l
wVnd3T/4s5+kYAr/9M8yEsorkaWnUl/y4BwH1XtN9ElHe3SrU34ULY7GRIyL6x54xFqMdiCmitfu
yJWx6BZUczc0pgRNTy66YpXbML9chzNdAiPXi5iM0QkSRsYAPhnbd3lA7cwwr121o2CPlmBuk2/l
ycOdKq7a458ofMvi3GAB2baa70GiPImn6ftpj1Joajd3wC82Q+cbJK+fT1TX4G3DHXPWrsMlU7ai
UJPyEHL+/5VLi/lt35MMgUMkzD1qQp0c/CNPKacW/mHXAYxbUOhPtGMxtdwFdd+UGPmDGQGJdvBo
qGvdJw5xvXb8OCvWG9mWcm1bKYrAOeJpLWKpRi9RORc0cToUR1MI5EncLIZUmWUOifkeq3MQGSEo
nBoTkE+TawFJ1Y/P3jxL/OBIwmY/s1aYLgrSgHbH4kCG/2G5mEKjneJ2Zqd0MIP+bWdJFeUXCajc
zAODvZ2ShJLPcH0iRFXQJYRRBtn5CmZOf+rtDm7hNobuYMwSKgh0EDb0BVOmFx35r+n19v+Bd+YV
NbVUiFYvFXAshi39M0890G2WcAHbxw+9eGnX+NzUD7YAlobWyHtHFJLC6wdxYq2Km1aYmw3deRSI
kZTDGpr/ueyaESuZoFABccfEkhxYB0B13bo0oY0swn7Wjjze6NiYGcwnxAPHgc/EVGTh+7807IfU
wcF+A/NvEb+kCVCveeAxChkX/p6ZBDpsq7WiiBj/i1Gw4rpinbs+Zqtwo6SFdA8aK0V3p6T1eMMm
UKQ2HOgcOHcVntUuwwMUvB/jQVf2VkJgxpNriEbtogBmpZijxLU7MQbfnAZcipXSjEP3MCFC3s+S
BV/hfFgOKkXKRFVINLwntrPbnAzgRbH0HRNo/O+1wbeVGnPMPzBTcXbZyLCtOnKUCHj9rjWxtsJl
tWwls8g41o5O6XZb0IwuO92KJFcj6QiZyDVjJAD4W4B5RdFKN9+Rnkv7BexrqG3EIX21Kb+SGy2G
p7N4LAd20oJTEMLOxTbXZjVP5KH7c6Svn9HCfU5xLSUWK6cPE7VKJksNqtAnt0OKk1zWihDKK0Sj
kUftU4gTdnxBbAtMY1x7Yg03GGRlUoE7KSjYrs2znqKV5ZkUlk2iPGjTE/5A7haH75Ce9Wkhkn1v
k4MSyYebZMTLV93pxsnaKWWeH47Z3jZChXjF9otRnxs0b5sVJ3SH0OsimynLYSrtfF+/JnzMLmc0
mao+GbyTcCR6UNfl/zD+Kr762u9n4yZlNwEs8BSC/6b5c2DYeNEKRdIXPCERxoXG/5dJCCxb3Lum
5XZbXovQgawC3LkCPp6hFKXBLF5JN3pF+ah2T0smzeibsACBE+kgfVxojFlYQP50PStM0g2WnZR+
nYE2J/2cvMga1SNCjX7qJ/8aqGD6OARkaLA/NlYEbIpV3PGiqbAn0OC12eKUl/JT6UoiLKXzwk3v
/xXeLhIqQ1A9b713otufm5Sy38X30ISaYgHNjyVLflhTqDXNxZDYaOAnZvpJoS70pIQr2SiwU/In
ackcTeHAwdFH48hqpwLha8rSxR2U4MX+oWP9iuK1ia9jEUr2NBihzGIYRdSuH46CfCAR7r/6Bj7L
Oj7Gkbv2MOnpsX3YXP7j7SLJt5KZaFDlOpl+ElzuK2FLl3ko2ZN4MosJHqRhH2PCz7M5u521yRZN
6vnB9P1LshaLP/NckzHbMokd/K65zexdqCoY0LJqoLIIKXdmy6RIJhMpIp9+jn35ySB+FL7sHq8i
VVCHjA1ulpLPd+B7XMSnIQKlRn9rpyjbvpd0oKYPIuq7mBOxKaztbtDZZmYHlVtXE3TdsW/lMbzB
eDDp065tQ4dpQzZGO62e8Cv8+W5uq6CwhT1t457tB7y7fXYDYEKtaqKU6A876miGUEA8QmymCh/J
O9cY4fR1629S+6oUbT2Jk1J4Z+wRu8VV/GZL15GSGNVf8t/AGXftKswUZGukWbqqk91W73WJeAiH
F5s2Tqfe6jfP04DAMq41d63TBzmYqbN6vzwc/BimZpHZvwXVkMWR8uJjmeKo3dW2ttuEcDit3OGI
Q+R8MmXVVc3ASKAmtncsvGn5RvRNu8aTrBbnrwj9o7xENL/aVp0lAsat2KAq7gVo19kmji+Rdz3F
r1np/rqgJmIT0372Ua5YCM10VTw7wiUa/G4p2Tx9hn/AVzOdUqqWIW3dIi3Q0aZd1lDDv8KQQfVI
MTymk+l/GQPavUCzPRlYkcDr1QQfZWF+5cWm8IfJZcJ01E3py2KohZkMBjeftrQ306dgf3n9h0kK
Cb989oTgudYBtSItzA6YAonjMEyjV/xT4R3yFsv4DX/i9jowqQudfggCfbEug+c3xinzBonZ+Wf2
DF8tweAfE3VmRYgjybLE7GzDNu8xR1IMB7T1Gqw+ZK89JbhJdvl0XwpDxy5b2xbrZYuRvG6eB42i
+CymBLY40f6CukCC3yhWqBjQGrtEXddh5Uvpfx2E0pTIVGkrVox1WT8lbbO0uyXeF/7JbmFEaa07
esihnBS5V81TtjXyPTmWRU3N3663VhbpQxUu4DXQOyFdmsJm4j0lG7CuY2weIky3kb6gxMXkNrtK
t9nyHP4J/cjXptTVk8vb5GFUUc1sZ+DEfAfk2fWIix/V8BSl2LphQjxgrIZbRQrmd3xRTHk1jrk8
kTiJ06xHrMnQhDII9AsYfslEcRTykSGQvNxPcUPEciIEA/Jz1XvPcl78uM8AMupfAA3DjVaoWA78
L0R75lQyUMrd4UNiSfBSCx+7iCOSQP8d3pBtfqly7tVDpFfmdfEwI5jyJRQurMZHCItSvOJuBIcj
ygqStC5pwrWyBxXrrASJuLCh4cCFBxXebfu7zz0MKvlccxRHuypfCyXFz/v2J5PKp6b8LajK+0ga
3TPnDBH+Yq7qFZvkVVzofxwCERIJ6KzpxHaesQUCzP5SxN9WxWt7+CAYOJvNC4UWXo1Jc4fbE2u7
D1V+njiMp6gLMR+ZoP4WWuEjlLLllPVl2GJg+pep/uXhtXWYImMuvg48kWGcPdK9C2KxHXkGqkpC
XuOAAuK88k7hH00FzbSUdLgYamzDWp63sWKOZQaICrWN2bbAPFoCk5KE+Sbp0rBr2VojaT9mXuSM
W3i5BnsZ70zLWN0U+O9P5HJOmBIBH701x1dkbuTm1oeFZcOrFtIL4JVewDo2wUsuQnKtcmbtiRml
QwxNAbVgMGFFHfi0yzFdLbQfa6Gk+KRBb7Q5yhfnf87Old0tJYSlzuzh23pUD0DmDvUPizHHlzPe
MV3zMNuq+YJBvHY3kjZe7E9uymvsO/0Wzz4evEZeA+/LWiNBhZeko4jar9Scb9m8Dc/0mrLjHoaF
7PWcZIlVIjDNqVGRQ1jzHkUbaLvDIaNXUt7kodWU6M5jkJWDyUl7w01hrC4ulDBSkbnj6bMPLlOx
kcVZ9PO3lPG9RQnh9xUgv/nUvKz5fn2vR5BkgFeyACfXMfK0KrSYBKacBTGL/EsAOgvjGM/k50Kk
Mihmbyynyz2Ewanzh49QCLIS8XTkHgzSOAR6/Od9QTZYiLcabRTZLBqf4uVvvFmqz4pU6ZCcXQOX
4YXM/ugnplkvotz7DBDbSp9BF3UuuwE0PR80tFkpvBOIJyFyrYWmQeCOZ96QCcN0R7Sw/vR3Zgfu
kDhGoS6vdjAsi/XLGd5euHs3gdWILRDOrhVx89CK6tfeLMNoSRzIFHjTyWLM685tY/pKenrEI7/w
y69V+4lM73O4QTl/l9ayu38QqE5hhMABRJ0YFAFSHGfFOuo8i9o9h/hsqbxUH2dCO2DzbU3HYdtm
hE3ce8Uk4fF4ubkC26lbzc2DMGii1GV92zV4MFCHxpMu0Sv7LkTqeXGJ7axrgjbzxTw3OePlRcAi
QjnvQXSvp9UvqqYKDsmUWtKa3kzkt8JxZgTZl27mW5w4NYzjXWHPO7PDOSgnY0yi2kGJFqqUGeAO
7fMDhZjDpW5by2wOgrqqdtSlYlvubNauliK60cOE+vtznH+7u7Cs41yGnVEFEJVzLZhwwlKUt2Ko
ChDfvCboXCg64XMdw5uL0auedKwmYcgW/JEcbJQsRUGLW1r2KaiU+5bGBoP0VdWtVkPHkLqzSzNM
D2/KFngHVABfSs17i4SftNwtw0NLAR7Aowy9Gc49+COK1iuyXbut7azRt+DEHJu0dgqNfxsi58oS
EsB/zKPEp17ismDZw5LtjMjAewvrLKDXk0aHJ0I0xDvQCmFQfm4/vq5+QmF8VC46bI3oSKqEVa17
GVo7duBR52Ij/oPSp2C/si5KXI70DkH6LF00LFp4xU5NnyxtpCYVlutw9Aq9JeGhW8LeVTmEUFgU
881UjKxGG7btcvmN6ONCV6H0YXx7gZGctyVGGv1XwC9icWv/iRXyJWSH0psVmAorNFrXAt5R/qjR
3vRvhvaT0cmViQvRvbfX8m/OiGpAWfiDpVELI7+4mi+grTMW/iBMq4d5KZnFaS7c5Nhiy+S8ihHI
8kUG5JQLzD/jk09SuyWBeMS5XRNLJYc7xPwugErJOUWp18ndGmHJUL9DQG/t9qB4Aphd6NJXDtlS
JmGuOJHYGk7rWKSX4B2T0eMXsUZT3AqPLlLCrPP0vXJwhoZR3Hzh21eCvSLO9F7OkkBji3PS2uXK
zn1xqtH2FFIVYHd8oGlBHCEER3LGyKJGWAMyujq6w/ITQkCb3A5iHcAp6wKj24wjEZ2k028T0gP5
hqPVMoiN1WZjGZg0xodm3lnvp/i4Jhd4rv44mpdY1QP/VWIdKJoL9zQPM1gxkXavFRkF1kD8oC5S
QTgby9+P6pPdz6Wc6DgeV04QExIH59POCwWd3lqh67vMbk6pXk9nOAlCKosP1vVfmHnByp8Sspjs
KEdGp4Hv2f/ndqBt9/tIyUp517afZulMnRLYap7JwDhBbN19QaRs8LqdPazZS48FaE+q9bccrhcJ
6XpLmHTQCOfA958JRBgBdjX3DHQbp5+YhE1VxS5dEELsoWQGsFySE5/w3/AMjacr5//3iibaYLBF
+VkNlD/2fuLJ0mB/1hvlyVnLXNzIqmKNyEF91blExCscnp1yFv9zMXzO7arPB+RXqW7nsVGu8MfG
IS02YtvgqyPiXWeKfAHzmmO/s18J4h9TyyJnP/n4LDL8xFjeIBu6YOGqQ9yIXtMlQb4HG7h3hYgP
deafsiWj04lF+hMc+7sffCMGM2tc77RM/v/cM1EC2FgdSqokVx5tyJfZfOEFO94dO1cdggpmwTel
ULC+Egj1uQclEhgpXNDOWSg3Kyrb4pObfAGjtsjqHO8s+Zl6mrUCZJISvL5FKaM6sxcK7MrYmhUm
7ta1hWFWxYi0pTzGLQXFFiEJaYBL6h5+uZHIzS7sBCvOflwAJXiCqeyILw31jKYEc4llBHnDntWy
2UyoTGXyof1TOT0a4iNh5XT6RM00ZFkm9WcKTyi6kNHUFf5Bfs9an28SdLQruUbsO7juB7q42bCw
inIHavjB7SisCZnKRSBQskXQtel1iMOtYiBg9IN1uRTFsPeL1KLZa8Yi7PKRpqIkahuuRedPVFk6
tRR95TmbCDOCBB3rwKeCiUL8fOXod5Wy1DnRcCogc7AOu+IF+HjYsdK3hI0SBKB6+Peia0J7apCz
6C+aYzAkKDrfUGQNtqLZ5vC7OlNhfumzgMoe5LbMjnivs8E+5glUzOyXl3lzahwIs3MdBZjb0lk8
WsNkv8BwvDZQ5wo4qSHj+mKfveHONCT2VcKPbXIHgM9L7rENO3aij1pfYSPo8JpzS101ZoU3sPmm
uaQPWWO2pvKN+UR4HZSTDR6C64S3UysngSsXXopl0MbNNll1Q9uBRdufVHw9ypYK9dOqSCJwIwPs
oB/VlofZzANf5qCgSoeO62ol4KtBEwfsiOvSquhmFBRotMcaBxoxHrxxczXumExazsWd7kUTGBTt
7HmSNRVzKwQe5bFKeAGXHIJBHUQCZN6UxayooIUqhmorlAHdyzW7RBj7sMHEoqoHuomhNuSuJwkN
ab6VAZE4qKSHDhznTHNMXOjmrclW6+cRoWg7ssnpFd699ehyMTBd6bmEcO+1Ipsea+Bt7XEugETo
GtEPR0rtyH66sOt7k7eNrYZItnVj5U4bfypgmhF0uXp6BiXwYpkHoysGQTsSwRsbx0/WDy/CbRIx
UrH2WQCyFjnTNsSdByVKHdESDJ8vw9bNuT2+iFn6cubfMnRTQLGoY60T7ONwUlRkeoMHxRSnhYpH
/diwJ0vUYt35Rew5SVNHJA5eybDIF58vFu1P7rileTaLv4CRrSMFb7UkzXVPaOdCXvqC229urH5N
PpKcMZcBvIPj9KdA12KQhodwmOMBRJ2xpHbIblH4FgzSOCQOKU16VAhJxR34jXRN0bBK1itXwR6T
BMRZPLG2Fj57FHkjya4XIJXAS1zKyWqJrsNud8rP8HonJrf1ZJNMY3k7E7Pjsh0ScP0MW6ch1zPL
lfP90PayRSy4QuOc7PU/YZX7BgdnG3A3Sjii5EdwUe8vsFL96eAN73pVjl0njQZvbqEPKQDHYeY6
I632BFxYprxwHZ5pTXU6VWpHFZlXXM0UP76QeK/2hkeONyHamKmxRFZWw+kSz2i2jV6S29IqvQmQ
m4Nt+DRsU2BBJREqqKc8VAMTq4zY0S5t8ISfBo1QACImfzk6WgXvTf3qxlSLZOoUG3CilmTQTDqw
sakhXMXDBSLBvpyTc6KVznbax3LsAzjAHZRy6TrPHnIZCcH6aD/fgrCZx392bb0OtOSU2IGl9iMR
71IQKxipR+ochyzo8PWqkzUPRdU8pSjQ0B0lHqWoH0aEN6xsM1PYdJRzd4Q+EqluF0cr5PAonqw/
NVdrbyKpc4yRTCTIudBedDrRKHiaRkQHECfyYe53KJmes/mqaxs7NbqFthoghDZ9+fBv6oNseoAp
u5lY+Q4anJJRIupqkxOV86stRqL4ZfmsB4vguMcS1Ma7xXxs7Jun+f3g+xJNnGjAXX3NZ4zS4OSZ
I1V8BlIOoFMntXevqcZOPr4nGcwumsdkuT4eari60sAc1WXdk/1sU9pCGR1WGVEVVZF8qlaFeK8e
0szyBd48IqeGL2nIFVQfRq7jnYePm+a+iaNoz/csUKNwWp0j+4JR5c2u4dYh3b2j5F3EcEQ73Ljh
roFUwzko26l890oZVstEMZ9P1hnVarYnusNh8m0nDhxZCh+3pEf01Nu88cp0GeZRPDOtJJ1kZtpZ
MRwbcckmE+cyEWcSbESmSNN4OYUyF99K7xntuCS7Exo45VYtjufdGQG92sl5iIQP8nwPE1u7AYSO
g0Tg3N7b+8N5EJSt0IxD6wNFaLIJmjuWYf2k0VxDcQdHWmUmTyUEx8395bw84Pox3u93EXnk0+bw
Ly0G+RMDwGJHYX4ZbqHuqaONaZt/uSmrAHfdXgCy+LoOcRUGOYtE+xu4WJCbANbkk9F5J+HsGg5C
G1/GaigSKhIgtSgU60cH5iV1bp/pahC/v8t6A1+FuJDZB2TsOie1V7UaH/00LXtj+nHFQw/ZLN6h
96fmdw7/JC/NOjU0eswjOWqXJOKSoWUfFfQEGco7at7SYcKI8LPiOQJwnONyvHPfbSW8xNnkiwtP
gS3ULtoWeQxjCYfwkOVf7ZMdUSWToBVIlaM2Xufewmc8qk9aqHRgNk8zMMPupbUfS4DcJEN4+JU5
Lgm6JjO6ctuOK6cBdgnAKiGgxxa+wxcvckTHfMT9T5+0MeG3LSTLiDXt0mdAGQQFwPdPQiVQGQZA
9sAsZvdiELZWpJBOtpYXCGdYnPCIQUSevh6ma4aPjGWwIcCSanWONnqxKoDobxeBPZnWgVCv0yM9
7Vu7psxu3OvgKKC86Y2q0G45mlLKtUnf2YnJgd8ErcetYyfWszWw0yE2EDarbz1AiRd+7/41RZHU
tmOyTVP6yUBDwzn8cdFsHV7wZmdAYHoeZqQiKo5Ayg0dN+/+FBSMa/9UyfDJGrFNGC9eUhcqNrbu
1/p9G6uAht69voiT3v6E90BG8CfJGLGeKBRBOH5faHzjmRJJUxo2vaaR3Rv3CUj5iP6pCFG+eYmX
bHqGNRxjTp5pZW3jUYWw0Kunfi1t9gpMoZtINvTv6s0Qz9q40yc83lnon0DQWXQg2P017znqXvPA
+F29E7yAWae8/2a2KGeEhrcxQ/X0C9b+n1WW6Mnt5ZPdNbzopwJgSbZPS0eoljRWy4w0TVm5FKCJ
yYzCFuNOA8m/n6pEN8debKBO/BIlAeQrO42q7Yx++KRNJKfZCT9Qwny6JhjbRWzxe7dVGpsWK0KS
bia+KGuCQvOx4dcN/0oQnc1A1BWiIF7meDZMR68Q+VGX3UuwvgwvZl7or+M7N2CXCq8wYuE1kTQW
H5p8m9dbDppHs4pGuz2iDxcbnlTdxGbI9scDBrUxRgBT5MedWGexh6ZBXKEwav7D4Idy/sAvuDzT
237JEWTYOJsKybYeMUFHRmXUQqD+Eh3umRrutaguI5b1OdajiQDVCEUNtMzeBYf3rW5IjqLzxRNm
z/WtZXmMDwgro/yd7pEB9TsIhke5tzxG0T/CmHiVgE+EclLGqZwIhjtcQoqz5+VTJmNfjkBxcf1i
epzO2cmhPjuj0znFqcNnhcF+qd5Hrw1jWpzo117Aq1J0DBFnAFm8h8dqZBT9t8gz5NhnHR6oDyUj
vno23s8UFaHmFbW94nUTT+LVSnPQGlQXWZaEFJDbdr1MY32DX8cjTLhyEyFBZoF0ZJi71Oz1k8RR
8Xk7VxAAYpLubkRV+6JfXfWWmBTxtgSxOvPsrFYNEqat/VeNfwlPyHJm7B5i/7lA8wdUQSbeUEsY
3z5fElaGAooI0+Cq9g5kFk/k+TkQNBFlDwrB5mqzvmT5u8mO5RpQRYdzEWc2zj2rMzVzslFUc07e
XFxvbAV1tks1QjlfsHaYSRN5QmoA2Sa0SjpGCt9qNH881yqC/GZjag8MnN3HzK27cD91Vxk/9m+v
Q1+tA7pzIBsEHhpAKUOPatOTxcoTk5e8Iqx07unTd7NMLDJ9DYNAUwjUcdV6A7GM/VicKvIFOQRS
fEoMaKXIovEFI/EQrxQN82DNhfXXmolddUpTCuhJKi8NaOL02Djcxu9VgRP/Ix8YNAJ52HQv9+Nn
q8qeSIIue66PxA72O/vfM4Mrp8W94s/QPO48fZ0e0BWfbA0kMk6Jy1q6IJjMpIDmgAGZj76F97+6
SvQSbALdOcnfktl0PZ+msVyr7TJSymTf6dcKYwb4zZgppAR1RVtWIvA1TEW7XyWMinpSmbxJPcYX
QPaUoVFt2B8kJbUq1Ytoo2lD1jiJRGoBm7Iz9Vgw7zPjENFbnhHr/HPCYbEQa2VOvnu7xmQtozaE
Mtq9SYjDdTMuOzupzAl6xMX8L1DDWrDiZ2wPjL7z61tGGIfyoLzRIiXHxRD93MAdI8T0oGMCGWlE
49YJWvWr+sxxr9TBUT3SdmqQVfuusfSIpCkdDVtx3IdgTVtb6V89CDKGRjvMuE3hFydUYBGmjOcH
EyIlFNVk+h75qFYxEVEjv1+GythSXu6NIHQThmeEjkwYgmvteYMyOdR2GKHsVgr+tb+1SiEI0q6V
3dB49NUHh8plVN49z5yAAiuDZKEyJ43z0uW2ixllQDYUwoVvKVx9/OKZjqeCuWjHRwrUezyqwGsG
DSmIjCuTup7uHuCaefEntuvNvbkRYSSUcw2r801NJ+uk/p/tvBtjIckX5iC2Rw==
`pragma protect end_protected
