.GT_REFCLK0(gt_refclk0),
.altclk(altclk_m),
.axisclk(axisclk_m),
.apb3clk(apb3clk_m),
.apb3presetn(apb3presetn_m),
.apb3paddr(apb3paddr_m),
.apb3penable(apb3penable_m),
.apb3psel(apb3psel_m),
.apb3pwdata(apb3pwdata_m),
.apb3pwrite(apb3pwrite_m),
.apb3prdata(apb3prdata_m),
.apb3pready(apb3pready_m),
.apb3pslverr(apb3pslverr_m),
.bgbypassb(bgbypassb_m),
.bgmonitorenb(bgmonitorenb_m),
.bgpdb(bgpdb_m),
.bgrcalovrdenb(bgrcalovrdenb_m),
.bgrcalovrd(bgrcalovrd_m),
.rcalenb(rcalenb_m),
.trigackout0(trigackout0_m),
.trigin0(trigin0_m),
.ubenable(ubenable_m),
.ubiolmbrst(ubiolmbrst_m),
.ubmbrst(ubmbrst_m),
.ctrlrsvdin1(ctrlrsvdin1_m),
.ubintr(ubintr_m),
.gpi(gpi_m),
.ubrxuart(ubrxuart_m),
.ctrlrsvdin0(ctrlrsvdin0_m),
.correcterr(correcterr_m),
.debugtracetvalid(debugtracetvalid_m),
.refclk0_gtrefclkpd(refclk0_gtrefclkpd_m),
.refclk0_clktestsig(refclk0_clktestsig_m),
.refclk1_gtrefclkpd(refclk1_gtrefclkpd_m),
.refclk1_clktestsig(refclk1_clktestsig_m),
.trigackin0(trigackin0_m),
.trigout0(trigout0_m),
.ubinterrupt(ubinterrupt_m),
.ubtxuart(ubtxuart_m),
.uncorrecterr(uncorrecterr_m),
.gpo(gpo_m),
.debugtraceclk(debugtraceclk_m),
.debugtracetdata(debugtracetdata_m),
.ctrlrsvdout(ctrlrsvdout_m),
.ch0_clkrsvd0(ch0_clkrsvd0_m),
.ch0_clkrsvd1(ch0_clkrsvd1_m),
.ch0_loopback(ch0_loopback_m),
.ch0_gtrsvd(ch0_gtrsvd_m),
.ch0_tstin(ch0_tstin_m),
.ch0_pcsrsvdout(ch0_pcsrsvdout_m),
.ch0_pinrsvdas(ch0_pinrsvdas_m),
.ch0_dmonfiforeset(ch0_dmonfiforeset_m),
.ch0_dmonitorclk(ch0_dmonitorclk_m),
.ch0_dmonitorout(ch0_dmonitorout_m),
.ch0_resetexception(ch0_resetexception_m),
.ch0_phyready(ch0_phyready_m),
.ch0_hsdppcsreset(ch0_hsdppcsreset_m),
.ch0_phyesmadaptsave(ch0_phyesmadaptsave_m),
.ch0_iloresetmask(ch0_iloresetmask_m),
.ch0_pcsrsvdin(ch0_pcsrsvdin_m),
.ch1_clkrsvd0(ch1_clkrsvd0_m),
.ch1_clkrsvd1(ch1_clkrsvd1_m),
.ch1_loopback(ch1_loopback_m),
.ch1_gtrsvd(ch1_gtrsvd_m),
.ch1_tstin(ch1_tstin_m),
.ch1_pcsrsvdout(ch1_pcsrsvdout_m),
.ch1_pinrsvdas(ch1_pinrsvdas_m),
.ch1_dmonfiforeset(ch1_dmonfiforeset_m),
.ch1_dmonitorclk(ch1_dmonitorclk_m),
.ch1_dmonitorout(ch1_dmonitorout_m),
.ch1_resetexception(ch1_resetexception_m),
.ch1_phyready(ch1_phyready_m),
.ch1_hsdppcsreset(ch1_hsdppcsreset_m),
.ch1_phyesmadaptsave(ch1_phyesmadaptsave_m),
.ch1_iloresetmask(ch1_iloresetmask_m),
.ch1_pcsrsvdin(ch1_pcsrsvdin_m),
.ch2_clkrsvd0(ch2_clkrsvd0_m),
.ch2_clkrsvd1(ch2_clkrsvd1_m),
.ch2_loopback(ch2_loopback_m),
.ch2_gtrsvd(ch2_gtrsvd_m),
.ch2_tstin(ch2_tstin_m),
.ch2_pcsrsvdout(ch2_pcsrsvdout_m),
.ch2_pinrsvdas(ch2_pinrsvdas_m),
.ch2_dmonfiforeset(ch2_dmonfiforeset_m),
.ch2_dmonitorclk(ch2_dmonitorclk_m),
.ch2_dmonitorout(ch2_dmonitorout_m),
.ch2_resetexception(ch2_resetexception_m),
.ch2_phyready(ch2_phyready_m),
.ch2_hsdppcsreset(ch2_hsdppcsreset_m),
.ch2_phyesmadaptsave(ch2_phyesmadaptsave_m),
.ch2_iloresetmask(ch2_iloresetmask_m),
.ch2_pcsrsvdin(ch2_pcsrsvdin_m),
.ch3_clkrsvd0(ch3_clkrsvd0_m),
.ch3_clkrsvd1(ch3_clkrsvd1_m),
.ch3_loopback(ch3_loopback_m),
.ch3_gtrsvd(ch3_gtrsvd_m),
.ch3_tstin(ch3_tstin_m),
.ch3_pcsrsvdout(ch3_pcsrsvdout_m),
.ch3_pinrsvdas(ch3_pinrsvdas_m),
.ch3_dmonfiforeset(ch3_dmonfiforeset_m),
.ch3_dmonitorclk(ch3_dmonitorclk_m),
.ch3_dmonitorout(ch3_dmonitorout_m),
.ch3_resetexception(ch3_resetexception_m),
.ch3_phyready(ch3_phyready_m),
.ch3_hsdppcsreset(ch3_hsdppcsreset_m),
.ch3_phyesmadaptsave(ch3_phyesmadaptsave_m),
.ch3_iloresetmask(ch3_iloresetmask_m),
.ch3_pcsrsvdin(ch3_pcsrsvdin_m),
.ch0_iloreset(ch0_iloreset_m),
.ch0_pcierstb(ch0_pcierstb_m),
.ch0_bufgtcemask(ch0_bufgtcemask_m),
.ch0_bufgtce(ch0_bufgtce_m),
.ch0_bufgtdiv(ch0_bufgtdiv_m),
.ch0_bufgtrstmask(ch0_bufgtrstmask_m),
.ch0_bufgtrst(ch0_bufgtrst_m),
.ch1_bufgtcemask(ch1_bufgtcemask_m),
.ch1_bufgtce(ch1_bufgtce_m),
.ch1_bufgtdiv(ch1_bufgtdiv_m),
.ch1_bufgtrstmask(ch1_bufgtrstmask_m),
.ch1_bufgtrst(ch1_bufgtrst_m),
.ch2_bufgtcemask(ch2_bufgtcemask_m),
.ch2_bufgtce(ch2_bufgtce_m),
.ch2_bufgtdiv(ch2_bufgtdiv_m),
.ch2_bufgtrstmask(ch2_bufgtrstmask_m),
.ch2_bufgtrst(ch2_bufgtrst_m),
.ch3_bufgtcemask(ch3_bufgtcemask_m),
.ch3_bufgtce(ch3_bufgtce_m),
.ch3_bufgtdiv(ch3_bufgtdiv_m),
.ch3_bufgtrstmask(ch3_bufgtrstmask_m),
.ch3_bufgtrst(ch3_bufgtrst_m),
.ch0_iloresetdone(ch0_iloresetdone_m),
.ch0_phystatus(ch0_phystatus_m),
.ch0_rxcdrhold(ch0_rxcdrhold_m),
.ch0_rxcdrovrden(ch0_rxcdrovrden_m),
.ch0_rxcdrreset(ch0_rxcdrreset_m),
.ch0_rxchbondi(ch0_rxchbondi_m),
.ch0_rxdapicodeovrden(ch0_rxdapicodeovrden_m),
.ch0_rxdapicodereset(ch0_rxdapicodereset_m),
.ch0_rxdlyalignreq(ch0_rxdlyalignreq_m),
.ch0_rxeqtraining(ch0_rxeqtraining_m),
.ch0_rxgearboxslip(ch0_rxgearboxslip_m),
.ch0_rxlatclk(ch0_rxlatclk_m),
.ch0_rxlpmen(ch0_rxlpmen_m),
.ch0_rxmldchaindone(ch0_rxmldchaindone_m),
.ch0_rxmldchainreq(ch0_rxmldchainreq_m),
.ch0_rxmlfinealignreq(ch0_rxmlfinealignreq_m),
.ch0_rxoobreset(ch0_rxoobreset_m),
.ch0_rxpcsresetmask(ch0_rxpcsresetmask_m),
.ch0_rxpd(ch0_rxpd_m),
.ch0_rxphalignreq(ch0_rxphalignreq_m),
.ch0_rxphalignresetmask(ch0_rxphalignresetmask_m),
.ch0_rxphdlypd(ch0_rxphdlypd_m),
.ch0_rxphdlyreset(ch0_rxphdlyreset_m),
.ch0_rxphsetinitreq(ch0_rxphsetinitreq_m),
.ch0_rxphshift180(ch0_rxphshift180_m),
.ch0_rxpmaresetmask(ch0_rxpmaresetmask_m),
.ch0_rxpolarity(ch0_rxpolarity_m),
.ch0_rxprbscntreset(ch0_rxprbscntreset_m),
.ch0_rxprbssel(ch0_rxprbssel_m),
.ch0_rxprogdivreset(ch0_rxprogdivreset_m),
.ch0_rxrate(ch0_rxrate_m),
.ch0_rxresetmode(ch0_rxresetmode_m),
.ch0_rxslide(ch0_rxslide_m),
.ch0_rxsyncallin(ch0_rxsyncallin_m),
.ch0_rxtermination(ch0_rxtermination_m),
.ch0_rxuserrdy(ch0_rxuserrdy_m),
.ch0_rxusrclk(ch0_rxusrclk_m),
.ch0_rx10gstat(ch0_rx10gstat_m),
.ch0_rxbufstatus(ch0_rxbufstatus_m),
.ch0_rxbyteisaligned(ch0_rxbyteisaligned_m),
.ch0_rxbyterealign(ch0_rxbyterealign_m),
.ch0_rxcdrlock(ch0_rxcdrlock_m),
.ch0_rxcdrphdone(ch0_rxcdrphdone_m),
.ch0_rxchanbondseq(ch0_rxchanbondseq_m),
.ch0_rxchanisaligned(ch0_rxchanisaligned_m),
.ch0_rxchanrealign(ch0_rxchanrealign_m),
.ch0_rxchbondo(ch0_rxchbondo_m),
.ch0_rxclkcorcnt(ch0_rxclkcorcnt_m),
.ch0_rxcominitdet(ch0_rxcominitdet_m),
.ch0_rxcommadet(ch0_rxcommadet_m),
.ch0_rxcomsasdet(ch0_rxcomsasdet_m),
.ch0_rxcomwakedet(ch0_rxcomwakedet_m),
.ch0_rxctrl0(ch0_rxctrl0_m),
.ch0_rxctrl1(ch0_rxctrl1_m),
.ch0_rxctrl2(ch0_rxctrl2_m),
.ch0_rxctrl3(ch0_rxctrl3_m),
.ch0_rxdataextendrsvd(ch0_rxdataextendrsvd_m),
.ch0_rxdatavalid(ch0_rxdatavalid_m),
.ch0_rxdata(ch0_rxdata_m),
.ch0_rxdccdone(ch0_rxdccdone_m),
.ch0_rxdlyalignerr(ch0_rxdlyalignerr_m),
.ch0_rxdlyalignprog(ch0_rxdlyalignprog_m),
.ch0_rxelecidle(ch0_rxelecidle_m),
.ch0_rxfinealigndone(ch0_rxfinealigndone_m),
.ch0_rxheadervalid(ch0_rxheadervalid_m),
.ch0_rxheader(ch0_rxheader_m),
.ch0_rxosintdone(ch0_rxosintdone_m),
.ch0_rxosintstarted(ch0_rxosintstarted_m),
.ch0_rxosintstrobedone(ch0_rxosintstrobedone_m),
.ch0_rxosintstrobestarted(ch0_rxosintstrobestarted_m),
.ch0_rxoutclk(ch0_rxoutclk_m),
.ch0_txoutclk(ch0_txoutclk_m),
.ch0_rxphaligndone(ch0_rxphaligndone_m),
.ch0_rxphalignerr(ch0_rxphalignerr_m),
.ch0_rxphdlyresetdone(ch0_rxphdlyresetdone_m),
.ch0_rxphsetinitdone(ch0_rxphsetinitdone_m),
.ch0_rxphshift180done(ch0_rxphshift180done_m),
.ch0_rxpmaresetdone(ch0_rxpmaresetdone_m),
.ch0_rxprbserr(ch0_rxprbserr_m),
.ch0_rxprbslocked(ch0_rxprbslocked_m),
.ch0_rxresetdone(ch0_rxresetdone_m),
.ch0_rxsliderdy(ch0_rxsliderdy_m),
.ch0_rxstartofseq(ch0_rxstartofseq_m),
.ch0_rxstatus(ch0_rxstatus_m),
.ch0_rxsyncdone(ch0_rxsyncdone_m),
.ch0_rxvalid(ch0_rxvalid_m),
.ch0_txcomsas(ch0_txcomsas_m),
.ch0_txcomwake(ch0_txcomwake_m),
.ch0_txctrl0(ch0_txctrl0_m),
.ch0_txctrl1(ch0_txctrl1_m),
.ch0_txctrl2(ch0_txctrl2_m),
.ch0_txdapicodeovrden(ch0_txdapicodeovrden_m),
.ch0_txdapicodereset(ch0_txdapicodereset_m),
.ch0_txdataextendrsvd(ch0_txdataextendrsvd_m),
.ch0_txdata(ch0_txdata_m),
.ch0_txdeemph(ch0_txdeemph_m),
.ch0_txdetectrx(ch0_txdetectrx_m),
.ch0_txdiffctrl(ch0_txdiffctrl_m),
.ch0_txdlyalignreq(ch0_txdlyalignreq_m),
.ch0_txelecidle(ch0_txelecidle_m),
.ch0_txheader(ch0_txheader_m),
.ch0_txinhibit(ch0_txinhibit_m),
.ch0_txlatclk(ch0_txlatclk_m),
.ch0_txmaincursor(ch0_txmaincursor_m),
.ch0_txmargin(ch0_txmargin_m),
.ch0_txmldchaindone(ch0_txmldchaindone_m),
.ch0_txmldchainreq(ch0_txmldchainreq_m),
.ch0_txoneszeros(ch0_txoneszeros_m),
.ch0_txpausedelayalign(ch0_txpausedelayalign_m),
.ch0_txpcsresetmask(ch0_txpcsresetmask_m),
.ch0_txpd(ch0_txpd_m),
.ch0_txphalignreq(ch0_txphalignreq_m),
.ch0_txphalignresetmask(ch0_txphalignresetmask_m),
.ch0_txphdlypd(ch0_txphdlypd_m),
.ch0_txphdlyreset(ch0_txphdlyreset_m),
.ch0_txphdlytstclk(ch0_txphdlytstclk_m),
.ch0_txphsetinitreq(ch0_txphsetinitreq_m),
.ch0_txphshift180(ch0_txphshift180_m),
.ch0_txpicodeovrden(ch0_txpicodeovrden_m),
.ch0_txpicodereset(ch0_txpicodereset_m),
.ch0_txpippmen(ch0_txpippmen_m),
.ch0_txpippmstepsize(ch0_txpippmstepsize_m),
.ch0_txpisopd(ch0_txpisopd_m),
.ch0_txpmaresetmask(ch0_txpmaresetmask_m),
.ch0_txpolarity(ch0_txpolarity_m),
.ch0_txpostcursor(ch0_txpostcursor_m),
.ch0_txprbsforceerr(ch0_txprbsforceerr_m),
.ch0_txprbssel(ch0_txprbssel_m),
.ch0_txprecursor(ch0_txprecursor_m),
.ch0_txprogdivreset(ch0_txprogdivreset_m),
.ch0_txrate(ch0_txrate_m),
.ch0_txresetmode(ch0_txresetmode_m),
.ch0_txsequence(ch0_txsequence_m),
.ch0_txswing(ch0_txswing_m),
.ch0_txuserrdy(ch0_txuserrdy_m),
.ch0_txusrclk(ch0_txusrclk_m),
.ch0_tx10gstat(ch0_tx10gstat_m),
.ch0_txbufstatus(ch0_txbufstatus_m),
.ch0_txcomfinish(ch0_txcomfinish_m),
.ch0_txdccdone(ch0_txdccdone_m),
.ch0_txdlyalignerr(ch0_txdlyalignerr_m),
.ch0_txdlyalignprog(ch0_txdlyalignprog_m),
.ch0_txphaligndone(ch0_txphaligndone_m),
.ch0_txphalignerr(ch0_txphalignerr_m),
.ch0_txphalignoutrsvd(ch0_txphalignoutrsvd_m),
.ch0_txphdlyresetdone(ch0_txphdlyresetdone_m),
.ch0_txphshift180done(ch0_txphshift180done_m),
.ch0_txpmaresetdone(ch0_txpmaresetdone_m),
.ch0_txresetdone(ch0_txresetdone_m),
.ch0_txsyncdone(ch0_txsyncdone_m),
.ch0_gttxreset(ch0_gttxreset_m),
.ch0_txcominit(ch0_txcominit_m),
.ch0_txphsetinitdone(ch0_txphsetinitdone_m),
.ch0_txprogdivresetdone(ch0_txprogdivresetdone_m),
.ch0_txsyncallin(ch0_txsyncallin_m),
.ch1_iloreset(ch1_iloreset_m),
.ch1_pcierstb(ch1_pcierstb_m),
.ch1_iloresetdone(ch1_iloresetdone_m),
.ch1_phystatus(ch1_phystatus_m),
.ch1_rxcdrhold(ch1_rxcdrhold_m),
.ch1_rxcdrovrden(ch1_rxcdrovrden_m),
.ch1_rxcdrreset(ch1_rxcdrreset_m),
.ch1_rxchbondi(ch1_rxchbondi_m),
.ch1_rxdapicodeovrden(ch1_rxdapicodeovrden_m),
.ch1_rxdapicodereset(ch1_rxdapicodereset_m),
.ch1_rxdlyalignreq(ch1_rxdlyalignreq_m),
.ch1_rxeqtraining(ch1_rxeqtraining_m),
.ch1_rxgearboxslip(ch1_rxgearboxslip_m),
.ch1_rxlatclk(ch1_rxlatclk_m),
.ch1_rxlpmen(ch1_rxlpmen_m),
.ch1_rxmldchaindone(ch1_rxmldchaindone_m),
.ch1_rxmldchainreq(ch1_rxmldchainreq_m),
.ch1_rxmlfinealignreq(ch1_rxmlfinealignreq_m),
.ch1_rxoobreset(ch1_rxoobreset_m),
.ch1_rxpcsresetmask(ch1_rxpcsresetmask_m),
.ch1_rxpd(ch1_rxpd_m),
.ch1_rxphalignreq(ch1_rxphalignreq_m),
.ch1_rxphalignresetmask(ch1_rxphalignresetmask_m),
.ch1_rxphdlypd(ch1_rxphdlypd_m),
.ch1_rxphdlyreset(ch1_rxphdlyreset_m),
.ch1_rxphsetinitreq(ch1_rxphsetinitreq_m),
.ch1_rxphshift180(ch1_rxphshift180_m),
.ch1_rxpmaresetmask(ch1_rxpmaresetmask_m),
.ch1_rxpolarity(ch1_rxpolarity_m),
.ch1_rxprbscntreset(ch1_rxprbscntreset_m),
.ch1_rxprbssel(ch1_rxprbssel_m),
.ch1_rxprogdivreset(ch1_rxprogdivreset_m),
.ch1_rxrate(ch1_rxrate_m),
.ch1_rxresetmode(ch1_rxresetmode_m),
.ch1_rxslide(ch1_rxslide_m),
.ch1_rxsyncallin(ch1_rxsyncallin_m),
.ch1_rxtermination(ch1_rxtermination_m),
.ch1_rxuserrdy(ch1_rxuserrdy_m),
.ch1_rxusrclk(ch1_rxusrclk_m),
.ch1_rx10gstat(ch1_rx10gstat_m),
.ch1_rxbufstatus(ch1_rxbufstatus_m),
.ch1_rxbyteisaligned(ch1_rxbyteisaligned_m),
.ch1_rxbyterealign(ch1_rxbyterealign_m),
.ch1_rxcdrlock(ch1_rxcdrlock_m),
.ch1_rxcdrphdone(ch1_rxcdrphdone_m),
.ch1_rxchanbondseq(ch1_rxchanbondseq_m),
.ch1_rxchanisaligned(ch1_rxchanisaligned_m),
.ch1_rxchanrealign(ch1_rxchanrealign_m),
.ch1_rxchbondo(ch1_rxchbondo_m),
.ch1_rxclkcorcnt(ch1_rxclkcorcnt_m),
.ch1_rxcominitdet(ch1_rxcominitdet_m),
.ch1_rxcommadet(ch1_rxcommadet_m),
.ch1_rxcomsasdet(ch1_rxcomsasdet_m),
.ch1_rxcomwakedet(ch1_rxcomwakedet_m),
.ch1_rxctrl0(ch1_rxctrl0_m),
.ch1_rxctrl1(ch1_rxctrl1_m),
.ch1_rxctrl2(ch1_rxctrl2_m),
.ch1_rxctrl3(ch1_rxctrl3_m),
.ch1_rxdataextendrsvd(ch1_rxdataextendrsvd_m),
.ch1_rxdatavalid(ch1_rxdatavalid_m),
.ch1_rxdata(ch1_rxdata_m),
.ch1_rxdccdone(ch1_rxdccdone_m),
.ch1_rxdlyalignerr(ch1_rxdlyalignerr_m),
.ch1_rxdlyalignprog(ch1_rxdlyalignprog_m),
.ch1_rxelecidle(ch1_rxelecidle_m),
.ch1_rxfinealigndone(ch1_rxfinealigndone_m),
.ch1_rxheadervalid(ch1_rxheadervalid_m),
.ch1_rxheader(ch1_rxheader_m),
.ch1_rxosintdone(ch1_rxosintdone_m),
.ch1_rxosintstarted(ch1_rxosintstarted_m),
.ch1_rxosintstrobedone(ch1_rxosintstrobedone_m),
.ch1_rxosintstrobestarted(ch1_rxosintstrobestarted_m),
.ch1_rxphaligndone(ch1_rxphaligndone_m),
.ch1_rxphalignerr(ch1_rxphalignerr_m),
.ch1_rxphdlyresetdone(ch1_rxphdlyresetdone_m),
.ch1_rxphsetinitdone(ch1_rxphsetinitdone_m),
.ch1_rxphshift180done(ch1_rxphshift180done_m),
.ch1_rxpmaresetdone(ch1_rxpmaresetdone_m),
.ch1_rxprbserr(ch1_rxprbserr_m),
.ch1_rxprbslocked(ch1_rxprbslocked_m),
.ch1_rxresetdone(ch1_rxresetdone_m),
.ch1_rxsliderdy(ch1_rxsliderdy_m),
.ch1_rxstartofseq(ch1_rxstartofseq_m),
.ch1_rxstatus(ch1_rxstatus_m),
.ch1_rxsyncdone(ch1_rxsyncdone_m),
.ch1_rxvalid(ch1_rxvalid_m),
.ch1_txcomsas(ch1_txcomsas_m),
.ch1_txcomwake(ch1_txcomwake_m),
.ch1_txctrl0(ch1_txctrl0_m),
.ch1_txctrl1(ch1_txctrl1_m),
.ch1_txctrl2(ch1_txctrl2_m),
.ch1_txdapicodeovrden(ch1_txdapicodeovrden_m),
.ch1_txdapicodereset(ch1_txdapicodereset_m),
.ch1_txdataextendrsvd(ch1_txdataextendrsvd_m),
.ch1_txdata(ch1_txdata_m),
.ch1_txdeemph(ch1_txdeemph_m),
.ch1_txdetectrx(ch1_txdetectrx_m),
.ch1_txdiffctrl(ch1_txdiffctrl_m),
.ch1_txdlyalignreq(ch1_txdlyalignreq_m),
.ch1_txelecidle(ch1_txelecidle_m),
.ch1_txheader(ch1_txheader_m),
.ch1_txinhibit(ch1_txinhibit_m),
.ch1_txlatclk(ch1_txlatclk_m),
.ch1_txmaincursor(ch1_txmaincursor_m),
.ch1_txmargin(ch1_txmargin_m),
.ch1_txmldchaindone(ch1_txmldchaindone_m),
.ch1_txmldchainreq(ch1_txmldchainreq_m),
.ch1_txoneszeros(ch1_txoneszeros_m),
.ch1_txpausedelayalign(ch1_txpausedelayalign_m),
.ch1_txpcsresetmask(ch1_txpcsresetmask_m),
.ch1_txpd(ch1_txpd_m),
.ch1_txphalignreq(ch1_txphalignreq_m),
.ch1_txphalignresetmask(ch1_txphalignresetmask_m),
.ch1_txphdlypd(ch1_txphdlypd_m),
.ch1_txphdlyreset(ch1_txphdlyreset_m),
.ch1_txphdlytstclk(ch1_txphdlytstclk_m),
.ch1_txphsetinitreq(ch1_txphsetinitreq_m),
.ch1_txphshift180(ch1_txphshift180_m),
.ch1_txpicodeovrden(ch1_txpicodeovrden_m),
.ch1_txpicodereset(ch1_txpicodereset_m),
.ch1_txpippmen(ch1_txpippmen_m),
.ch1_txpippmstepsize(ch1_txpippmstepsize_m),
.ch1_txpisopd(ch1_txpisopd_m),
.ch1_txpmaresetmask(ch1_txpmaresetmask_m),
.ch1_txpolarity(ch1_txpolarity_m),
.ch1_txpostcursor(ch1_txpostcursor_m),
.ch1_txprbsforceerr(ch1_txprbsforceerr_m),
.ch1_txprbssel(ch1_txprbssel_m),
.ch1_txprecursor(ch1_txprecursor_m),
.ch1_txprogdivreset(ch1_txprogdivreset_m),
.ch1_txrate(ch1_txrate_m),
.ch1_txresetmode(ch1_txresetmode_m),
.ch1_txsequence(ch1_txsequence_m),
.ch1_txswing(ch1_txswing_m),
.ch1_txsyncallin(ch1_txsyncallin_m),
.ch1_txuserrdy(ch1_txuserrdy_m),
.ch1_txusrclk(ch1_txusrclk_m),
.ch1_tx10gstat(ch1_tx10gstat_m),
.ch1_txbufstatus(ch1_txbufstatus_m),
.ch1_txcomfinish(ch1_txcomfinish_m),
.ch1_txdccdone(ch1_txdccdone_m),
.ch1_txdlyalignerr(ch1_txdlyalignerr_m),
.ch1_txdlyalignprog(ch1_txdlyalignprog_m),
.ch1_txphaligndone(ch1_txphaligndone_m),
.ch1_txphalignerr(ch1_txphalignerr_m),
.ch1_txphalignoutrsvd(ch1_txphalignoutrsvd_m),
.ch1_txphdlyresetdone(ch1_txphdlyresetdone_m),
.ch1_txphshift180done(ch1_txphshift180done_m),
.ch1_txpmaresetdone(ch1_txpmaresetdone_m),
.ch1_txresetdone(ch1_txresetdone_m),
.ch1_txsyncdone(ch1_txsyncdone_m),
.ch1_gttxreset(ch1_gttxreset_m),
.ch1_txcominit(ch1_txcominit_m),
.ch1_txphsetinitdone(ch1_txphsetinitdone_m),
.ch1_txprogdivresetdone(ch1_txprogdivresetdone_m),
.ch2_iloreset(ch2_iloreset_m),
.ch2_pcierstb(ch2_pcierstb_m),
.ch2_iloresetdone(ch2_iloresetdone_m),
.ch2_phystatus(ch2_phystatus_m),
.ch2_rxcdrhold(ch2_rxcdrhold_m),
.ch2_rxcdrovrden(ch2_rxcdrovrden_m),
.ch2_rxcdrreset(ch2_rxcdrreset_m),
.ch2_rxchbondi(ch2_rxchbondi_m),
.ch2_rxdapicodeovrden(ch2_rxdapicodeovrden_m),
.ch2_rxdapicodereset(ch2_rxdapicodereset_m),
.ch2_rxdlyalignreq(ch2_rxdlyalignreq_m),
.ch2_rxeqtraining(ch2_rxeqtraining_m),
.ch2_rxgearboxslip(ch2_rxgearboxslip_m),
.ch2_rxlatclk(ch2_rxlatclk_m),
.ch2_rxlpmen(ch2_rxlpmen_m),
.ch2_rxmldchaindone(ch2_rxmldchaindone_m),
.ch2_rxmldchainreq(ch2_rxmldchainreq_m),
.ch2_rxmlfinealignreq(ch2_rxmlfinealignreq_m),
.ch2_rxoobreset(ch2_rxoobreset_m),
.ch2_rxpcsresetmask(ch2_rxpcsresetmask_m),
.ch2_rxpd(ch2_rxpd_m),
.ch2_rxphalignreq(ch2_rxphalignreq_m),
.ch2_rxphalignresetmask(ch2_rxphalignresetmask_m),
.ch2_rxphdlypd(ch2_rxphdlypd_m),
.ch2_rxphdlyreset(ch2_rxphdlyreset_m),
.ch2_rxphsetinitreq(ch2_rxphsetinitreq_m),
.ch2_rxphshift180(ch2_rxphshift180_m),
.ch2_rxpmaresetmask(ch2_rxpmaresetmask_m),
.ch2_rxpolarity(ch2_rxpolarity_m),
.ch2_rxprbscntreset(ch2_rxprbscntreset_m),
.ch2_rxprbssel(ch2_rxprbssel_m),
.ch2_rxprogdivreset(ch2_rxprogdivreset_m),
.ch2_rxrate(ch2_rxrate_m),
.ch2_rxresetmode(ch2_rxresetmode_m),
.ch2_rxslide(ch2_rxslide_m),
.ch2_rxsyncallin(ch2_rxsyncallin_m),
.ch2_rxtermination(ch2_rxtermination_m),
.ch2_rxuserrdy(ch2_rxuserrdy_m),
.ch2_rxusrclk(ch2_rxusrclk_m),
.ch2_rx10gstat(ch2_rx10gstat_m),
.ch2_rxbufstatus(ch2_rxbufstatus_m),
.ch2_rxbyteisaligned(ch2_rxbyteisaligned_m),
.ch2_rxbyterealign(ch2_rxbyterealign_m),
.ch2_rxcdrlock(ch2_rxcdrlock_m),
.ch2_rxcdrphdone(ch2_rxcdrphdone_m),
.ch2_rxchanbondseq(ch2_rxchanbondseq_m),
.ch2_rxchanisaligned(ch2_rxchanisaligned_m),
.ch2_rxchanrealign(ch2_rxchanrealign_m),
.ch2_rxchbondo(ch2_rxchbondo_m),
.ch2_rxclkcorcnt(ch2_rxclkcorcnt_m),
.ch2_rxcominitdet(ch2_rxcominitdet_m),
.ch2_rxcommadet(ch2_rxcommadet_m),
.ch2_rxcomsasdet(ch2_rxcomsasdet_m),
.ch2_rxcomwakedet(ch2_rxcomwakedet_m),
.ch2_rxctrl0(ch2_rxctrl0_m),
.ch2_rxctrl1(ch2_rxctrl1_m),
.ch2_rxctrl2(ch2_rxctrl2_m),
.ch2_rxctrl3(ch2_rxctrl3_m),
.ch2_rxdataextendrsvd(ch2_rxdataextendrsvd_m),
.ch2_rxdatavalid(ch2_rxdatavalid_m),
.ch2_rxdata(ch2_rxdata_m),
.ch2_rxdccdone(ch2_rxdccdone_m),
.ch2_rxdlyalignerr(ch2_rxdlyalignerr_m),
.ch2_rxdlyalignprog(ch2_rxdlyalignprog_m),
.ch2_rxelecidle(ch2_rxelecidle_m),
.ch2_rxfinealigndone(ch2_rxfinealigndone_m),
.ch2_rxheadervalid(ch2_rxheadervalid_m),
.ch2_rxheader(ch2_rxheader_m),
.ch2_rxosintdone(ch2_rxosintdone_m),
.ch2_rxosintstarted(ch2_rxosintstarted_m),
.ch2_rxosintstrobedone(ch2_rxosintstrobedone_m),
.ch2_rxosintstrobestarted(ch2_rxosintstrobestarted_m),
.ch2_rxphaligndone(ch2_rxphaligndone_m),
.ch2_rxphalignerr(ch2_rxphalignerr_m),
.ch2_rxphdlyresetdone(ch2_rxphdlyresetdone_m),
.ch2_rxphsetinitdone(ch2_rxphsetinitdone_m),
.ch2_rxphshift180done(ch2_rxphshift180done_m),
.ch2_rxpmaresetdone(ch2_rxpmaresetdone_m),
.ch2_rxprbserr(ch2_rxprbserr_m),
.ch2_rxprbslocked(ch2_rxprbslocked_m),
.ch2_rxresetdone(ch2_rxresetdone_m),
.ch2_rxsliderdy(ch2_rxsliderdy_m),
.ch2_rxstartofseq(ch2_rxstartofseq_m),
.ch2_rxstatus(ch2_rxstatus_m),
.ch2_rxsyncdone(ch2_rxsyncdone_m),
.ch2_rxvalid(ch2_rxvalid_m),
.ch2_txcomsas(ch2_txcomsas_m),
.ch2_txcomwake(ch2_txcomwake_m),
.ch2_txctrl0(ch2_txctrl0_m),
.ch2_txctrl1(ch2_txctrl1_m),
.ch2_txctrl2(ch2_txctrl2_m),
.ch2_txdapicodeovrden(ch2_txdapicodeovrden_m),
.ch2_txdapicodereset(ch2_txdapicodereset_m),
.ch2_txdataextendrsvd(ch2_txdataextendrsvd_m),
.ch2_txdata(ch2_txdata_m),
.ch2_txdeemph(ch2_txdeemph_m),
.ch2_txdetectrx(ch2_txdetectrx_m),
.ch2_txdiffctrl(ch2_txdiffctrl_m),
.ch2_txdlyalignreq(ch2_txdlyalignreq_m),
.ch2_txelecidle(ch2_txelecidle_m),
.ch2_txheader(ch2_txheader_m),
.ch2_txinhibit(ch2_txinhibit_m),
.ch2_txlatclk(ch2_txlatclk_m),
.ch2_txmaincursor(ch2_txmaincursor_m),
.ch2_txmargin(ch2_txmargin_m),
.ch2_txmldchaindone(ch2_txmldchaindone_m),
.ch2_txmldchainreq(ch2_txmldchainreq_m),
.ch2_txoneszeros(ch2_txoneszeros_m),
.ch2_txpausedelayalign(ch2_txpausedelayalign_m),
.ch2_txpcsresetmask(ch2_txpcsresetmask_m),
.ch2_txpd(ch2_txpd_m),
.ch2_txphalignreq(ch2_txphalignreq_m),
.ch2_txphalignresetmask(ch2_txphalignresetmask_m),
.ch2_txphdlypd(ch2_txphdlypd_m),
.ch2_txphdlyreset(ch2_txphdlyreset_m),
.ch2_txphdlytstclk(ch2_txphdlytstclk_m),
.ch2_txphsetinitreq(ch2_txphsetinitreq_m),
.ch2_txphshift180(ch2_txphshift180_m),
.ch2_txpicodeovrden(ch2_txpicodeovrden_m),
.ch2_txpicodereset(ch2_txpicodereset_m),
.ch2_txpippmen(ch2_txpippmen_m),
.ch2_txpippmstepsize(ch2_txpippmstepsize_m),
.ch2_txpisopd(ch2_txpisopd_m),
.ch2_txpmaresetmask(ch2_txpmaresetmask_m),
.ch2_txpolarity(ch2_txpolarity_m),
.ch2_txpostcursor(ch2_txpostcursor_m),
.ch2_txprbsforceerr(ch2_txprbsforceerr_m),
.ch2_txprbssel(ch2_txprbssel_m),
.ch2_txprecursor(ch2_txprecursor_m),
.ch2_txprogdivreset(ch2_txprogdivreset_m),
.ch2_txrate(ch2_txrate_m),
.ch2_txresetmode(ch2_txresetmode_m),
.ch2_txsequence(ch2_txsequence_m),
.ch2_txswing(ch2_txswing_m),
.ch2_txsyncallin(ch2_txsyncallin_m),
.ch2_txuserrdy(ch2_txuserrdy_m),
.ch2_txusrclk(ch2_txusrclk_m),
.ch2_tx10gstat(ch2_tx10gstat_m),
.ch2_txbufstatus(ch2_txbufstatus_m),
.ch2_txcomfinish(ch2_txcomfinish_m),
.ch2_txdccdone(ch2_txdccdone_m),
.ch2_txdlyalignerr(ch2_txdlyalignerr_m),
.ch2_txdlyalignprog(ch2_txdlyalignprog_m),
.ch2_txphaligndone(ch2_txphaligndone_m),
.ch2_txphalignerr(ch2_txphalignerr_m),
.ch2_txphalignoutrsvd(ch2_txphalignoutrsvd_m),
.ch2_txphdlyresetdone(ch2_txphdlyresetdone_m),
.ch2_txphshift180done(ch2_txphshift180done_m),
.ch2_txpmaresetdone(ch2_txpmaresetdone_m),
.ch2_txresetdone(ch2_txresetdone_m),
.ch2_txsyncdone(ch2_txsyncdone_m),
.ch2_gttxreset(ch2_gttxreset_m),
.ch2_txcominit(ch2_txcominit_m),
.ch2_txphsetinitdone(ch2_txphsetinitdone_m),
.ch2_txprogdivresetdone(ch2_txprogdivresetdone_m),
.ch3_iloreset(ch3_iloreset_m),
.ch3_pcierstb(ch3_pcierstb_m),
.ch3_iloresetdone(ch3_iloresetdone_m),
.ch3_phystatus(ch3_phystatus_m),
.ch3_rxcdrhold(ch3_rxcdrhold_m),
.ch3_rxcdrovrden(ch3_rxcdrovrden_m),
.ch3_rxcdrreset(ch3_rxcdrreset_m),
.ch3_rxchbondi(ch3_rxchbondi_m),
.ch3_rxdapicodeovrden(ch3_rxdapicodeovrden_m),
.ch3_rxdapicodereset(ch3_rxdapicodereset_m),
.ch3_rxdlyalignreq(ch3_rxdlyalignreq_m),
.ch3_rxeqtraining(ch3_rxeqtraining_m),
.ch3_rxgearboxslip(ch3_rxgearboxslip_m),
.ch3_rxlatclk(ch3_rxlatclk_m),
.ch3_rxlpmen(ch3_rxlpmen_m),
.ch3_rxmldchaindone(ch3_rxmldchaindone_m),
.ch3_rxmldchainreq(ch3_rxmldchainreq_m),
.ch3_rxmlfinealignreq(ch3_rxmlfinealignreq_m),
.ch3_rxoobreset(ch3_rxoobreset_m),
.ch3_rxpcsresetmask(ch3_rxpcsresetmask_m),
.ch3_rxpd(ch3_rxpd_m),
.ch3_rxphalignreq(ch3_rxphalignreq_m),
.ch3_rxphalignresetmask(ch3_rxphalignresetmask_m),
.ch3_rxphdlypd(ch3_rxphdlypd_m),
.ch3_rxphdlyreset(ch3_rxphdlyreset_m),
.ch3_rxphsetinitreq(ch3_rxphsetinitreq_m),
.ch3_rxphshift180(ch3_rxphshift180_m),
.ch3_rxpmaresetmask(ch3_rxpmaresetmask_m),
.ch3_rxpolarity(ch3_rxpolarity_m),
.ch3_rxprbscntreset(ch3_rxprbscntreset_m),
.ch3_rxprbssel(ch3_rxprbssel_m),
.ch3_rxprogdivreset(ch3_rxprogdivreset_m),
.ch3_rxrate(ch3_rxrate_m),
.ch3_rxresetmode(ch3_rxresetmode_m),
.ch3_rxslide(ch3_rxslide_m),
.ch3_rxsyncallin(ch3_rxsyncallin_m),
.ch3_rxtermination(ch3_rxtermination_m),
.ch3_rxuserrdy(ch3_rxuserrdy_m),
.ch3_rxusrclk(ch3_rxusrclk_m),
.ch3_rx10gstat(ch3_rx10gstat_m),
.ch3_rxbufstatus(ch3_rxbufstatus_m),
.ch3_rxbyteisaligned(ch3_rxbyteisaligned_m),
.ch3_rxbyterealign(ch3_rxbyterealign_m),
.ch3_rxcdrlock(ch3_rxcdrlock_m),
.ch3_rxcdrphdone(ch3_rxcdrphdone_m),
.ch3_rxchanbondseq(ch3_rxchanbondseq_m),
.ch3_rxchanisaligned(ch3_rxchanisaligned_m),
.ch3_rxchanrealign(ch3_rxchanrealign_m),
.ch3_rxchbondo(ch3_rxchbondo_m),
.ch3_rxclkcorcnt(ch3_rxclkcorcnt_m),
.ch3_rxcominitdet(ch3_rxcominitdet_m),
.ch3_rxcommadet(ch3_rxcommadet_m),
.ch3_rxcomsasdet(ch3_rxcomsasdet_m),
.ch3_rxcomwakedet(ch3_rxcomwakedet_m),
.ch3_rxctrl0(ch3_rxctrl0_m),
.ch3_rxctrl1(ch3_rxctrl1_m),
.ch3_rxctrl2(ch3_rxctrl2_m),
.ch3_rxctrl3(ch3_rxctrl3_m),
.ch3_rxdataextendrsvd(ch3_rxdataextendrsvd_m),
.ch3_rxdatavalid(ch3_rxdatavalid_m),
.ch3_rxdata(ch3_rxdata_m),
.ch3_rxdccdone(ch3_rxdccdone_m),
.ch3_rxdlyalignerr(ch3_rxdlyalignerr_m),
.ch3_rxdlyalignprog(ch3_rxdlyalignprog_m),
.ch3_rxelecidle(ch3_rxelecidle_m),
.ch3_rxfinealigndone(ch3_rxfinealigndone_m),
.ch3_rxheadervalid(ch3_rxheadervalid_m),
.ch3_rxheader(ch3_rxheader_m),
.ch3_rxosintdone(ch3_rxosintdone_m),
.ch3_rxosintstarted(ch3_rxosintstarted_m),
.ch3_rxosintstrobedone(ch3_rxosintstrobedone_m),
.ch3_rxosintstrobestarted(ch3_rxosintstrobestarted_m),
.ch3_rxphaligndone(ch3_rxphaligndone_m),
.ch3_rxphalignerr(ch3_rxphalignerr_m),
.ch3_rxphdlyresetdone(ch3_rxphdlyresetdone_m),
.ch3_rxphsetinitdone(ch3_rxphsetinitdone_m),
.ch3_rxphshift180done(ch3_rxphshift180done_m),
.ch3_rxpmaresetdone(ch3_rxpmaresetdone_m),
.ch3_rxprbserr(ch3_rxprbserr_m),
.ch3_rxprbslocked(ch3_rxprbslocked_m),
.ch3_rxresetdone(ch3_rxresetdone_m),
.ch3_rxsliderdy(ch3_rxsliderdy_m),
.ch3_rxstartofseq(ch3_rxstartofseq_m),
.ch3_rxstatus(ch3_rxstatus_m),
.ch3_rxsyncdone(ch3_rxsyncdone_m),
.ch3_rxvalid(ch3_rxvalid_m),
.ch3_txcomsas(ch3_txcomsas_m),
.ch3_txcomwake(ch3_txcomwake_m),
.ch3_txctrl0(ch3_txctrl0_m),
.ch3_txctrl1(ch3_txctrl1_m),
.ch3_txctrl2(ch3_txctrl2_m),
.ch3_txdapicodeovrden(ch3_txdapicodeovrden_m),
.ch3_txdapicodereset(ch3_txdapicodereset_m),
.ch3_txdataextendrsvd(ch3_txdataextendrsvd_m),
.ch3_txdata(ch3_txdata_m),
.ch3_txdeemph(ch3_txdeemph_m),
.ch3_txdetectrx(ch3_txdetectrx_m),
.ch3_txdiffctrl(ch3_txdiffctrl_m),
.ch3_txdlyalignreq(ch3_txdlyalignreq_m),
.ch3_txelecidle(ch3_txelecidle_m),
.ch3_txheader(ch3_txheader_m),
.ch3_txinhibit(ch3_txinhibit_m),
.ch3_txlatclk(ch3_txlatclk_m),
.ch3_txmaincursor(ch3_txmaincursor_m),
.ch3_txmargin(ch3_txmargin_m),
.ch3_txmldchaindone(ch3_txmldchaindone_m),
.ch3_txmldchainreq(ch3_txmldchainreq_m),
.ch3_txoneszeros(ch3_txoneszeros_m),
.ch3_txpausedelayalign(ch3_txpausedelayalign_m),
.ch3_txpcsresetmask(ch3_txpcsresetmask_m),
.ch3_txpd(ch3_txpd_m),
.ch3_txphalignreq(ch3_txphalignreq_m),
.ch3_txphalignresetmask(ch3_txphalignresetmask_m),
.ch3_txphdlypd(ch3_txphdlypd_m),
.ch3_txphdlyreset(ch3_txphdlyreset_m),
.ch3_txphdlytstclk(ch3_txphdlytstclk_m),
.ch3_txphsetinitreq(ch3_txphsetinitreq_m),
.ch3_txphshift180(ch3_txphshift180_m),
.ch3_txpicodeovrden(ch3_txpicodeovrden_m),
.ch3_txpicodereset(ch3_txpicodereset_m),
.ch3_txpippmen(ch3_txpippmen_m),
.ch3_txpippmstepsize(ch3_txpippmstepsize_m),
.ch3_txpisopd(ch3_txpisopd_m),
.ch3_txpmaresetmask(ch3_txpmaresetmask_m),
.ch3_txpolarity(ch3_txpolarity_m),
.ch3_txpostcursor(ch3_txpostcursor_m),
.ch3_txprbsforceerr(ch3_txprbsforceerr_m),
.ch3_txprbssel(ch3_txprbssel_m),
.ch3_txprecursor(ch3_txprecursor_m),
.ch3_txprogdivreset(ch3_txprogdivreset_m),
.ch3_txrate(ch3_txrate_m),
.ch3_txresetmode(ch3_txresetmode_m),
.ch3_txsequence(ch3_txsequence_m),
.ch3_txswing(ch3_txswing_m),
.ch3_txsyncallin(ch3_txsyncallin_m),
.ch3_txuserrdy(ch3_txuserrdy_m),
.ch3_txusrclk(ch3_txusrclk_m),
.ch3_tx10gstat(ch3_tx10gstat_m),
.ch3_txbufstatus(ch3_txbufstatus_m),
.ch3_txcomfinish(ch3_txcomfinish_m),
.ch3_txdccdone(ch3_txdccdone_m),
.ch3_txdlyalignerr(ch3_txdlyalignerr_m),
.ch3_txdlyalignprog(ch3_txdlyalignprog_m),
.ch3_txphaligndone(ch3_txphaligndone_m),
.ch3_txphalignerr(ch3_txphalignerr_m),
.ch3_txphalignoutrsvd(ch3_txphalignoutrsvd_m),
.ch3_txphdlyresetdone(ch3_txphdlyresetdone_m),
.ch3_txphshift180done(ch3_txphshift180done_m),
.ch3_txpmaresetdone(ch3_txpmaresetdone_m),
.ch3_txresetdone(ch3_txresetdone_m),
.ch3_txsyncdone(ch3_txsyncdone_m),
.ch3_gttxreset(ch3_gttxreset_m),
.ch3_txcominit(ch3_txcominit_m),
.ch3_txphsetinitdone(ch3_txphsetinitdone_m),
.ch3_txprogdivresetdone(ch3_txprogdivresetdone_m),
.hsclk0_lcpllclkrsvd0(hsclk0_lcpllclkrsvd0_m),
.hsclk0_lcpllclkrsvd1(hsclk0_lcpllclkrsvd1_m),
.hsclk0_lcpllfbdiv(hsclk0_lcpllfbdiv_m),
.hsclk0_lcpllpd(hsclk0_lcpllpd_m),
.hsclk0_lcpllrefclksel(hsclk0_lcpllrefclksel_m),
.hsclk0_lcpllresetbypassmode(hsclk0_lcpllresetbypassmode_m),
.hsclk0_lcpllresetmask(hsclk0_lcpllresetmask_m),
.hsclk0_lcpllreset(hsclk0_lcpllreset_m),
.hsclk0_lcpllrsvd0(hsclk0_lcpllrsvd0_m),
.hsclk0_lcpllrsvd1(hsclk0_lcpllrsvd1_m),
.hsclk0_lcpllsdmdata(hsclk0_lcpllsdmdata_m),
.hsclk0_lcpllsdmtoggle(hsclk0_lcpllsdmtoggle_m),
.hsclk0_rpllclkrsvd0(hsclk0_rpllclkrsvd0_m),
.hsclk0_rpllclkrsvd1(hsclk0_rpllclkrsvd1_m),
.hsclk0_rpllfbdiv(hsclk0_rpllfbdiv_m),
.hsclk0_rpllpd(hsclk0_rpllpd_m),
.hsclk0_rpllrefclksel(hsclk0_rpllrefclksel_m),
.hsclk0_rpllresetbypassmode(hsclk0_rpllresetbypassmode_m),
.hsclk0_rpllresetmask(hsclk0_rpllresetmask_m),
.hsclk0_rpllreset(hsclk0_rpllreset_m),
.hsclk0_rpllrsvd0(hsclk0_rpllrsvd0_m),
.hsclk0_rpllrsvd1(hsclk0_rpllrsvd1_m),
.hsclk0_rpllsdmdata(hsclk0_rpllsdmdata_m),
.hsclk0_rpllsdmtoggle(hsclk0_rpllsdmtoggle_m),
.hsclk0_lcpllfbclklost(hsclk0_lcpllfbclklost_m),
.hsclk0_lcpllrefclklost(hsclk0_lcpllrefclklost_m),
.hsclk0_rpllfbclklost(hsclk0_rpllfbclklost_m),
.hsclk0_rpllrefclklost(hsclk0_rpllrefclklost_m),
.hsclk0_lcpllrefclkmonitor(hsclk0_lcpllrefclkmonitor_m),
.hsclk0_rpllrefclkmonitor(hsclk0_rpllrefclkmonitor_m),
.hsclk0_lcpllrsvdout(hsclk0_lcpllrsvdout_m),
.hsclk0_rpllrsvdout(hsclk0_rpllrsvdout_m),
.hsclk1_lcpllclkrsvd0(hsclk1_lcpllclkrsvd0_m),
.hsclk1_lcpllclkrsvd1(hsclk1_lcpllclkrsvd1_m),
.hsclk1_lcpllfbdiv(hsclk1_lcpllfbdiv_m),
.hsclk1_lcpllpd(hsclk1_lcpllpd_m),
.hsclk1_lcpllrefclksel(hsclk1_lcpllrefclksel_m),
.hsclk1_lcpllresetbypassmode(hsclk1_lcpllresetbypassmode_m),
.hsclk1_lcpllresetmask(hsclk1_lcpllresetmask_m),
.hsclk1_lcpllreset(hsclk1_lcpllreset_m),
.hsclk1_lcpllrsvd0(hsclk1_lcpllrsvd0_m),
.hsclk1_lcpllrsvd1(hsclk1_lcpllrsvd1_m),
.hsclk1_lcpllsdmdata(hsclk1_lcpllsdmdata_m),
.hsclk1_lcpllsdmtoggle(hsclk1_lcpllsdmtoggle_m),
.hsclk1_rpllclkrsvd0(hsclk1_rpllclkrsvd0_m),
.hsclk1_rpllclkrsvd1(hsclk1_rpllclkrsvd1_m),
.hsclk1_rpllfbdiv(hsclk1_rpllfbdiv_m),
.hsclk1_rpllpd(hsclk1_rpllpd_m),
.hsclk1_rpllrefclksel(hsclk1_rpllrefclksel_m),
.hsclk1_rpllresetbypassmode(hsclk1_rpllresetbypassmode_m),
.hsclk1_rpllresetmask(hsclk1_rpllresetmask_m),
.hsclk1_rpllreset(hsclk1_rpllreset_m),
.hsclk1_rpllrsvd0(hsclk1_rpllrsvd0_m),
.hsclk1_rpllrsvd1(hsclk1_rpllrsvd1_m),
.hsclk1_rpllsdmdata(hsclk1_rpllsdmdata_m),
.hsclk1_rpllsdmtoggle(hsclk1_rpllsdmtoggle_m),
.hsclk1_lcpllfbclklost(hsclk1_lcpllfbclklost_m),
.hsclk1_lcpllrefclklost(hsclk1_lcpllrefclklost_m),
.hsclk1_rpllfbclklost(hsclk1_rpllfbclklost_m),
.hsclk1_rpllrefclklost(hsclk1_rpllrefclklost_m),
.hsclk1_lcpllrefclkmonitor(hsclk1_lcpllrefclkmonitor_m),
.hsclk1_rpllrefclkmonitor(hsclk1_rpllrefclkmonitor_m),
.hsclk1_lcpllrsvdout(hsclk1_lcpllrsvdout_m),
.hsclk1_rpllrsvdout(hsclk1_rpllrsvdout_m),
.s0_axis_tready(m0_axis_tready_m),
.s0_axis_tdata(m0_axis_tdata_m),
.s0_axis_tlast(m0_axis_tlast_m),
.s0_axis_tvalid(m0_axis_tvalid_m),
.s1_axis_tready(m1_axis_tready_m),
.s1_axis_tdata(m1_axis_tdata_m),
.s1_axis_tlast(m1_axis_tlast_m),
.s1_axis_tvalid(m1_axis_tvalid_m),
.s2_axis_tready(m2_axis_tready_m),
.s2_axis_tdata(m2_axis_tdata_m),
.s2_axis_tlast(m2_axis_tlast_m),
.s2_axis_tvalid(m2_axis_tvalid_m),
.pcielinkreachtarget(pcielinkreachtarget_m),
.pcieltssm(pcieltssm_m),
.rxmarginclk(rxmarginclk_m),
.rxmarginreqcmd(rxmarginreqcmd_m),
.rxmarginreqlanenum(rxmarginreqlanenum_m),
.rxmarginreqpayld(rxmarginreqpayld_m),
.rxmarginreqreq(rxmarginreqreq_m),
.rxmarginresack(rxmarginresack_m),
.rxmarginresreq(rxmarginresreq_m),
.rxmarginreqack(rxmarginreqack_m),
.rxmarginrescmd(rxmarginrescmd_m),
.rxmarginreslanenum(rxmarginreslanenum_m),
.rxmarginrespayld(rxmarginrespayld_m),
.m0_axis_tready(s0_axis_tready_m),
.m0_axis_tdata(s0_axis_tdata_m),
.m0_axis_tlast(s0_axis_tlast_m),
.m0_axis_tvalid(s0_axis_tvalid_m),
.m1_axis_tready(s1_axis_tready_m),
.m1_axis_tdata(s1_axis_tdata_m),
.m1_axis_tlast(s1_axis_tlast_m),
.m1_axis_tvalid(s1_axis_tvalid_m),
.m2_axis_tready(s2_axis_tready_m),
.m2_axis_tdata(s2_axis_tdata_m),
.m2_axis_tlast(s2_axis_tlast_m),
.m2_axis_tvalid(s2_axis_tvalid_m),
.gtpowergood(gtpowergood_m),
.ch0_rxprogdivresetdone(ch0_rxprogdivresetdone_m),
.ch0_gtrxreset(ch0_gtrxreset_m),
.ch0_cdrbmcdrreq(ch0_cdrbmcdrreq_m),
.ch0_cdrfreqos(ch0_cdrfreqos_m),
.ch0_cdrincpctrl(ch0_cdrincpctrl_m),
.ch0_cdrstepdir(ch0_cdrstepdir_m),
.ch0_cdrstepsq(ch0_cdrstepsq_m),
.ch0_cdrstepsx(ch0_cdrstepsx_m),
.ch0_cfokovrdfinish(ch0_cfokovrdfinish_m),
.ch0_cfokovrdpulse(ch0_cfokovrdpulse_m),
.ch0_cfokovrdstart(ch0_cfokovrdstart_m),
.ch0_eyescanreset(ch0_eyescanreset_m),
.ch0_eyescantrigger(ch0_eyescantrigger_m),
.ch0_eyescandataerror(ch0_eyescandataerror_m),
.ch0_cfokovrdrdy0(ch0_cfokovrdrdy0_m),
.ch0_cfokovrdrdy1(ch0_cfokovrdrdy1_m),
.ch1_rxprogdivresetdone(ch1_rxprogdivresetdone_m),
.ch1_gtrxreset(ch1_gtrxreset_m),
.ch1_cdrbmcdrreq(ch1_cdrbmcdrreq_m),
.ch1_cdrfreqos(ch1_cdrfreqos_m),
.ch1_cdrincpctrl(ch1_cdrincpctrl_m),
.ch1_cdrstepdir(ch1_cdrstepdir_m),
.ch1_cdrstepsq(ch1_cdrstepsq_m),
.ch1_cdrstepsx(ch1_cdrstepsx_m),
.ch1_cfokovrdfinish(ch1_cfokovrdfinish_m),
.ch1_cfokovrdpulse(ch1_cfokovrdpulse_m),
.ch1_cfokovrdstart(ch1_cfokovrdstart_m),
.ch1_eyescanreset(ch1_eyescanreset_m),
.ch1_eyescantrigger(ch1_eyescantrigger_m),
.ch1_eyescandataerror(ch1_eyescandataerror_m),
.ch1_cfokovrdrdy0(ch1_cfokovrdrdy0_m),
.ch1_cfokovrdrdy1(ch1_cfokovrdrdy1_m),
.ch2_rxprogdivresetdone(ch2_rxprogdivresetdone_m),
.ch2_gtrxreset(ch2_gtrxreset_m),
.ch2_cdrbmcdrreq(ch2_cdrbmcdrreq_m),
.ch2_cdrfreqos(ch2_cdrfreqos_m),
.ch2_cdrincpctrl(ch2_cdrincpctrl_m),
.ch2_cdrstepdir(ch2_cdrstepdir_m),
.ch2_cdrstepsq(ch2_cdrstepsq_m),
.ch2_cdrstepsx(ch2_cdrstepsx_m),
.ch2_cfokovrdfinish(ch2_cfokovrdfinish_m),
.ch2_cfokovrdpulse(ch2_cfokovrdpulse_m),
.ch2_cfokovrdstart(ch2_cfokovrdstart_m),
.ch2_eyescanreset(ch2_eyescanreset_m),
.ch2_eyescantrigger(ch2_eyescantrigger_m),
.ch2_eyescandataerror(ch2_eyescandataerror_m),
.ch2_cfokovrdrdy0(ch2_cfokovrdrdy0_m),
.ch2_cfokovrdrdy1(ch2_cfokovrdrdy1_m),
.ch3_rxprogdivresetdone(ch3_rxprogdivresetdone_m),
.ch3_gtrxreset(ch3_gtrxreset_m),
.ch3_cdrbmcdrreq(ch3_cdrbmcdrreq_m),
.ch3_cdrfreqos(ch3_cdrfreqos_m),
.ch3_cdrincpctrl(ch3_cdrincpctrl_m),
.ch3_cdrstepdir(ch3_cdrstepdir_m),
.ch3_cdrstepsq(ch3_cdrstepsq_m),
.ch3_cdrstepsx(ch3_cdrstepsx_m),
.ch3_cfokovrdfinish(ch3_cfokovrdfinish_m),
.ch3_cfokovrdpulse(ch3_cfokovrdpulse_m),
.ch3_cfokovrdstart(ch3_cfokovrdstart_m),
.ch3_eyescanreset(ch3_eyescanreset_m),
.ch3_eyescantrigger(ch3_eyescantrigger_m),
.ch3_eyescandataerror(ch3_eyescandataerror_m),
.ch3_cfokovrdrdy0(ch3_cfokovrdrdy0_m),
.ch3_cfokovrdrdy1(ch3_cfokovrdrdy1_m),
.hsclk0_lcplllock(hsclk0_lcplllock_m),
.hsclk0_rplllock(hsclk0_rplllock_m),
.hsclk1_lcplllock(hsclk1_lcplllock_m),
.hsclk1_rplllock(hsclk1_rplllock_m),
.debugtraceready(  debugtracetready_m),
.ch0_txmstreset     (ch0_msttxreset_m),
.ch0_txmstresetdone (ch0_msttxresetdone_m),
.ch1_txmstreset     (ch1_msttxreset_m),
.ch1_txmstresetdone (ch1_msttxresetdone_m),
.ch2_txmstreset     (ch2_msttxreset_m),
.ch2_txmstresetdone (ch2_msttxresetdone_m),
.ch3_txmstreset     (ch3_msttxreset_m),
.ch3_txmstresetdone (ch3_msttxresetdone_m),
.ch0_rxmstreset      ( ch0_mstrxreset_m ),
.ch0_rxmstresetdone  ( ch0_mstrxresetdone_m),
.ch1_rxmstreset      ( ch1_mstrxreset_m),
.ch1_rxmstresetdone  ( ch1_mstrxresetdone_m),
.ch2_rxmstreset      ( ch2_mstrxreset_m),
.ch2_rxmstresetdone  ( ch2_mstrxresetdone_m),
.ch3_rxmstreset      ( ch3_mstrxreset_m),
.ch3_rxmstresetdone  ( ch3_mstrxresetdone_m),
.rxn(gt_quad_base_serial_rxn),
.rxp(gt_quad_base_serial_rxp),
.txn(gt_quad_base_serial_txn),
.txp(gt_quad_base_serial_txp),
.refclk0_gtrefclkpdint(refclk0_gtrefclkpdint),
.pipenorthout(pipenorthoutq0_to_pipenorthinq1),
.resetdone_northout(resetdone_northout_q0_to_resetdone_northin_q1), 
.rxpinorthout(rxpinorthout_q0_to_rxpinorthin_q1), 
.txpinorthout(txpinorthout_q0_to_txpinorthin_q1), 
.pipesouthin( pipesouthin_q0_to_pipesouthout_q1),  
.resetdone_southin(resetdone_southin_q0_to_resetdone_southout_q1), 
.rxpisouthin(rxpisouthin_to_rxpsouthout_q1), 
.txpisouthin(txpisouthin_to_txpsouthout_q1) 
