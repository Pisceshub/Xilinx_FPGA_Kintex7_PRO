`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15952)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9JQaMgpupSUIgDmsbAQQ3DIx8z3pNa2pGEVlZCP/TzE0x8ycv+pSJiks
r071EYbc4hdeCHe/16wjR7f73cbFPXhgyb7dmJRm0CiWNkMgcNk5zJnG4pSF7gjokzyDd10x3x4y
9fI9QstUbOZ7kSeTGMMfh958r2Le6r6MAm2PlSW+P3nFy92THIqojBEq57b32NwfrMx+1UUnv8O9
5XoOvHRVchFETuXHMTEghaEU8NxQ8vv378pKVTPyuyf1QIcIf1n1mHPdWcJcgvVg3mY1fvOuiRfr
XM98AkMuG2hFjqSYQcdtBFI/ZzLMg4/G9AMcfOLZYWJMunpf82XXFM/7vORUX9l63Rz/y2jvBSGR
0wi/kjiONB4ix+Hb21fssY/ciypTKcDLRAx0dOWpkyAYLaOAb2t4dbHWbO0Jm2hko/gYR23/frX9
tgJoxlD8ifujO+LcAdczZTE5C9/XDas5syjdHuLrkEpSuYNfsJtHA2KjcY8PBuTdqSVp/DSVn5j/
OtJ9nj06k4svzyV6yJ8IGVbX77c/R+TTrGXVNsJr5yObZLXemLBAmZJBH/qui1/NwrYhFsoDd/0L
VV94EExN02DQG5IoSH9a2BZKZxoZXlQEkc5cBPMHeFMk+SRvxQuGLmH1yxXgZpA1jlx4CyY34i8c
EuXkWJnrsTU2Iiy6Wr6PO23w70vUUxOtV22w4Jm1zSi9X/PHoNzJio4roIi5pQuOR4REDr8Z0U4+
EyAt520TNUiMdh81irX99wonpr+FNmP6bFViBMY9k4NXq+HIB3p9Kju/NNwMsU/qLvENh5NTgsWR
MNGwWhGPLHhPzTm10GBK28hXISLyq6bD5B3MfJJhcItIiSHavfcauaGSOCGySZPpy2Mi/bITJ38d
PEzYeNwnrJv05FmELHOYWfC9ZtgEy/YFFBX1L6taYp+ik+klEFUskybEO/11vzLN+06ooV0eNbX3
UNNnemRQ8oCFHnZVU4ErzVnbxnc3YpyWhQmWHJSlsv4BZzbif8YVc0erlrUDbgtu/8CZKWfYuFdi
AUQGEaocIc2a/3HWcWRtmutx8LxOAFubM1Gbf+gokSBREmfibfSEDWb4Pk0eLO4QGtHLoHNooa8N
mv0qrIxk8ZohMh4Sr58+yKA0Ju6a4PwGsaYv9SwwkLWzzQQYnAG9Kk4f3yrBwzLADu018OEVuddG
sCEIqsuyU8YRIDb6M7P1rGV+J8Kd2gzq4qUxqZw0FqzaxjTwXSpJ0HjBSEDhTQOSPHLJ+9shK/Xx
ivI5K0LEbFW1GPKf5eelns1yfi3UiuEElmAYLuY5worSwL3/b+kAKkid4l3uBZF9KvnnzOjQ2goh
IAozgK8sWKda9xwKu9Z9clJH+J/UwoMBHNFcJ4buDHBM70ENSSV+a5lKHcWzNkpGCQlu2SPEKU0w
Vd/v35MRJ1w0bK8F6budeL4rd4rTkECYqz09D+2jNU6/wurV2F19GK8yeX7oP321591OxspKmJJm
5yK/VI3nwYdR02d9mhO5NfDGqoH3NIZDDP4tVhBtPfE6aMP31HiegRDwGOqhCs2Gu7DqAP5JHwjg
5JHN61SspGdduXLVQ1vWh8MngHUWZUFQlCc6yBtbY5q2+2bNgcnklaCAhGtcRszHnaOkbLUL+bRZ
i3pJ0uxsPoZ/mZTIx1q2qrjh47USwRtcmuk5W3WYCpr7WLzqJWSGheoFQFORVHIT5aDwEJ0eiZRF
FakzbSL6/i2/7b7txPCvcJgVm4+/nQftbGINO5JdcdIVnybnstMLD+7rWrndUN7oXrpIfygnruk1
pet2bVYzCn99f5tYzM8NXv/n1JiweiOaPo1s6734gIpGL/zFIXSFsMlIyaXKK5FrJbEf80MKPXp/
8Jfh7rWnSUCnFDYs3CBiBz1C/mf4JV6m7kL5PXagBpJRejIszyfpaBtAmKh1gVPZO8fnch1Xw+dD
mVSWPC///w+GZDADqlKif2KpMN/+unv88cL/vYvOJPfnFAKWwlmL5jGTMqIXJIyWpCuLYurA2Yju
hxNzf1qSPCYnkiqvyw3FYv/IHEmD4OO+Q153jCt7YeR3lahuRITUxM3OGEo8F5qKe5Do65GZPgvh
zEMwyOBf22buSU34qfgHCc+Jl5U8aC/Raka3Yj8+/RXeJeJEyFBUaFfhANPWM1OgI3H467L9bQEy
DdUHbMC6/BuiUbFFZx23y8NkOhCEEXvntgdq7cW1yZBibUs/GlrQo2ENcDCVD8RhQ2pSdJO4m7AZ
BLAWwCQQic7Pw4wm58AsAWwyHiF900Cfx2UzM+cd4Jd9/Q4ZwLRNKW8AW/ftfxTDTdl5Jg8j13dz
2bxljTzj4orHnVNHL75JXIT0037motosoP5ZJo/0tUIFjaMC/m2eTTAOZeqsPNGtSvrDdk/VMt6z
iF9P5OzJx0S79X84tAQ/G1udMKsfvqLb0CsjK2I4H3uFlx0/qHeiEXkQs5s2t3rOg2keVHg6rxI5
k/K0A+XoSZRf3LJn6RLUXx2cyhl324UzGVb+S1iDPoshmJiRM/JSUHAWWeQUqaQFWR3WQuylPzfS
9lY/Tqs84Hb/PlQS6SGqcVK3XD5c2wWf1/oyQchAwYCvlt12WjcrTDTryhrLg3S9tYL+o/s6sWvT
yC3pm+ACAwm4rbEWCNuSb2zUIvJ5aNLWTI3ib5DsatTLlSKskgadn1puvLsyZHFDliJlq161Yxb0
+c5UMibO4SNtSC6nq7PhkPdykutAWrwVIhG67AnCoUfY6WPehv3D75FSJTGcH4YHLuyB04eXg9Da
oOcfc1tVs26RGagGAz7SxaCUmdaAayohxIXaT6Bu+zV5L9md2sArkGjHpD4NI4bLMcPubRV03qJV
TK92Xp0mNCpvE+/enXl3vYNoveKivQzXpTVNKiQQT5ju8LgG8I3bS4F3nuQOg2w+Ym5lbm57Llb3
yC9HFBJGEOcBhhHtbuYiQ+5Q+UsCv4luJVU7OT/GmAVqMoycIEJtYmJm07Ng9jCNYpgSWtyCUxY6
muIus8lrWf2TxepHha74OfoE7XvZ0kyd3UkiVhMFCZ5DXLcG93he81WmQchlp1v5U0dAPaldIxC2
9AxQKDP7zXiMm5djlflPe2+rnyqdUtVJviUR7NhDd9y8Wj1e0ZtQyViy8tMsYRYY0k3+QYWpsJzp
xWm8jdT86TGflJSH+whRkXGCbU++ghw1H+cepd5GQ1HVWX9fcqhzZsgdZAvAOgpyEra/dbh3f1ER
oGBVCFT/ot/ZtDRNYganQnB5C7n12DbkYCvXfaNDw8TUoe18EE74ZneYPiQnIjtcXK27LOay+F8R
qkciM+dSEWfJFJ/h5aEfCVqrob5gxqCHDKcCFXTgnk1drs5EACL7WEHV5GQqHbeH401Bd17ZozZa
eToUduvFTAoqbKpoeXtrDN5eyLO3pEv+N7m+Xscvqy8Vjq/knPBGHJmf8JEZ5ex2UMYytKBQ0cgL
k0zud7oBLJ78ZfPKApVkKfTXxldxS9edK7A02YN7+Oz7rOjhI9j0tp4LXg6N8Gxr8ynD+DAc8Anj
mcZJgQnHEbhgeWCicHFtbIY10sU5hQq3Qwm/wpWq7AzisBWZl8SnuvFaaKQ+U0NTQ1gFryo826eY
TjcEcf9LzNbGEvItBNx7QwaaNC/wSTKgRJ50DntB8BXA6n/e2oGl9Uil16cZ53fYh9EXH1M5Peyk
edzFUNMDTPYtDhVJkMjIgvI+bFENcBC3oXvt+lxuQTPyOQrY3t6BXMyCyu+wfipLZ4mP0v5vrOzX
01E9jK0XCEKDYly1PAQOBGzCJ35j7leoKdAjfSxbIc7k60puV0r7xqYEPxte5JRWQkIfPWhou22Z
LSMvP+20KbXzaoXgTzr66wt1a12VHr3Za0ZkljnJLWiFjzf8r95KQPahOf3nIT5U94a7TbRwbGGK
oA6/RDGIawR3GCczTSxkwMBE2Tphz8ED5LZ6Ytuu2ip0mMMuaWTNpycuZVf22+grN86llRWeitIH
7t40CAqdlDiBAn+itgGiK0QMHckRp4X4RIQP/nH3zSt93usxEAMjGYZeywzlHwvU1tfGclpptV5J
bkvj2PK+nHlgFEa7Y0RfhXL9JnMpydsoWGdDVqm9TdXIp9JlCxhZIilb+97AeG3GHBw7yfraHfGu
vlVHrHHwTu3d+Tc2utVZhJEUObmhmSJ8Fh0rmdtciMLvUvUGtKOwAGNE8L+JSzXcNS1/bek9wKZ3
JyV5o7PNMyJxSFzruF3L1gSIJrSTAZ6912ycILnI8HMUe6byiLUz6SOhNc5MGtQAkdyzHPQcYwyP
fGGqDKCq16yb2s+HEdTRzae0xhpoexjTF3UN2hILDcqM8ErvCG/MJiBzU3N+z7aPH6KQNksDCJrr
PAtQzPDs7kGqOj2FDJQuxcLPYyZc3SfZCIpTP4E2wObBShxeJWhXFoSdk5QLnfJjB4o57blCXyyx
TTtBtr+R16GhU4UfLmhvEAtt0/Keb1QWE4SRa3e9QUhQ950+MXOtC5+f1S65xbKRQbKgnQqnR8ZW
eUR/wW9jlu+MFLRXwcr0LTU8n7cbIjs3BugFRuh2OdMnBpJjLVDVIcO1zah5QeQYRQoHwxG2iRqV
GeNW5+6VF5eoZGo8olQ09o+xATZm0ETnCvveS9OUTJHGFnttm+cPnlFYwUy3V60LEnt1DqWXVhw1
X0T185pf3RSH97jh003n5CaHvTmZn4wzGDtrR9oAO8meVCBLjYC6wvdXoWivZLqIh67pDsFWfvOe
bcMVE/8tz2AEbiVYuORAXPHX6S3WGouxzoEjfGyw06LSuX/npOkGLnIXa8QVDHJk4Sdk5kClNoGL
/A5/s4/na3R0dcPDxTYjnBmM4YctJhIDFMKPq9kVSpcdTpc0YEnqdYKDDV2EbdHRi07YQ7wNXAeb
TdUVbL5b3N4NpJRJHa9ZiGHUfn3P6o8pO7Fz3fhE33w+3QtXuP8zL5ad3zdlUUDSBGsDfaoxyJJK
ADf9/GMeI5S3worFwQh93oAtPA1nFheiSrr/RMJ4k2J2qfqh+8m5ELM0eKrqRRp5LPIUY0tMBcVa
iC+/D2INjvKGuzJTkQEuqzRFp1HQ3AUPUYekLrFL5PuYpErMdF1I6zGZVre9Zcf3G4wxvyawasKr
XOU+aD2+rpolbUF6ZxNtT44M1N56VhMHKMdq8+qFlIpLJKmjjgjsiMVt4YeHlpRmmIb7XTKiGm13
+8nen48gbNKxq463pxJ27PhmNT4NfoBecU3j2+oJ4/Sf9Wlfc5qY9ejHH510i5xfhX27CEE/dqhB
eJghhZq1pNhu+5gTDVps5V/r4Sr96/VbnMuZ8xGJHh/QLpWxokrYzkWW1ytDmEp1qoTBB3ogwVje
X9RlKuiSUAnhUkED+N/e2r4HcYf+n3KqxIVKFA9Xl8erxy7BYQKn/jK+O86UJfrbwx0wJ1dIX4kx
L9elTRbKVeaOLbqsZdM0MB0KT195RhEvpQAfCX3J9ZIWBCtgggXPte+3aonmOS8MyKXUK9IesDBB
gmdfVbVz/cm4dJd5v/8mf+j5KaiDY9szQC2BQ2xsA4UR1rsXagvqzn9SJAqyzKfTSDRF4EtAsX0Q
Z3LuVfRvRzdQQ5c11+PGcVJBikl4V5ImQeP4O8z/d2d22roz2iNl9owyOtMPTVibnF8RnNTvw8xM
OT6y7Sf1Ve2/Ky8/op0TCHh2osxZQ86udfhnMX7y6JDg2OCM7QHfpTWq40mjD0H5PvcQhNJqMXDw
1YZHTv+LDCJWPVEC5gb97t0C2anQXOlc4yhKzbGucy/g8KwgZqut9SOTi8UxnZLMRAxJ7iMX5Kq8
TN3/OaYc9E6RpFpFeeo+ya75WqNfUPVZloGoDH3lrrdhCe+X8TJfJvcU07vN9Txjc0rLHxNrXUWw
g08xpK5fxcOz63TTs8vnS8Kznf+flo1fRxooDJhgYaqnEyEYM2/Br7H7gNgOvfMn/DUwVI24JDXS
Kb36LFjzSACXqZdpW1d8jq1Ys81DOg0fdbK+01BpWOoh34JmqvAv+hRW8zOkK8mwg+H4uuVt1l2f
L6LpZ35R8B7lz8Poct8fYgTn5xt+wtQw2SlkRA909Bz4tAd8EED9aZ3C1kLhjE7Eo8mEJ0lqZ4Dz
4xuFzHlcfvjcdC9uSagUcikNHijrdojlXBYv8O4cED/BmXYohRSZhPyuQGCqnKz9LbyhrNpa9LA/
Q63ptXFhj6QaWAhLNzjEMW/EGPvfIIp0CyBJmsmh5hijqG7IbLNNvZ+YtiZqc6VSyQsMa4+uiNmf
NyJ88kB7HU9tGLC18yU4Otw556tOwc860iOyttPfIcoH/EyT4YuRpIDi9AlaK+cxBNA6aohM1oia
QKFKHz3jISIg82g4wEIAXXLUIyTtBF8cRfftcZc2ViN4Bt6WAaWriY34dh1YAiKqSepEHvTZ98pA
UzfCXtnkSBH5kEXMzhjG8/Uu1uqX5JC93/ay2oQqoGDh7dmdyvOAusnhzFJv4+bASr4ixQ24NjWi
XhvL66SxKV3/KQO8wApSReihAjL0dBbv8yz9pJGU9I/BsvjlBmxJ58475Akq8xYtS50mD9PmFLqw
KfRFIS+1EiNwOClU2EYpVKm+Q3ZX8UNWJgBEmlGHatvlfScGv2LnyO5JarhMbTaYLU0RBc2f4cGK
kOWxCNXzt6awBGklUlVXsPqfu+whHwQ7xG6AWTTA96o+OH82H1pAEdUhwi3sTzcmc2mPQmaC3RKi
bNhPOmIvos5Zx/A4FkZ0YaxuD2h4oJb5OpwdcF01KMFvJAC+aQJ773RyMpPYjoR6RoEUg+a8N65f
ZQNPyNy50FDmd5WuoMrbiWj3oi9KhoPEMsfChzvqNNFPlhr4u4uTjDGi27JHfHWNRqZ5zsEpRopk
pWSqIgRXTCAEyCZ7QImzqk6sI1IgT0TL1vy1l/4pfVqsMXOpf+z/2Z4AFtdD267dYWtXB1Ph7L/0
FInj0MtCyZTV8uwxX0nxCdYLIKhODTQfmSybHFmCTHx6cJslX+Byu7hQ/8NYZj+5b1jhLkv2iO/i
L/gdUlz0VEdETb5ByGTXCRz3rxbphbAqnhJgFOcHw2j60xhbGdC+DrG/je7uB5uZ5Egvi0GuE3yP
Jn05YExnwKHAm/SNkXY58j4u3s5Fk9u7sspkp/hHKEacFApSfPp9sjeYMPWAJcxUok7sgAZijQYa
wJsy+W637rqggxMP3frEMxCt95fmfPm+ounRjtuOco/qjLj6rnfs6wL8bWGK0YV7puSUWJEoTA2o
UD9dZhv85530tgVNLvp+WjMkYiy0Fe+e3LE4ETslYA+Qh1YKA/QQZfPYV73LVhT6lBRjJECXlj5j
5TNwN5TDifQV0CjQbnef0m4jrIfTFsvxO+OnoHgB9QyrTBd6Br/lyjxXWv2vGd1Mrj29w0UewkMI
nPsiU4TFrnXptl/rlzd6l4zWTkh+ybaBZwZKo1X6y0b05ZqkUQvfaUZPMLate+4K5wzkfQrirnv7
rntL8SMWzhqShRuo4hd5ls4h9g48yZljmsWV2bl+kuHcJm10veiNGo0YGl5Qj/MDGH80FG7x9PNi
RFyyp0HPaQ8wwOKUGgp6Hc/yNhOkm8eDJiSmGM5e6fQl5qaG2JfUAnf/5DgeU4EE0vUMuX2AQ89n
8jxASuZqljAum5LsKvqrN6TvfwRMBF5f0FZwaYIZcyYO8VsHE0L3ILMm4nqQVTwiWI5G0ddqpAVS
DoXne+tv4vvPIUs/KbW4uwRe8bsrqwqF/Nv/f67ICV0eTUOgSmL2iOOn15rVmORxjD3hmgZfoZYX
fFoTVpQCKoMYDH2EzbfsFDHUjommjozY9pWbJqR/YrZdvB+FqueVDTbhRa1N8YJ7RaY1C0d215u1
urm6pzbDv6hDnRE6gMXyUlwxs/gy3DyNibMthuS0p52r8vLX2WzZow8e4lsOQEyl44ydrHDmUpTn
AHyxY+rBc6qT4LcubDNdPFjBgP/TIbos6IPKFS3LZl9BMDOPMNU9QuD8KMDSS+F1Wnco7RIq6RRO
v4+N/a1VNG/UngpO/ntrfwuV+Br0OzCTdOuAlOqcuMZUSdxrX8HgqZ/KvesL7kvPUpOFbg9AfwpX
Ticbf87j7Y822ejLIo2QsTED1rGsyZmvrHENRlTu2fDOb2/D3y1DSe+rXbPbkWRRF0npyCkyTHck
MWSFf9opBFjGHFIXB8qYKd5YeeXgUt7Xe9RI9lUUxWNw9DhANCD28xgc3DQj97SzjmCVkQCsWdiE
1z3qhBj0aRBxfkf5hIx6nOl5RrkADTJNX+U6xLDvd1i6PSGlhSZ+sIfUwWQ+ojYpGB9Sq6d4Nvu9
TFF5oX6vslBedhWAHmXOXZu/hRtchbSdO9gG6A4cV+X/FbHCX2unZv5FT3RI/RUOmHFFi/z0yj3G
Zyc9IJVDHbYR+SsHQTpMwd6OPoerC9Q94n9t9u4pvzD9PD47pqVFJy5/yGmffQNWAxxUyxoU1gOv
I0eCA4tHsEAi8Rjd4mzScYA7FAuESW3GCY/xcADBDmbFoW7of94iT19wE7dQ4ngDpOv6MLRVbMgo
DE91KKAZb01xQgsY8iN0jpXLFpsA/sV8eR2zQBWYmvHmIAPyuVdmZx1QARwMw0uEfYAKAn8NQYaW
PiIVzmpwOsT0Hs1ecPLEZpb1JOMBy87/SIWYcW9BKr619Za45gMNnBvWhUTzNOMjXwXf3tIn39RX
Rj18/dIeXvwu5JNQuGWuz7OulTYy2s2kgPVRCRZGfT0TKEAD/2sk/TX9LnW6teTTU/xy5iencKb6
jKn1zx74Jwz7d8HLb/wlpjSPqayga0hA/rNI0ikFVogeL9Qal67zs0gv798yidILiwEQ+vp66xpq
1T3moa6RTdnxQZmrmWuav3snXdZXTi/VjbhnCRGzOaoRLt5rLdIR4LurriKII+1AsdkTkUohlwGd
yWICtdUznYlPMxixl7g30AC9Q/jfwdGJvPkMxLofAYwG7tb6WvPBU1w0vJ6T0diDMuGHMsXsoYxk
jxXSHTkAAERsO7NjKw8tlvUwnMzAwBtcsjHIAvqxp7KkKdupvez7yM4KPwAaiSctCVYLZeJrh6qT
m4iLay2AOTg+gBVq6uXTT+o5ijmOs9HHlT58MdF2jha0O3gfm7wq5ejQtTuDRU4hqDvhrCtDAVyf
A98zZbOTR7w5YTUeJaZaa9lHmlpvw9Pgv6eOeGoczljWFjuEAsLF1Q6sy9KYVC/FzEO31r9Jgdw+
9PnWQyesk8KdNJ6quarFulQVU2MPFK2IfiRbw6HyredaFtu6ICaGjFCHOPukFdBO3kOGGWwUYU21
YLT42arSIMaGaHNOkCsaVP9UAmaPCj4BX0q37iHElu6KuQfAnnH46dJi4LCqFyB80txVdmzUCZuk
tTReFuHLeUSC+6wEJIRWIqfk9A5brHPtXJuxVqZiRi4IL+x0YGjgoROeQhrvc3ghqzLvs4PEaloS
3Y2aVHv3dPcrSGpl2u41a6x1907hUntz5xS+uWyLufLwXmslWNDcNJ8daBTOPiRusUWeC1bzKAsU
Ilvnqf58u0kpox2bo8pWxg82kt1WWuW7wWKx7DzXoinHqmA6spVHfm0a2XFtD4zvPyM4NAsMaHUP
pZmDFEMX3eZGxIDKGrL1Cf60ByZMXCqQplrEkutFxWPzbhUfh9TmFdTcTZlHHTMeFGdKCxsn7EqJ
Bqs0Q0Oox6DIQIUC0Nvwi/HQvYqsuWZopV2aq+N+b6TinvptKJjrG0YmYlS7fVZ9T4U4K3IjobsD
KFZVUqBV/9aVavQhClipcCoiDgEkqihnd1K4S3KiRuIIvxER9lkLnwlAKfjUnC+407/s4QoEJFOm
aneIUF5rFKx5/qdzdJjXGgYZIr25qHWhYz6+A3g9QrhZA0r2psHQT69o4Qgz2+MrkCAcnWSzD9XC
v5yZE9+mPQ5gOFJG+wDkF6WWSLyj/qNJBzhCThQQpKk4WCQetJDPNpQ764x1G2uzDLSMfWx3XoOg
WAmGA52njUBvF62qoUi/ipAduNKG54dacDz6skl2qcOyBdRPTW3lHlLYQ2BRYcOuiUp+diDAW1wD
2g+brSdIgEEeoBBk6baRIhAB7K40Srx/4wew8GLC9HAzjeUprsN4C7eGJ1Zl1lv98Vn/rMtGQJFp
PcTvgquLzoWXNp4IZlT0FsiEz1wPQpcjl0tr5MweFVzkpgRwMeeWopH5BwGHH5thwjaC+jtd4U1J
6I5JWuJTElENbADn4ohd2nt7L5w1p+s6h1rl3Denw9KMIPL001uXXZi2L8ATiHZSVsbSN2tVfVKg
CnL7DivZCvPHDfY18kV+WryvBEJnv+I8zdc05h51IjbLcg7uPBj5SZ55n4sKNA2AWBG0E3tspddD
XCO1M1zpV65eBe2RPnEyBITCTyk+eMYnTvfQMtbg2YLL0maDPP8ppa6YZxGAIufOPs6tgrr4UPW+
xsk0etLGfGqxzF5rxfSLgZjlZrqHm6gP+j9L7dXykiYyqB61ZuPXrcRNQrm+ExvN5CZpq4uZhWu6
quPwwwws+ivs1N0YKJspLTeA6W5zvEoK1A6T3ol3qMTUieHiB2NHHmJxQRqGQ7HKlYOGldwVumSA
K3oKolaFhvFLjl0rWVzd+vXtpKxw7BJmP0R/tEq+DCzcau5LSfln4LPEYE7lAiNHlZVH4SfIpDWy
JD3PJfZzs5mykbwLUSmisZSRwlqcIESy6ETqajmeI+1yQScLvoGlv4SDV1LFrSMJTsruuJQOuP5X
PyXZNUQz4H/UNuLza0BPBPCeLjuACQiYldxcppydWS+6mSDrutLpqi6vkVKQdHPS7ShsSqiIMgW9
5LLBzsYJm+mlb4q4k+XwOwgPKoUvmWK/9hcgHoHU9Adia8K2GUWLaLONEbKOq/0MdVp8vkVIoRch
kNzov+FaALoNIGDEIN93GxKtmo5WOj9N3fgoMLponYQqKntioRH553XHpmQG92nNoyIMZzMCVXti
uXFZJP9UGiDfpDSyUqfAEAPxCIF7WOG8oocwDY35Y3zZwVW9SNQt6aRTg7HBj/m+Ma9TXVTiQVLN
7GY/YxlQ5l7yrEbW2Qcb+Pfnnrqud3bGkE56OLB8NJCdlZp6K3ShLP/+QwL1ZB3LuD5JQJX7feYz
VIgm8OHxTfdZr8ZGeVklLUAG+65uva7l6mDeFgvJQ1HCSQ8Jh2GBXtKn9DlNpdArqwGv7xvSNTWt
xIGe08IukJTctWyZYvz9U/vI04dTgfJv8zEHaEWsOd6c6JJkAMwL0dNlGpHkHq6f1gdCCrKF4rJu
5sBIEpzKQCoomwShBZb6fw5VsKSzP5Gf9lZDYBOy1mgtbLEvbrOnyEchGQMx+9HRrs5U6YdLeh6A
o3HQZLasTlKyrfCkW914dWwpXS7QWmOfC8Zl3AhaqqDc5wHPGiFzPJxIwlVOoHHM8VYLi5Z3X+fq
R3UYEl9mVk62idhrvmzZEZ4GVaCqKtaNVbXYRQ6E4A0ts6qi9k+QxqOJLNo0euNkqYy3MZT4iUEu
fFwQhpchDqQXdIlB1HajXkqQ06iLh+UE1abXe4B18ovNjxNBQixSyTYp7vTRBthc1pQXUjg+6658
CMPGUrIMZBWwlDldB78jnuZsyyeCZoEqYZfFoWVPtZIIGOtihrstV1JgE0HZfWO0VId9Si8hOtmE
2Xy9fUvIdQF5aNP9iLDpfPWwURoXqQRpuP+nAdtkNBhWtGLQ34Sbt8pM5eNL0JEM3qnpnlBtjU0R
P6Covk0Ek97NcGz86J782zx0afbuaIaJwEAk9m4CZs+5x+DdTrmbh2pNRfPYtALZuInX5j/9xwEE
UACIBX3yJHWeXo1Pi85KsZvAnqspYVPunypr3UmAbzhDsB5UTDjHfrMpnWH85A7cM1BbMyjMqeTq
Ja2AsIsO5yOwiFsBQROrRLtlZT+HOSolJHxYjGWR1QQFQ53U1xlCG18JDrKYh9W5Qv9hvSJWQxYw
mpUG8bK4DC+Bz3mzw+ltZdPp8qQH6PQeVCGZQbUUemV/TnoKp8cQaS4Qh8KbOV1AND2gt0T8dse6
0Jbc0jw1OzZUlKgOtbstAq3/lMSo56XJ8iz97LuEKjOv3gOoaZ+3Cu8lfRTHZYruAT9k7E0HvVCL
o1KqeLUQWPF1CBgQY34KPYrgmca3aRDl/pQkku8OS5Ib+C/qRDOBO0MconuuXSVlXLYOgM4umNZe
AltsmSDG9znLB2ZmRJpJN0ThGEdu1p+CWZY7NHwADyv4CbyfyWF6ig9NXsNjBfnUj3qVekkRatIb
RZa9ivkzXBNDzm/Z0u+oE2l6yPLniKssTLuaArNOblNI5L0PD3p7os7DAf7JxPIR/NfG83JBS0X+
V499owv8SsxHQZnXrSj3ElkCaEkUP/mbrlr7o9qkjQ5HhXVcoA5dtNWL9T+9bixpQST/Dv2292f7
gB50wo6fOWI16dTeDn606CbjuQbZ+T4VM6DrQj/8cT9IVEVODgVayJB3wEepw7Jwdwf3QylRE8GW
aqp3fZ72lC22I/Oe1SlB0B1j36Zz+7R4O7TSVoHIxOIZz4vhBzgr1kCcVsx3i1/6Kikg577NZzr0
4NLSOez+As77UemPX1aT4zErQ3UrNjWKNrwG3r91nKJji1i0Wzf4IbtuiBJAieL63yEsPOjU6Ie2
KexyGemGGGCrERIK7J7nIYHQ9Bb7jDA0meS1tf6xxfUa3P0hq0SvK0iV7HFUjlYbA88L9K2Ebxgl
TGGdiG3dt0RkcEojp2RE9Hd8s4puhxQYBwKL66SmmHASsm3kpl17AQNvYQ3e/euWj01M8OwP/YAJ
pEyUuXtZHOJf+gjqLlPBpeUwfeBCxZ16H8QzzO8R+KhyVASeXuQdp0OlxvsEjodzzltJiDW/0m8n
0HZnAf9XiPMnuog5OaW8YyGvz+Q9CM0Cvm7JoVZvCc/MnfiiZ7xA16nrY56Wrz5NIikMfnpzisjy
aFtiV3V8Tu4yuYmLk8i8b6geQ6vjUqi+GORUi476uAuz7zS+3Waz0P38ZXPbmA0/9WO78Mlk071V
mcNxjlgexJehBR3R/MJGOI7sXNbO4XAugozFFZKR0OpOQhKFsmFHGBg4de5NwuiA7LpSuOGKUP0n
ShRjCPksZAoI9D6e3NVN/n/PjwB1Ao16CUPjrFdOly0YmmVMUxi8kMxQH7q0HqUqQ0CdUTklD2zs
Ir23LOIGSUSGJpY1VnsDZFGYpDMyz2TthiyAouHkjGE0J2Bp9IW8YidR3Q0ER3vc1Nf1ACJPbKSh
gdabjIQGolrQsCIMfAk6bhA1L8kVtsSZdiFJHBz3/DmIcuUM3vLYJCrDoCG5aO4hFpKbOVDoDBbS
ud+94GdCGN03jE+c42h3T1DGBAuviOPihV2na+TiAeLv2J3ZPC6n4yQi17Qxu4l3kgo0olcYHqkY
Y8FZt95PM77wvd2ilAVzDmnpECZZNtAehteo2qeZsJ/PCl2343IZ58Keql+1Gplef38yoMMwehyE
cU8+55TSzavYxU0wks+5Jri+MYdX7e1GinaT3st6eElMcUz4VsZCf8m2ytD81q5nBjASEuw4bfhb
H0+K01Oa1xvF7WPd6ZFJtj1b8IsZ75f3dVE0gfBR5CQW04JuUlMwbNggv4mvTsbLza/yj4mdzfcR
4mv589KEEfUwOTZ/aLs7jA7EEpfM4lVJEaSB6Q5zsR5V+SAk6WIGUXC9LiIuUcMCFqD+dyrpaQmg
6nbUUA//Wig9nsY2lked5p8Ri95SnIiFfaMdxRdH9//j8JB9bVOh+LI0hPNWDNQEoEVq3pOhvo6u
BD5eI3NkClB9fCgxSknq8CUcxGBHMoPNzQ63x1CAFnwfqSTiG19QLBAfd9uVUAXRnkfNxCQsT4fi
+N3ILDBF+k1qH30Rn96tE6hjSMWcDCgyAYX33LPzWgujkkOeHGwr22gvLyZt4DPKdPhQKrRf9ykc
fZAnXX36x6IOgowWg7cW/yV5tO13fCpW9eGzWh9n9ZvzqfZmvvZRClZEGdusPp3pSZp4x18S+BXr
uYPGmezjFsCtzFI2lF+vsTBTc60Wd7lI3TwgTdYTEmecSztCVoDfSXzCnjnxZGdvOs7z+IghEJ1i
8d0LH+lwgWkG89W1dGgpBlvf2JcWFIGL2EgFqszdKPIdR+YT0uOlVGryVa+s/5GrmWMji0sZ5XrS
4RtemzYJT3W6DYhxr761WTmsFEjw+g7Wx2S0LYzU/sZihaCccOILGKszdTDyLRABCf+brqiKSXHR
cgeUFtuf/B7WQL1S79WCl+RzncTaT2XrDPnLWPP0FCBF7S5w5aMGSQPizGeMCd63sagELICsodQm
MS67wuFgOYpG7L2V5qFdq9j2K76VWh/rxFOuuxClpYgO4CnTILPI94HQK3/xF9V1aAoK5HwgBjj5
KId4MfAu7ywUwb1D3g4/MyQm/0nGXjFrchifYhp5sHGoTmSF6tF85sT3hiQgaEf8fLg5xE6evH8D
wpKcZH861gTqz2f0M5jkocyu3ExD+CBvsJM64Y7uQKyVof80UUNRXp4hwn5eucODc1JGL6pVxA/i
Ye1zBFJdVm/9PtxS6tEFUle4tb+5jbyv7oP9Z/hA2epXqdCKIdI3yGq3uvlyq0oL8R6n48O1UHid
8VwV5P3MP5DJwuwY9prPjh8YFR8DXi8Qarz+y4ZD+WxzSte+ukhOjqXhQonFtN163R/O6obHUc2f
cH6AF4k80T4Oh76CUtXqbbxGcOaGs2avHYqayfXzBm4T44l6zidE5oqkPxQC2S8IF8slluYz4CCQ
hBhXWK/pN7QscFMyWCLHsCfyn5+2oOBn60wFxBW0mkbcR7EjgJe/g5xPwDrJBlPVFRW/muaqf20G
7cqZ1jgOXJshnjU/hYCX8T+3mA5O7s+eZ0Bosw/FvNGRqPX07LiuZPw9f1K6os5o2S47hFhWcMqG
jZCVC/Qg10e4CQjZ4FFOXcJmXSg5CkVMGZLYNOeLkNppU68sGEqWUBcODxV9GDJURIDfawMZvEO3
ojPFhTQAp6rwxo0cKZrnkEEImP/MuyL6v/tPYskVdLzLxXreCXHKrBB9+8OC4hnd23UYTXT1V3nZ
PVHBpzX0zmG8sZVpgrtQRJUOSexdZpauQMnF3FcY7ffdrQNwrpNDgGtPbffLRHeTqBnvmIKihH1J
Lxjib87esTrKF3olyBcdHTAsIrnhxW7g6QwtO/cHDx9kDA2+EGY4SEIKPL7Zn/9zKPgqazRSbiOE
ca/W/noYLkpA2CpSVglSr60q7GpaCow8XrvDQOe1AVkhKlLR35x81ObSj+D8e9gQrR/WKClRzbV1
lUw/TwTIh1uRAGJEcj1Obm2IPVCyz3lTr79B8XrX9pvUjvn+ixl9qf8uwm3kprjn4k1zDCJnbsF1
ZDNfqDgdgZgD+orGEh7hAFnMx1Vd+kslqSsXpDgJyq2k56RNrZt3ZN7UGLLnAXuKmqPl4xe1JWAF
7nLCK2x0ro7IyXXlOdzTnMxg2AIRpnhEIcOVodoc4ablLeeAKKEL2AV+KFoT74A5GOoBnmyjvOQi
16rEzwlzPtco8UksGxQzguL6Is1FYIfghtHPPxTYAy2bh3n7+P/TGlrgp6eU9TJ22vs7zeRxJI7m
a22Oj0yGVwK1Dzi2x2oNIFM4CN8XtQN4UZ7Lo/znAP9qQhG2Sgyl9E0Rqy/26ax1XrEoQLPEaAms
zY3bmWzlF8tiZgJMn3rsKSlJMiACTZYRHoMg6/TMko+/gmrsdL9gUWa6FoJtuk32xIEnhSRB8jW5
WULU951m5R+FcOuHRcI2Zc5WV7a8Ur86hzVybC10OCwSAWl7V2Ldzbtsx84PpG7VFXRzBpaxY1pI
2MAqDFMbEu6JHGsX09WoEw2Idp+I1QmcB/78G0+Voy9yu6DlrfjQ9sGPxCD+NNV3qoBLhR8gHOkI
Jv3VBgKkjUiwpZsPE2uAcIPQmxFsxYjbTTZSJjb5SnbbLSBu4zYfIRxg4x939sDw2kwbu5bSWl9w
7x4+MwDKOGmh+R8CTmOfCNuas6KkpJNr1+IVlp/7TaCtJA/W5XH2tZfK0ZmQ8T5m5FZEzhbufcLQ
QuS98WyOH/oB43GE0NqphombLkJbvQxy1hioMpYcwDzN/BHNRevpWydO6eowpx4Wmkz5KxA3uUnB
y/2frcdxBLucycfvv7h4eaWsR6axrUj7xWt1v4KuVFUQI4wfSM3mVZXG7LMDLR5LLdlwTYg2jHgt
VB1zunqkiKBsdlpCAjCGlHZYaVpmELdSvFFnS/mygXJXlWrCNLxy6cr5ccNaBiwIqAYdV/yaIr2R
wrxOtSSTv+vJOC1CW1T6F380XDpmzKTbuh8ce2pdyo+4csHxBzzS4QqJ0Fhb3Z9SvhVCdZwyW2K8
CgKyqcGtE+XFjl9CVwGQGUJBhw8btsvYaZ+j7EzFSZiDyS4OUOYidWHG5WM0T/kg3rRvH8r7qdbP
0e2zHPBD16JRVCV6GwUZjOJQQL4wa0RtyDwxtn9sCQARQMMAj9oN/Nj6b3Rg/Nu5rVsNMt6y1Vqw
gzpOIVMXVXOuk0J4JkDqK5i0v6sxgXDmejc1ILmBjj5GjYETpuh0XW0dD1X0BXu6hX4AGxjEYpDf
9tqLaH9PHTEA/EFNQEwkYUlWGG+HmDYrOYvMhlq0SfxZIECbtKr8iiC3ME49sFec769lwzqYzCF4
TlNG7ISHNOB/P7gsdCqwRgBAF01DrFLwSxY8OhGC2CdzY3LOwPy/phpn+gEoqSjMkZZRFZIZx7ed
J8R0Joo1ZlMTYFRvQWaMYyGsVtdv0CB86qSPeMXGiKeY4IqLdIMP5H/N2UgGAV0yTtUJpxjmjAu4
5l6I2PmeABrBr+S+j7gdKdx6k4Zh6W8vu0tvD3tjUtJduwgVXmo8f9RNKtHer//Yv5JwjVrY6xn0
GTWvsMzg95W8ovLVUhNLZBrRkp3x1R/dday0Otcrci/1o+MnlesH0FdxVcKbwIk+STSzf1TvCflG
o4Ywkrth7ho4MFb6IpDGYdr7zZWs/b0+fRBsB5RgAk1O5wNM6Tuk+zwamrk9uHl4myvpLqqA0wTa
eunBwbC2egDPZmX0kMaSYrgVUqs9D0R5jkfagUdbhaKLIRmkW6Ng5lpbUBnUyW5jnV2ybM1mFStG
zb/ETxtrmemlKm4aX8v/C5MsJFcToa6mPu1BmA64l84Pi4HjDhwASkarUtk/hT311uRC5LpS/0J2
jz+MskmniE2kwTW0OmxSW9oqUU/5tGfgeaxxwC4cQ4M3GKUe6y5BWcNwr6G9OMz8MDdDHO2Vo3rJ
dHWkf5oiGtWVULgpGg/dx104Yc5M3prHei11Ao8LqcmVLyIoLKTDpTHb1sBzeUsAUJRMo2Ql7eED
vvOjt8O80EzilL2RUq5Mj782ZNS3uLBFsqZfZtJhjILoda3MZVgXdnMIcsQ1L26r2w+ywHXwFeTa
Jqr2qj+Vdtr0q3hddVh/x6XzCzsYIJjy4vOA5dL7Xo/GCNfo8HaimCRrqv1bir2Re3LadwIAfjGY
erCt0IC03/oVaC8QZs7gdMSOQro0npZ7p6CHzlz9qdx3SQwhfEgnRjJDA1/5hKqFG3yyDK4Suc00
fc1VpiGlfsnnG1s3tqB0P/29J1/Cuog3NiEnsT1Mh/lF0UoOGfkbUt6GvZFJYF0HyPV6/VjVKH0w
4zz9k3ZhWy5y2aFCprapT9jK9xuhG3eAv0VKcgldF1LNvb7QuUbhbcYNqIIU0e5iT1ynBCIb6KX/
UGIwUwUlcVBElVglnV0s/2x5W2hu8BIF6/EE2K4VZ+BwkcPSRzWqDg12+OuHtOaCpiNQ8SWozIG4
bcJ4dQdzrqkED0NmrItEg+etmiCovnmvEk3g4Zyt/ZmGQ0HOTXJMvJZMaPkNxXQTIcYzLbcWCZe5
pihU4FXep5SiMAkA3VabfOB6xjqofhVnikRDByuj3jt38qCwF0gB+YCmUxEOru/xozgBAIgKg9es
L5/q5YnhiMdHOjfatMvhHeuxOh0wMfHexT1TEn1YWFJ7x42mPIMAFvn2l9RSs5vmWlAFoLiXZd5b
+vvp1923a1rIajOS0uCl/ORXTapXK70oKqupIen80GacpY2jsXpfuMvvT3YmfCEn+YhG0scBRYM1
R4FvVWJlbH/coMA1+Vxh3HyLbN9pQck1qra3CR1Lcx+OC2ZdxxZRmu8p7jouzqoWZX8Ui4wDvSiw
7I4qS3jF09nvoFJ1G+jXqZijujI/dNIoU63FdYsDBHCV5KF8MMlx3+sSmouvoTr02LVaxx2hK+W8
JfmILhcRYm+K1p68mK89TXYA++E8DJ2sWzROfvfZFsbxMgsH0ckUmU91Md2GXhAK/q5KqeBm7E1P
g5aSIIkqt7d51XByl0KmdPZCix8cXWXAVmtoNFcWQd0NjGEZ0iFPyFhhstDcO1YIbofSS559sL2l
ypLiMoxiWqeLlkxYYlfdR9vhtR5ShsEEcZt2WAGmfG7rEcSO7mdXaeYqL4uGOrR7Yejy6b62b+ZF
d9isGqKC+Z+dyQpjmY/frf08YVfDGMHM2/OZj64sldt4n+dHtl3pK8cU+cbfhx01b86VHvzpRleg
2nei7h5tzIU8OE8/6fvuHQaAO8MIMZTTzjGsJh+aHfxsMqEBjPCo9r2CR0AoPEgqJ6sK6bd8Azml
UxvSJHwWW12zsgG4tJuOJ16JnrqmC6F9+C+pHu9vuUBFkOcCtZ3LXK4H6Dd3iMDNNDaiyUJWse3H
OAg4M6SB1d2P0bmygU4S7dRNurCBSsn7Vt0TzP9tyLcDBCy3LbDD4H3x+RbaQdUt9oBmktfmC8A3
+E4RC7A/W2FnQ+89/xeLJ5eohnaGLA2EL5GZuHtduYY7RcUBRIgtIXzGNvWsAmYHWnw+5Yrybte2
0HZW/SiHy99985jcrd3ciuAzqoG6jMbqM4TLYkAjQpz/Eo62Z+JEDrY7rPfcm6xiPYG9DgCr1q7h
nKPnxiIU+evuNt8syk1A+6TZrQBSpO5AEfhmZvAcye62oYSUGBKy/s32Ko9jtJ2vHxPKcvJZeFBM
CUisUz5sNPahG8+4HOHU6aioj1zDyVgoyYvhj5oQFFQ7bOd41AjoT88JLLBTFJLBuxWUeFdEltvz
okfzvOXVT0OM9uNwYNmyV/677uwEzH6Fl5gQeuBFgpiO+D/A8QzyGsPQ9vXl6nEAmtO6ISuz/Ggq
h2Pkz7bnr24jDrc6Eh+yCojHxpHLZNjIqIl3NUcXmHdTfzRkYV6Z7PdFATeI7msTHY9hbGIuq5ry
zaQIFr+rsPoQXTcyI88GvWWA33omCc4wreImb8/lt4itNlazL+TaG4YBZgE4o5IKQai+8FsknUNg
BWDNN+bwKWz0jvLzbwOn+wPK5hlxfUlqQHHvbinFRKcGOpIa5aGGnPxKPiLtwz7Vv1GhNr9WVs9c
Nv2ki9uG0lRgCy3nmFymioUmNkl0sTALGeNwhhpSZwd5+IaqChlAWYlg5iqyBK12ZX2fcrdZhNVO
Tm/eH4mfn9ROBVyipeewOBdlPKcDsUpfzLGmKi064RXAZI325tO2L3MqJhr/hndZHfAkPQHmxIfE
PxINfh173DgNrdk32VsRlU0yZGsxEzpPvLHbdQJ5vGo+QrS+NOFqvUn/Yjty+ITpNBD0XpMC1UqQ
pbn6lXnmG5F3UCXE08UkvY4DeDiGnFDDLDFIe9r3Y4UXQ49ygyzYfh76yohEfOpOGu7Tj6T4hDVT
b31kRtnh3FhzDMwpwjbPt+GFXxbtQ1N45gHnuiKvv5l/nZ9QdU7SE+y02ZEnkV9ZljTZ8HHdfU0M
25hJqSR93jZpS1tEvJ5QGY6yOJl/LYJrarpsjT1D6cqJ6qQZgrVTFWSRIU1ZDQP+a/S8Pva0fiAI
fAaxX4KB3d0ResvEV569/NzDZNLwe85wnr5bZwhj8+8J+Yrozm/83fzYplcB5z8xJ+tywwvTo1rw
1SW9sY02kfeqJGsYCUN0slIZImiXAxG1lwysaUTFaQhhGV6zG1plrNEHTk3DqtJ3U3d6OhfhgxNU
cx5a1tOsjaNm6Raw6LNIz06NRCuJwnWs/Lom3DBUTd4zqqISB/f8Qc8kTug0fcQIs4AG5bk6OAvj
1PWCZdWEZ5VRCQ5+1aiu+ULmJTlBxTuJqpvGSlMoGwvGcUjL1GwVCWV24Yuq/xQVm2r+PFyIwqzR
FYSsmaTm7dG9wzS/42SCQda4v3ylHIkza0GhIcwtmzwvWSZ60MRYEuuyy6d6tfntHV9Z3FZtQqxF
bSX2tND2AS9U3t50Rn/I7dH5E8wviq3240aGmjtNg1Tt2QuIsidujSZuDXAu7ofREQUpulvb5Qpj
HLRcW8GC7xDweZuY/DY7xLF2NiaTwQKQEIUA2wD6T41dJCzX4D0MoyEC+oucf62lWEgPvgKZ72OX
g7CUnfKkblsWjrbKvs1KizBdm+bR5iavKL26WvTdGH+zUjgBZFDB+WaJ+z00l+Yqk5RjYm1w9pLr
PnKeuTTY6KeC3UxPnBTmv7nE5+1P4ph+IQ9Qi1+AxA0R+ahYGFvVzcl7X2tEtAe8e5SBSQKxOvGy
B3QvdHvXHLfrd6ijy4qdELrQcfLlVGFF8swy2fAujIi6zuR6IvkAuUvY1OLDEQr+a15hCrPiehWd
O3JR6Qm2O7Tz18SMR8Rm27WQG692qSSExawN5ENcUKdKQjUXDtsobcgdf0JB5KKpb1NoGbeGwLOr
EEHysZu3QiG7Sq8TimVaIrvkZQUmjaZ+tn7KR7ycrrArvGPkYHto8WTQx00jDF/yFXFvOwSyJRiP
WpxmYtN6VsgyyFOR3K1a8bN1hh61AINdsr7g/XLTN+UbNtuSQVOPESh+HRJhN3bUCmSMzOjw3uD1
cpWkmOjKR0xsaTCUlbfhA10HXY/CImkyIp7JdIqC/WZipUnPEUefJuwQBjYf+JQJT9QN5w0JWvR/
jSnwTv68dLxTPzZ7Re4sXoohAnADveun2SWfPRn2lQDsGexAcz4AVcF1r+ypES1hzYU/jDADHJut
ZOu6AAdVWjjqJAWwnuRpFdTqfkAxc/mLw/MFp8rQwGTpvMmmCWyKkf86YQLUjDuwO1KmGwkMpcAF
mN1rqVm/CK4QD31OGMILfkWPPe410PsE8hUIEJlyGaQ3/EyrA1NPpgfQffv/kszdfgPwCWWm1k6D
L0QMXYHNfBBebPgS/4TOi1VQ92HjYi+utqGWGn38dj0hEvy2Zqd3Wneqn666uT8fnw==
`pragma protect end_protected
