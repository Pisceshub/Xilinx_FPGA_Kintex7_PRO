`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34880)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3Nxgd26/+Ei/r/WT7EdxPCvx4pn6JlvOP5PB
h3zJ6hx7BRutXu7DahSdf2nKX100c5VDDL/OvWRFYnrR4tM4gjRDAHZ4hCMgMDxlkh2nBUfLz7C+
+N68wH+k5oyLxmg3Vn7U4G1waMF74kCOvAXflV8pf6G+dkG7BtKInH/Rp+mrIOAda+DsfvLe54D2
gfY1zsqLvLu8ZkEFtYEPq2kjUCk3mYKeSqvenK4zFRsCsHZMuJoECVD4TDjNfKun2YfG4tfxXsiv
nIDaOW5t5ecLGOlnAeIqZz1hi7eUoiFGnnKmNbNCpxdZLpJU32U6063CEZ5GLrCCCtLbA/2flBvO
sMeKuhby2OjsoNGkxnLk2efcGvNCENq3jPT6dk760NxyAG1+nqR1aDF6xSPxWIgjOnxQJf3g5iKK
Tc45Wo2hRFg76d6TopXIZLd65605RzQ7fUdXSr8P6YEejEQgETqvcfNDc06abyk2aF9qWu5Mldjy
X1tuq2gq4vn95oPBzFe7exO5tCKWXOwh/R6D3/8Mq581fgcSpx4zSg0HTTALk3XLmSENo/PZovuG
2/ImUD2zbYe/9e1CUOEf3LCB58sYLde45gwc4YtNZEXCSlvuaJlqY/TfmH7B5G8F98tomDjPl1Ad
XLPv6wFP0hxIitK+eAOVdYJWK04xkBAitQl/yKaXcLqjUaOEwRgmBiV1IQw4BjtgFSBzRIoBQVU1
TR/Xh8k7QdBRCYpsWhB/gyHoTdNSSsRtleEIMgb2FUsKg6bS75H7UF3txjlATBUi3T0uzbKLCZBs
Aj7QlX1NMuAW7e8NtNgRYUWC0GdTr3/Mzdf7/RdLPs8YXF7npb0rm0Yxs3sVfjWt5CGWdW800zzV
CfVDqbAd9CwZDuPzX6YU5ia3By3BHfOlN/SML97SguCA/V6GwEpPwkY6hgRVwE/LE8cmpWq1ZZuW
PZ32D0eTK9wasap+50Spup3oezwLL3biO59bSewk2BtThkYtaO/Fm9yvk1PbXp9U8Mmvet3RnJyY
4nZdsTBBzjbGsAgR1YFAnp0jWTesBskmlvS3e8g6E/2G2hDQZzKH3z7ph/bd+jmR1l5dClt2wOCw
ZHy2+6fEBO1tZniXnFZ+8ZtFhE6NzMNW0fUeuRZeEQbcJlxVoZB03GB+GTrTFCFcC8wZHTH5mX9u
62wBYL/cenesW74Rlz6RPpZMO3dugz0x15IS40U2YsW09mWUsSQ/GcdN+qQxE3H/dTQHirnRxJPC
VWJUx7alJs+f33wK8StlLYJo3cWGykvBJmiF3q8KEitU+GnETMZPDFk7ElN6Bog/I0tj5RlTIJ2+
x/dtFQGpl3kXdOJpNjTHACZUHWHmudNIzT6ETw3HGrk37LcFfwUxVqMQvmk01bFAwSJcLK9FidVU
goeXAuFKypp3hpft+UvlQ8/085YDzQfoNqIsz3uFQaVHOP7BoxmfXuxP4IQwntXFFIGKUtW/WsR0
L3e6B6+ezDwkQHxX5Af9ASo0caQMkR/2AS/IjsxrA/nwlUqGo5m1gmvOSS0pi+lOJCeRctvIt6vX
V2KCQbLTbXngsRoaVCA24e/DIIP4UgnUbNXQv5PRuPaLMSExTmqB6dqEPZUekdKptmhROUh3/509
jb7zApZUA08rsDwb5AjZcwYzUjFg9PgfRhL8YBz6FJznxVKDOLdjWDYj5AD2pI4xixK6VNBrCffd
eLM2xvbUS69HVAEqST4m01+wzQd1KksJs+sO/9sBX/XYSsP1BRcpL3u8QOJS+n+0jTSKmXsjpDCO
1PFVpJ9rTmzIFP285c0CG/XqS4ZKHj56Xq7yAQwBZCH9+d0Ro1vciN1+V4SZoRyZNZge+MpuNYKj
+c/f2lXmx2aVCkcCUdGdt2VeV2YRgktc7YOgPy+/gsw59lin/NQtiKo2OMELeBwAmrWMapOPM1M5
4zgVW3ZmxBo9hc6ykVWAIeBecHbBRuf15TbqcSiE+G6XnVRSpzD+i7ZZpfvcHFHCn6BZsLs0/lHW
AzvXRxjsXJ6/baIEIpqzmCxPDdg1xKbleuN06HcCUT8ejbEA8yfwX6VSXVkxjaaRyEgTx0nJX0He
JYNX4t+Zvh9cDKndVwJIdv8ZT8KEVTNUGSo6MyFsKPiAJEPfKb8M3ws2qvGjrz/F8XP1RWkjFpgy
xDF06Yj/g/Hg/mzZindxvVXvlQO4akzhZoZG183PsuAybu7U5/T/8J5f0/xKdME1kMxzJ5dWwIYW
3Vhmi5QAkyuTUD6SsaJ7+b0bh0eWvwoMX0TO0wdBtJcN1FL+JMfNlgrWKgR0zXFZabZmYBbCTp9g
rQdEytAS+86IgfplZuE9okYX+9TZubMI8cujcw+Tqlbkj4IHirQUZnov6xKJrZ7BICCpNcRyQ5Pp
m8j0QTszd7Q1kSYP69vOlF0CLUpDH/IicojWl2jRVEIZ0Qvb19/vW3Gpf+3GxLuSOroCikrQRBNh
Ej427VPykvO9h2SHZUscs0LgY6WTm3n9PcUHmFh8QNAAbRRVUmsQjA/jA+lGt2ExYMO+ebZZaQe4
szIoOswJ7Anq78KiqaVFVAzl3nlJnelNDvQxdtIdqAZGuxucpLPux7f/eOwEWVcEk3uxGrfIwZuX
/fIN5L/zjo/rF364B9Lv2WGQ7gHSvGFJngo2J65JnyXTda9EKuJmB7KCKI5ZVlgP77MqogX+mb3t
bzWacVZQkoFJPczKyB5P4/p8JFrxhWHmStAgxxzDgq4ytszKhBU+0T/uTUHgwP1vmycREc8WlJSj
oOseS+XeTLK8mnhQiZkgB0dyztA1mLezGJApYPEPnLc+/nC0mxQU+O2/BZ5zIAxVKDtQ5iPmgZKs
idZxAXQvrUsBN8HWFb9LECIGRcHerB7LO5HsZw3lpLeI+m8DGP8cFm1hwlNdwp6kwtya2gXqtYhc
eGqvKwKdPoVvnHqt5ED+LlrzTFxbjs8TFSr8bFu+/FqXg/gHbWPOTFjKQljMs5P06zWhzn/MesQk
y/RXec2Ug3Zt/93JIZ57PyIbiIRUav93QoxnzMHQz/a10kJgkmuR4FUwxshlcmbqhXeSEJSlykMl
bXudrH+2y8mpjrcNTTKCzx+6FZEg11SanyuvuoCBCehke3Lzz67tMtTtr/Rf9xMSxCXuYBtpoykI
aRFLjX+BIWEVZvGg21MRhvmvD+ZAw5KUsbWkYoJ/AZ8rcv8QETrxpOXAKJj4jSyZV9lyyawLeBfC
4Uot3CJGfy+wYC8ja7lF+qK3+Z+tJd0TPUnWTGTEW/5x2cpU4XfR2OlB7AOf3ACONfYVCz/cMd/5
kWGiIXvlU/EyxehIU+6gymJ41xl0y+EOWZ36qc/mfVAFtLtnkOpnA6fxcjPuas+gPlwLFG0LgCH/
C4iR4FKxbePZ27PQ9nrbFTKCXv+VW5FwSZvzuJ+1Fhs2B+lV8XiwM/0Fijv4Ucc6MGX5dgm45/GF
oJ6X8jpCtAiojkfrHkIvXRWC3qvpHSF5Ivl3lsf+2WkaK5Bcgz5MRaBh5Wjv7BSQQ51Mukh/F6Hg
siCiqg5+CcUcz8+rtn7Yv/dFEfJ53tfjXHcnbgOX/hFd73+y0kR735XuAD+s7LwPKY/2dyx3rxsA
LJOsr/3bPVpRZasS7OuCXKZ6WhNOuW7uVc+6xyfkMlbGZgB4xSsMRApQc8rIOpMO8Xk5VwBt53Jr
0hAT/tEKHWWKs/x9I3rTG2g1zPnTYIUaF1SJ/NbFU5Ua9+hr8RE+oKZOC2tTOyqsyGeoImGItwzW
hGqCSBPMHh2fsgYvlZUxBAcAn4oEsrUERnI/2qj+gm9wauz11anL3+oV3SeS9c6nBSQ3dObbGWMb
NRVeoQhrlg4HYpVr6QPSEgspURwpnzuXPANYyHIVPeAL+q62tuwrDotJXJ07d+QXQ4RC0bhQ+ZCH
6hB2xlwlwUEuk+5V5M14W3KjbQnuRC30U4w/kmzrAOCBfucxMuffTdI1SM0+xkQ9cX4Py5DrHBDg
Xk0F2LGSIndMBjmUe9juX4pwCQQwm31HKdHX0j4kBYEyEUOinxFovuNkwW1KoTw5/omXs7XSJp3G
NLN643BBsQraOA+Z82T1Q2yYUrx+S9j01LuMD9z29MZy2rrF7MxQYpA0Twdjo7GcMwG0yJ7FZ2PX
IRmjcwXMS6AS1oVdZ/KGrLrPVxQzxIYuyv5jxktBd3MqepOWGgcV1msEbU1Dwb6YBUZclZ4dXnKg
+iOFJuby3H6G1w5Eg7AVBUADNJHfTRBueOkZeKSAXrihNY0oprekHhGmBVtzNhSBGtLSeZQYx84Y
mU0bzBwLBokXm56iKysHkNwQTm2Nc9nS1PRVzoOqQbe+oY75DGaX2wT7uijC/tBw+SgqeG8609J/
GAg7yevrjxKAElbp7FDlj4lM1uuV+RJFrDfYsnfNoY9bVMnYgIRnrllVWXLCvEML4ElzL0ttxySr
ekhSm4q64sGpEBCVjZzWlN+SnthSyGA8wI6ghacQkZXqY+hfNRzRYwpsyOTkSl1bHPUUhxnr9BuY
LD/oN45xISiQ0HPHnKeJElkmCOeDcV55EeZlTRO7xaQNSHW91lCWV4oVEGSFOVCYORJQ/dtIrpZ9
TNZNP55yE4nt/kGb7AEYCsRER6+lRFhm/Dlh3P0qUHsVeV+lI6KcWuYmf6WNK1yaIa+Sph6x2ngQ
Rb6scS4mlQ7F7q1uCZ8l6NYEc4tjtftaAe5V3SWuiTXpCtJcga7zUszHX+vkBHJI6nBDfMlma7HQ
P39teJtL49CCCK7yqMKi50/V3cytq6lq+nDpxuyT4B1FzTOvAi0glrZ/gkcRScBCtCtETiXSkd0n
FDTXSolbn+3YqbJyLqjs/0rU5GLxDK7+QdK6tJZui0QV8SrT+ohqRItYYPX6HUmR9GcYLJ/QCzND
CTfDIBvE+A10SWrZbFCci4WSjzih3AbEsb4anarEAj0oiBBChb5xZfKv6KPhZaP/I+HHymG5LObK
kkjgMDRe4SXJFsrLigIHoccfD5xHbrb63uwh68x/iggDpar6iKu5MKgJ/wF2iD/bfIKczlgwd41B
J5EhDX77XHLhYD77A0UDQPDSlcJB54wClS3qYRJmpsqtnHSDJM7tAlBFeYOdJ/wZXbCDrv3iMNij
MSRtHOxKJ+mmapB3Gj7JGNWJ4C53AkvPbJScj9Eywgo0ddcU0Qz/iMVMTq3ozaayorzHyQGrUeeR
0zC2fzJRupsuoIBYFv48RmmuBDCQ0+7E9reXJr5oV7MaDyOxMLv06UW6IFmGmm7vUxBs1Go4/Mmm
OMYux3wAfz2U1FawFn9pzIZFuALmsKB0WE7HEh8hz1RbCsiBCveCIpT7mAnB/TR2L5cCQgln0JL/
g7ougYhrIomWgkbzZPHwvZgrD5CpiU3lKL+3znG3PuU9UwDxrsJfFIhZX5qb9FlO0F0LxkMtuZV+
mROMlwD72zzeSZ6VhwT/OZUeAKxcICfzQpJS6JZ5QWx99klvS2fuKh0s6xa9hpxLQiPRDiY9wgS1
TIdFP3CaTMW1ZiupTKr8AFjG/BaiPlIEftwAzwWrOUt/WHL2XtYysfdI1snd0pj3htrgXeXTG2b9
IhopQA1iCc9cImsn4NQVW4QRQE0Ma/FpgWN8MQ5xiSzno0kdNapGOJoRuNFc3esDgeXwisKUnh2e
UxfHN0NfCTlAL2BernjjmkHuRPOXNE53NHt8dPwBA1Z6QEqqc+eftF3h3og4uddOSLr4B8jy4IU8
AigoxFSaYt9Vr3Zofgjn3dhKll7jRkwEI2dED+gIkGdAMTUIHOjCiM+Z1dUEP3d0O4SW3hg1z4FR
MGlhM+kt1ze9RooDE68FWSkb85E2HCr61keVdY86biyXuufWardVKj1QKAoCweXMO1MA5NmLeGL1
QyY2OjPaVEvFqn4I611xoOow9MEn4Hd5d15tkOTpyneHgsJ48vI4ApjZLMmY2BUCfBPvVj4MnXiJ
8y3ZBVFibn0frxQLTzDjcRCKNe/u+eUMccBQfVqUIwYlpBPF/9nLhWIGYTnCXvcfUBCjhWobeflk
NdQvZyky1RjMlBAyyOfHUFifT0SJ3e4UH5Od9tpX1vyVbI3w9dIq11dUgBkSinKP1K3UGbPKnRrk
jfrGTduCZiJoO/RYwNP45xkvyjBMSYwqMnGeX+jVrRiedQH61ceo3njqOa/qh44B2iG5Lb/NTSU0
WeCxibJC7s8PBN6SrLv5uYyjuqksaZ1BQwJglpLiCsPzYwxBGwNf24Q1t5Nh+CKmaOSRNr90FHl5
EY4S6nzT1URdnQSXJOTT6L5MALBcwqBzExlcO/7tDGMB4E4V249awlmczM28JF2H8svPM9KXWg5q
UiPPAhUNgHOLAlJHW7t+W5tmDLz6HSIrvur6F/T87yDWzVtufYnOCVkY/bEUM1F7jVPKe+58iBEt
t+fOVvI5056qjO84XmLJNKUVtnydnjUNoGLh0LBHSGGzJkQd30mxJnSQyFXXXQR3+gBmBEoOBhhg
crjRB6qW+gQhtMhsIDQlFkkBeQODBbYT1t8czOD58VkaCJ2dpGh+588WBtKxr5GG3tmjdBwXjgDO
cz8MFNmJzlyWuERnlWJWn2KEPeMuG07dCV6puXZl2/7yjLs6MhAbJsYpT6vKfPOAmuRKCw3EaE2N
mGftv3lzpCELXqPNbDg/XDtw6FcpRi2buMbsD9MPxB43NgkN75HvgMRV/N8OMStrKbnh2a57aXF7
eUT2MaZ0kHd5GTPg8+Aft9dGAceKangKF7Unu1p2hcSzDOlJ3C0/G7m4prlhq205w5Vzcv6TgBxk
82sOYqmKwfYLKtlpCK+C6+ejKlnDnBi44wayVpplSHDRGLA7P42oiW1cS1UMicip7SGFh3+Fvpjj
g+BnMw4DvIsQotFlYz/ELak+L7qf6OLPNmw8G8kj2guf2ISzyq40xDtjip2tAf99xz6tJslbK+qS
5wYsACuNAIZZRKEjLZx3Imi76QRTtKJiHHoP/F+HLYMRs/ENKQw2KxyBXZ8lzYt76eI2VpmVbvtD
4mq3/MMqWPjpTLd0xEZcCTXhpu8WHMXxaMGJxFj7XXwboqsyHBj0pkyKiiaOFvpLMPfJ9g8JSijL
C5zUd33DEhSVymkXoiq7iwB+vbiF8hoAsLv3vLL6/8YVzPVnpciFZsFPIleLRZrHbWhEAo/x7Shl
Xy+65u99D11V3uBeaY2fZAMMSfN9gIn+0LLqL50KFbTnMJzXo5HDzj+AihPLpwrWBZXZnRF1OibZ
pfmZkfUcxUaNYWQ0KuZGh6137YuCgfjTo7OPO/UWYZscBg2TEQgJVFMic6t0an9B/SAXGdmudRu7
5YmeeLeY6xlGG3xE/B/ROhdUaKn3tOriNjIaz46RiAl938ptq+CJO+aFUNJIdjK7OtQ7E3vsF8gr
9HqQ6ftHLym1zpmYRSy9TkHH6qml/zGb3llRB6ogUFjXCED0WTcl51lAxKbpdV1HpMwnr4lu1o4X
7qjJMmwNuIdWjKYrsaJuONzcP4y06eUYH8CbJqut2Csc0EDzEaxJwHn3pRXwRM6r9auPsNDJCe3r
Gbk2O//uqjsbXDXdSfLRP44nANJAuPzxkb6ORmBSWokT0N+4uAwMafgX58pYcOEuaO0bZH8wT7t1
Ac5COs5lptx2LSxQiVD21I6FRp6cHcrSrXtjAySc3wXqQb88o5YdXWe2l9LkNPKQlRFf02ux/NmG
8AdFONQ2yT37meQZFwYgUHC1Dlazks5S2OsXKw5/HympwoXIEjHf8RCfJqt9myftyh0XhAcZvXzu
x6EvMGb0f7EZnyAbvxBFZuOSU0Hl6g990GeLtjmQD8WbKTICtcD4FWc7nR4HtzztEveNktMhh8rS
8lgUU805lvQt24yXLe024v2iPMitmxb115thZsuHYDXQAgGKtKfWg0zJDH1dunrbFIj5CAAaIbFK
ho4W+gbQ5ne9k0aDMvRsMYeFzoln1sySMTSLtZVBt/Fa4kD3skBy3np1dpOy2EEMhIX7ns/Z8Prk
TfHZCkWttkooRdrbE6Sjjws/QB4yUcnhw1wraMW5rxRwZVzTieirrd6msK0GFQNvaHuX8QaFas5b
178WRg4qVPNJ/zbP+iMn7tJonBrYd93jChN81EzcmuvcnKG3YwvZan5bt1chpwti5xd3izCNUSD3
DSUCf2a6q/IZU3gNvQ1ATwDj8/ajNb21jEv9QD3XyttKod/UvMPmVNIYAwZg3nIX5UoQX+yjvFq+
W4N85yBcmktJQzolmiL/3c+gzDNOajMMkmX8z45M/J3/dopxwhu5uhBtTugJaMPWce6LwHjvLFNS
R/8V+VwEdIuk9b11lvET4lsGgAztUK3AZ2lCNlX5R9v4cx81HRMn1aIWKxp5ScJitAmhAbIZJzOS
ImbkEVXzNqDDvoGT4M+4QiiT4Gp9cKiZsnOShLBEuHPqm/8Dgiw6n13/EnP9nW8pfE/BnmMYqYYf
SQinMliTyNTT7Ix5ns6VPgwz6AXU0FV5MFX/Qz/QSguX/HNfgGMIIoIqLlZZQO3ikrmxVnx4gqM6
NFzkEj6dpdveHEffsXFl/NhYkUT8FGcfrrnGj4ZYm8wkmzFYsU0yMwv/O2xc39yfuJu6Xe7TJmfW
10PeX5+JAGKWO6T0yoNj2+eXpJrJK18EWOm4lh8EKDOnabFXBkBVPeBnk2tfrYWfgEbIaXG0UpTQ
29nxa7TGr/f0kJwnT0c6zagmrNd/Jvig7la77FV/RTwfDloQkNeqJhElWz1VDMuAxDnAk4bKu6VU
nEMJF0c1SlWs9nDvfy/emRYe2B1O+8CQW3kCUs9LRSWxAyxrUD8jVvPI7zQzDgS51d4dQBTjaVY8
Tz/qQXKbZW1bClk2MlKR2TgR2Au/pnavq7Pia0s/HhRz/6t9PDjsd1TxRudYK6nNAhAl0Px6hfc8
YzwOtLCmnY2mvyt5GMWnrwkjYd+E/uO4AqWIt7DMPnrbO0gWiDsrlF/kMszaXM09YxYmyKqz54jH
lFPswvblrttH44mzxKuV8ZdGCO0BXToB+UiJQLLR5xGEOwZZ5CSx+BJXzprZnYyox3UzY1n9o/S9
dOT0/sFR+/S3QyTg+n/Qjeh6qChiIuGnVQCPPQNLC8hAs5u02ZGo5MQMBYFSkIo6tMpuSpNvIHZk
+DnMT1vxDQQGWuEbDFJyV3W0aRZUjBL7XwxTJ8mFubSGrhRkqbpiIm11ZWtvaU7wIWOJzl/fR4iQ
SyvcUnCfFykLjgNGn76KZg73Aw1/w4Auu8SSzQliaTbTFK/HSbxFpvpXmwWi97rlUckexg+z24wr
7GQa8lbG6xjXmZzzZ927mEv7tYwlakFbVrYFLK8DSh6yM6e2zGhVTZQUrlIsLWtQuDpQ3EFW8FkG
IE4noFXBa/R9ZaDYKYLO24wdQRyPCDleWw7+zhAEQ8UYsXXa6qF5rVxjtXD2ARcnrEpbLlKVJvsG
K3Ml2J3MaCVqNboBikwWjfsBl7N39pv9x8VcM7l07JRocP0hJvP17qzsnGpBCI6mfBouVnOeHKTj
M94e5EDXuQ4laEWm7q4e9uCBbcg6uh4Iz9/gFw2rt+jUPb2BEBG5z/tG092axFxBqUVEyMob8mQG
Q6UfJApp5pygQtYtPQmIa2Bf8LoOioG+tgWd/LIz78G0kP7GszBBpz3iAoMyGJuWmoNr5y5O0hgG
spggrBM81HsPCz7VY/G4Xqu1XCPbT46aPZoyaettThX8s26kbkQ0Hr8UnQlp8uiU2K0tgwznNCsj
VGtEhwN9ttZQcyFazVeJURncah6gLTBZ5uIrB+nwQyHJL0qpD4bvQu8TD7o9zTQrTP5DNhmISBAW
G+DA4e3wIKqJYt2CGyAwaupbJcnXxK8X1pLf5Xsx9JxE3pPDq06DtJ/vzQ7Czn4wrrx5bPekO2/w
x+GCWlAj1flvJzxaNOmlqtPmkSGDNfVnM5APOdD6JBExZ/gE9Kqs2W2TeITBFXJHGdKsfEwDpcUu
1mP2cGcGYc22YTpZP5VLSc/j5FnaEuz47E5SZWQSBeYf7WYNJ09WnJBCtn5e1ZlFRdAVlQFS13Re
sCOL+lZBvusH60lTLv0TExxvyovDZvKVzSsI1itauY2bL8zIGdttUXLU1JbdkwXyTfjWvqxsQzcZ
mWC0aKwexg5fd9yfdixUcFeL/I35BrxAht4fnIkw8xo9jnsDn/VIkjvIx3O51yaCh9KJisWhwj/B
ED7ZTbQOXhFm+1GJdTu2V/Jo64b1SGFwUx6pn5ajApYYDbHb64S2ZW+xyTBHz94F4zt3svAfLIzQ
NBYW99tg5qE2aombfg2TnRcfu4dJ/OBlS1qDuc98bMOOOj9Rv3xZoe6eZjnI1ZgAx32g6asfyyKx
1fDpjxhRwkIWFE+BFsc/h3avGfnnPJo+ewCIE0T9zko75q01Rnr5TvhCo6hHfTUBPjgyGjcU2RNq
iLdm2E5ZCnEwS8iCXVHp3NUrHyn5eXem+FlJuosjP8oUZBTcEkhiJLKiV6CyxC3EIlfFP6yrURN2
U6aQmhlsqZ6Qzm8t74vLhC+QhWkN1DB6OPuL+FC7PLVlVLKATvZnd8q9ctQ3Tc9EUU+9jjcT9XJu
9qEYXt0NuyiJ1tgLVXZTN4t3br5GMWI/yGU9ZCPtBkH4KdjAJnboGUeE1DyPKQLgk1UGtsAvqUKm
7P1JksSk+4WEop33OHxy+emNXvUIfCS1s7c7x3MCx2/wP8ENIZfBOKCM/oMLj2HSAlJqCD5dLIpf
DGpPSIzhXoyggkjk+cfm9xDl26SzlA4uLqMtakKdYhaF5deVXpwawC35OAoSB4GIan3NfRzduKDp
acKpVjzrf6sfYoiyXQo6tF5dz6JCgwmCLCl1tkl6tI9TySI7opOyEMRyTbePE8HvqalO5BfCOKUp
3F9ZuMKBnD/w0Pb2b+cfKtXSkDRwIySrC8OL5CL3J58YsYgvXmIfZXHHVx++NBH1WqeX4qKvtfWJ
rFP396xfW9AmtbRnJGLZWvozzZj7kiM84Z/LGQ2C6yxQNxw6HRPTnmGUp8o01nS9NtBhVrA5mD9I
zzed4pqpu8f6/3trI+yn/bYUIO2Ikt5bOrXo1raKkuO6206HTniM4AMyP4xZh0VswKpE+vGjsfp4
aDCoMWim/rxwNUuDjO6GOwKh490dPV9y0yoqxFMvdnUmvDSEUmLTTFdiSfBtQ9uvlmj9b3qdnES6
VVklxrpuXabHYNfUkfV9Q1QlfEaJwMd16OgVG/FEbRp21KBjIHk2bfKgzvsmjJ3XIoJQqnqocLM3
d8lgzehWduX73UV8vRsy6W020wR8TZS9S5csmCL9kpGhmKeS+mATfaQv8njfa2Gpq0acBn2slmEC
Sswq+rxvgnf78tJWIdunyjSwtG0gZD8fV/YZBoz6B2r50TKLVeZy93L8sITATEg/AwAuHEJj7ELS
ZOpzgXt5wUsOV1fpmWfIGT7jLBW16geIou8kpq1xfznlNU6GhZe87mbaZFZE+kQyW+5we9Xr6oTd
vdu/EEqrqR1wWSKhM1wWNaX945KnrsUPtzuB6BrvhpC4hp1f2837DAQphmjVjGLyUcdbrWPTqyLk
Zj2ryBTfQXPHMXz2/l8RA1N4S8zX6C3Bri62a9FDSaqcx7cQTJnfDFwHXh3+/D3QXIMCQeB1arWA
sbnGgG6gAMun3kTZByDXh2iuQtQtDiY4o7JiA0qB1elPfWAkKacBGGbhxoUxDaAB5cYPaC55RAJx
mN5VBkrEKaTiTjFM/3V5htQygqfMetyw62pWMC3eizZIUAMjwXZB/5PsPu2wBsDZbycCQ1o1hEBG
vU4BsI/qjuedZ7DWSlhToYrSBioZBdCBv8k++rMLGsD3MkujYyjQXO87rAmQ7Y4cOHAlsy13vo12
q4yBRlxn55FbNj0F3MquDw7vZu+o6GnXQQlwkLQQgEzmbMevXAjfVRSjN0MiMf9zQ1zcxuignUh8
OB2UbBy20A1N5IuFKgIAp3huaS/k64I96sL+SKNC7mDkGqWc3cRwuNPhE0TMwjEFnscx6w/mZwB2
mhw+kbIIBPdsC5KlQwbZMuwI/CfN3I1Z0MqaD4Wh3qylHY7gq2v/Iyyjh3nmK0Mc8+nottKzMA/m
WeMmmvovDNpC51CooDE3eJe4+TJcwGqqaw6FUlOt/EO3bxvlRec0pLyEjG+AnjoPQ9MsyjF0OJ8T
cwvRdAA3LvYx5xDW3OFV4JzMq91dRFwbAb7Gxnrz8jwhKEAE+2CsxnnBMNP/CDx+88PJPUDR4Gqw
TUTcVtq+mWGUPEVBTwOz0fTnyoIUe6GvxrQKWgbd8+auohsZn+e3m2Iqi+SmYhXSbnzk6gSfyjHY
u2YerHVTUg5n54+GXnB1Oz2gz+NGntfUjWjdv1icQ6Zsa0Zau7pLXqTAJK8FXm8y3xvqYnpZVvv9
Z24XVH6l84OU+W67fA62TdRJNeGabReFOv8DNGgwtNUuOz7NB85dIOEYVB8wJtyfjYhpG52kUjnl
A7CmZycY7OyyjLiIMoN8w1J8EBgMjPVqjBHOx9J5ezuUvJn1xva6qiqlQLgcli2U/TFzIOTdkM7S
k0Y3kTI5VhXl8lxcg3v1bnw1FAHnFpJTD2nQXgUaIkmh34nQVpNt0exunesTSjilu4Uzru+V69eM
BWUEemxPKIK++AFJLKbamNXYHpWEshjyaUht+s4AXim3LSGkw8g0WT/Z3nFFWfoFck+Rke1s9TU1
OC/8cg7OTFiwMKVMsIGFbiO+7sYkMSZU2cEILgtL7qIja1JKaGqJ9D9OulCGMsy/A6CMPC7bxPY8
qUnygedo+ZIrzeSuaPo44sdG1h2+3pwchAIZlGFwDdOgT65KQkaCrNlP0j1cYbgWU7HOOL+d8OT0
mcTTR+TUOQ8StUubUhhwCUNTQ7gKt1xFf1Tj82beIdCa2kRVZQaTIYx5Xl06ySmkDEHxna7tulID
rTR8ElK/0d7A4dImZRVGuCK/cLBMcqPbi7byGrd2UpzO+HDChtSA6Y6Kia4Kjx11dziVFz8q+FHR
bwLCCfqujuKtaWceQAVHL65F3c0TlVx78w9RB6LFhFkBr0QYVTBXyj5aUmxiY+oc663HM6etIX7b
55zmLyJnrVHKCs358RvD7+81u5Az2bVRLZGdtm+DGBymGsFRlqD9br00JNeSP/XdM+0TA0JpvJf6
Xc2H/r2faoNKEai0Cax4CCeAWMDK7+qhtJQ026tA10rB8/eXvhKpLVyXRbyElgiVdzsB2haagqIt
pMl4ihZVSezFk94R0F4UDl1E8Skqg+5+KaetuzRcBlwOktS53aJHBvYkfkG9sC+Uyyy+B4F9qxLr
k8n5BqYqHQwSbWdxwztjvRM5/nZ4Alt14PdX5txnwXPWa+s4ZhsVY4XxMV0P2M+btnuKt/aTgSuL
zlcFusOcl3/38LwAeq+5T35FpcSIXbIHrl7lvUnBY0CdJeRE2HK+MExuBZBxD8NK0czKDQq1mF3Q
qphEQ+XshAYNGNPIZHuueOHZTZhc9SnX0E7Ps/gYxabdc7AIF9mUY2iYhPGY9D4978vGX6AFa9+g
fGAS6Y8O0X3FUESBxHU8yYFD9t0KFus2cba+U3H4YjedHvKSfWJLpgtf2xv9gCE324P0vCq09n0m
gxDs32LFtykyd66l88yK4f4GGS9FhSBC/RT3fm/w0V9XzaQ8ATw8Ryqm8x6azJSfSv0iF/rwJmQl
DbEzYWGngb/l67o7CznzaD3a7NpZRgRoduUO4Hu/pANGrQGOAJ0wnJ2V8f/JAs7DwprvYd1MtyTI
pIn9ba/cUDywp+4qynsVkBn620nPKMZKLBf+7tSaosBZ7xqHpnOyVvmCE0JJITHLyg6Id82rNdiw
Rxzl+SkRoJuJ7ilItjEfyM2jYCN2QkQX1zVDbgIdD7j8ZXdZlZPsb9Afkx3i4H/v+0oh9axqv1EQ
2y5Gy/EasZ8upV2tNDPB65lXYJR9bH3KABCa+rcnZZaOMZy5xlZXKSbpBi9vYnGwhx5hZf6STMIn
k+DV9+/qb+bAxeBcdqsV8mfMLrjEBoTGw2CbrEOoXjrDt1d/5W+ogw/sVpHZkBLOAG0a2YfQ//Bx
4z021C8jEgsIvqVMOk5XWEHrMIcH2XpnZu7o1aCrUTEkJ2qV+3e4agTk6VCNF1IYCwwKyEJn2Jbz
M/ALFFkKVVdx/+nWIq4CaLeOJlTlaPbY+SsPe4rDRJ6t9Z8YLRyAUAKGsO2/0PvuL2AQJe0BR6OG
ywgUCOO6X6UnFDwTqNED9wBp1BuGpRhv19g76YzKFu6mxwYST9ZzciKSLZ7EdOPt+Qlt47MRuyAQ
S6YQMbRxsT2B+1pzITdy6xfRnnKyB1Vl0XsQbg5DOdEN18ecjg1QKYQwmxFtEyEoVmZsY8nLlMgd
GusGGNG1pr/MGV4fQRHVBQOew2zTTL2MbGtuvMRP0+e/DAlVK5zwaXId5QpE34mKU32/wSaZXzll
05B7fl8LEc/zQHUkMrE45jtzdWnJ3KmGur8SxLw1WPwt9DmkoVoW1515hW2AXRGX65Dmk0kE1WGD
W7gHqjl9NOczbk4sL8TZNmqd7XKbDRi0QTm7SmPxPJwe3c76hIWDVUkbH3txWi4I15Dnt40Fyohn
h/sd1EveVsW0Qm4jQvi16LA1Z0hdrVdOPu3QDt5DVEEZ+fuw2rwO3LORqy8mFXYEk6cLUtBW1RMk
yWYRoh/hvA/QqO+3R5cPCO3B8Xan4vYoTJCJvsa+iwQ9WWcuBFX4uhDCdUIcOWdyXsEEZJleU9Cy
kPjy5rEww4LvzW2P0lLWmPx1/l7CVQ8fcizkciVVKGVLoHfHRd3Y0IAHU1sZJRn6Ym9jzpNqrazb
2tR6MV1LonDIQVG7U7OSLDgiaFcsKYFiB9l5n1U+8ekU6KvTXsHwSKgwvuQ74hynvWQbmmKRB4ZR
Mlu8QKyq7nEpzpAAfZkxe3Gg8V9VLJF13Dec07D7msWvvUA7vZNG8U+P1sOkk2ZBjbW4Bjpa+kut
1w2wXPB7DFG9ld2gPkgoMUQItx2GqOnje85qm7fjNzsByLvimpD2cxZ+HndXQZc5jJUZYS3xL7qs
THHrR1ss57TP+d+MKM7RLxxbiIKl3tBo2tNNblVe7yuRTkQE/PiKltYwH2v144BphQdkkMaFpcmu
Z8ox4EagcK0VTQ8+XNW9BfhZZCU3L/EsBsoAVOFvY0xz3/6Uroo+UiXW2AJu+7LWE+g5yiYdxWhm
+dxIm+rusjAPbL2L9UpLh6mTAJwi5DINjiPnxdzDKatDzRr5uGAssOyBuGaANv94Tp/1Veg8aRUm
F5bX07DK/8/Es5UurtAo5EADzLVqx3Wmqwa/lYxxTlkxj/01F+WzYMToRt6vn9UMGMkz00xVGl8G
gcsTwWAxM9ZDdJM841VkNUFSjnKpoc34kTr3ebV8/Xnf64FNZ8lyAbWi8FaACOdUWOt96vnz+p7n
4AGP6ssPWf354dBj72ZjvVERGWyFb/dB1jsGgnD2f4iAi8AFHPC8BAqIoozkBqjNaF4wjZz8xR4A
93GiFQiTCxv0WrqBBeCBEv57hC/xR4Rgl4yvQfGVYpgTybkWgMhcB0MeOLhYqwUEo8tlhqWoCJkH
4mCD0tUdLxwz7zE/6zqlXM0cjpRQJzaSsXMINQaYDz64+4+dr7JO/ulqlABFOL6ALVAO45eK+i1q
uqc+0z9MuxJaARPsiigPHELwCz0bU6ZJyHaVh0aRw443+2w13g+Kutr7l2ivuc12IIP380Jxrjpt
gmwtI2r13Jd6qlmcn0ID4rO8Ceg81Jj5bZkuhrI7fyhqSXBuaU4nHIR9a3J+raSrp1PaBaPeBwFl
AZdmRLhc4QXKgXgTzTDs1Wj46Vns6mo8JAWt3M3hU0E2jPAUgALvNY5YUd5LTZR2nEW3bBu/LwSo
0UBcellGXMvJsrOsK3Rat35wn+MLaW9ChbyPjwaNuC5igeFsrnCbFqqOSlD7n+y/5xl5ozDupae6
l2+3iEv/dpcQQx6DQ/97xrG6JhRU0k5B5pnKBA7WXjH5MHzskQekLQdqVKbD7uLe8aJ48mCxssJF
GUIPWlekU35pGebXeaHldEX+N7w1y3Bcu9OKYtlhmBzMFzgAyOKjfmtsi8m9FraKMm2BRYw7AWVC
xWRHr/FoIE7iJXZzX2LHfXGUiseLJgWzRBI/pcgSLpGatojPa+f6iR8nwQneIeDq5lI7XFzQnG+d
EYdA3fNVdTXJ4aJlVs/CKCCdwj9Qrg/Z+eT/uUdn7urHjtam4OdTqY0k3kLOXTCI2TssOHnhzr+L
t6m5JsvHAUHsGEARC3WR2LHDar7Q+pGe39np2xM23Oj+jwkrqVcZshSY3NWOtsKEBnslfBenMbMZ
5zj+ZMPhMFRV4a+xFv6V6YYotzs1sKWKTyUcJbmGkOHWl5aUDuMJZr5uJPpKniLpAjdD5LQF7wru
zgNU9e6dgxAQ8c8l/7exB5GRbtCI3h7t2ACWYCfEkGmpbRTX8i3qk/JFkuitzfKGnge9085tESnn
jfIl/MBE3Z8jh57OWvB69eDTqAfoGkW32weeKjG1uv9RJlFppfPAQcEwtrPAS+SuCYIPKJVciaHL
CCMlH/G0efd9fPM4dJlKruIZWdiReB1HiFKmv8iN0cBSO3iXcoEsWOKUt+gt77TPfpa9LkX3XpZE
fLG3fWJ6G5SzmeSTKF7H1AbA2Lc2+gJJL1IKFIF1CLDrONGDzYU+JAaLpugAKClSuwVhXma9NoX8
DMSBbItSXB0BVIYK6k+gQ1QQ8sr8kWfKCLpXGFuCPsgD4UPJT+x8o9QhDHgvVnTM/czjq+BT7Ypj
g+n9p3V4u7bZ/FZq2AZQcoUEmet67eE4OitG/2qkI1dJRyQj4sVZWkcs4NpwwSgKvIN++na9K8ph
IVDdoRXSh2+Ih7a/C+5gMh4h2Qgns1TMbq35dLP07D4nw7Wnhm2WF4sDB2vD8kK4l5onjV1jEzir
Vf8V7geVH+l/tku5VRX4h7ewUNwcfi58QYVHzmgeg7OelyZibfv2ErmU+3t2DEgeqY6SPIPf6FGP
HfTx13ITlRklLq7cCGtgg0usWj7kln0apzGt1lTAaL//VU22tfP6lHXKXAKAPbwTg3sWQCg9aEhO
6tZnTG4qwvpYVZZXzBshro7Hy5RHy7iiDE+6p7DgdKiqU+GZ7Rq7Ht0h84d20r8BeboEXshONblP
NgucXGpb6Z3tX7F9CpTFbuEbA3cWYf1Q3pSqV4mt2fIxspBIfVhxwdLHbldrFx7f566RQyOdHBnG
A1F4nlfGuhcyNjoze1JnMapq0pYsAS/0NZt+YJEoEKlRF96pkGgNGY9+wRIoEbuoG60fOakGb1fN
tJd2PzO4BjZNDNjSnZCJBI5ZggQXwmYE5Dt5/kqI00PJKJlw4Rf7yWSpknUtKvFbb6YjqPIWzy4e
AcLKFZSHQo/IWG2H2pnhH/jBdeinKjOh5IKZxEecjZCTaTJPAQ7NYJdqcM9boRyJ+W5iJI50oTRH
u0nNRX+Q8It5QKw/dlP1eC2UQR2uqgI5J0zraZA3CuecmrP0ak9Iu2nTylpf4o1QAZ/0gkTcxjoY
K5BLWovMK1HuLB7pCz++6Nl0AzMnYjEmBaG01QxknevfuMHUNsf9uFFA4vn9ObHcuxrCw6c3yHMv
cinhoKh7lSQkZ9cQe5RAMTDf8vei2g5b3b0+vmIkul4t7AW8x7buLMBO+78plLusZbX81A54EbJ5
pliHF/kPuqmWDs9ljP6kE9H8LY18SExAYqxkF7E4DA7Ws8Vnx44ar2LGI4YbCw/MUytceyGwXJoK
EVITjH+xlrJgVxaMpm5kwgWyNWUKOW3RmfGVli+zby6HqAc+TlFvTNbUqZOYuNOUdpG25gYAr+yA
2qiereXwrO35vExBkL7MwxP9xtsfLIEVhTngD3sSrDSjxRP+IeilnZ8/lPk05cY94sz6CJLghpAx
zk7w4La48IaLlZAzJ7pFc8gMopRkrB5OoaxgaBdBDUkLy2epI4meAV7pWwECTwwvTuogeMOMQstX
TETWh0JV36YGWkQiisYgbOJ2PrBJlBdgQvJlvF/Rx5NDZQhOintbQ0WfnyjBrZQ0iD2ynj9Nj2Ew
iu7XobepJAVjbCEQ3ML3IsJNEbppRbHcFlKI8q/nu+8Odv8NSZjgIOFPwyKJ0I0f8BNbnI3lhd1N
bZmvFT9aIc2ak6eaaI6Q18O7bgxKohVXXkzmnO/67HYR1OZaWrExVH11+uZb9l8igewrQp6Xj0qF
EM84ASqSBKxxk5g+2PifRyViwtSDoYsWA/0jOOdInoTw+084DU12i57M6rseThyE+vUPJbO8xb6X
ce8ZYf4Z0xhPp3qOI4HGoea1n4YRmx6O1OV4ugemzetgriTkfxbge07N+3mDj91PJu83G/jvRnHd
q/jXO2CEs/ZOyghpEH4MEVcfJTJj8genr3RtRNX9ZjTJpMbJ6MblEXgnwhuDovCec3JF83LflRYQ
bNbRbswcNkJTKO0qHIw2kzXRR8xhIeNhK+I5Awa9EcYMnsA6yTQSVQTm5gz7HfCOi118L1FtFJU3
84RG5EsPVh8wwaS5HK6qoS/YnEeyTLp9TmLQa43D7xiNMRrz5aHP5ZXN9G9+IqNSFFeuem41lFBM
4KPSoP7H2t/EDgxOZ4ZKJ5y+FresQcIqSiAKr7ufoj6hbiEmMNvOqeKI5UN5bPlGPhHKiBKim6sh
GzEiE0A2cOBUpZg7Z167ui/Hz0KIhh2UfM8LKVrAxX9zLiEtMKXpGgtGmJWvE+UIu1oVo/RD6HKO
6jZqnL6iAFxHPbXEjpVo87+GtncutbJKQBoy4hQK/qSmAKevpfgK7URLP2TSo8OnUnpDGel5U4KL
nae5SqyMkV2yWnld5NC2cWr3X3pJE5QhY0LKoYa3oRXQDxCffhRULk5DNvHlX9iXs1G2kr49yo13
nndHtQH2F4GEdepvCgFHAgfwysJduDaHG68N5MlmT1zCX+nFvBpxEAhHkQPO/DiInPr9hGyFByxd
dRKyNpj1vi9wgKGJfen1mmtvxFb1QJpzSLSPTLbmDbr8fD8lSR1NcLHHmylriCkV+UdUNqNTHRrd
tZovQIGeFmvwMXONv01q6By8vB2ucGDNVfHZ6Csr+3yyMleG8TnWKmhudGUwcGosGiOYrxi4lEZD
OqkhgX4UMA1pPiFV+9BMO/d6KaVO71vuPtawfKqQY5gyHwAKO7NQag3HiHQP9OOan/m5gXLykHl2
eQvyIaDJEU6N3sYpe2O71TEJGO2sgVs2hHdAG7hVV9ifExi9YsHWH0Ssze+BNMCo3AZ4gTnYarIt
WNFsZlkGV9enAEeynLi5SMnqH+89ewRsfgtgHmLyrnfUBNtw6R/KJMX9rUsORV+nk6GM2IFf19b9
g40eZm3CRCFluPCdrZFHNKhG3EBkbf9+C0kZ2kb7VhCWdD1tsFm8SNj5G5/WqIt4rma5/1zSF6bW
wYuUdErc+MQgaJeg/G05QScfgtfZM/RlV09Jc4vFmQbtSp9MA7k8sROhq3gxZ5YDhC6KNal2r19o
vzuP9xK4cQxPtXBVulay1rYGAPjjLS/ccTqL0387CfjX8Eca2G0pQYwgfc7vWRlqQ4hkE69tedYe
63UYvzzd5eytnxnDzXKyWrrf/q216wnI+e8L8h52Lg9fqQE5zLE5vgTIeNJrrfW90yquPD3FHbdo
XvS5iP1ZjIWtzVkKKJFfk3JaG297PzbP3TFzmVtgf3FEuUHpcB3TSeL4tzPo5668t4fhXvMym8Cx
9GaI1vELPgsOo5pylAKMNAzXXdI0EIYo+vUY587DG74g0RWuy0lHTPM44yKb7uleVqayp3GCmi71
huF1XGtWuYUSzLWTMz7ejJXaKoXX7iY0KKch/b9sI4R5MeSBZSoVKeyc5AgQ2Zca/CVAAkHG0zZw
CGL8Zmt79t0OUUsrxerQ4JDWEQAsbEntjo7C4Io5/J9DiHctk+YpnQnmK81J6S7oZzqTMuGPEGVD
ig9Ye2W2D+yVwES98Cz5lN6o0vhlGtEgx5LYUEE4zcrL5elFExknhbNzB1YiB19h1Gny4tJHAH3D
zTLkOS9wVwd4xYore6XC7dRWoHAO1Q44h3CmoNZBiOjL8V1pSquoy+2Db4/y+/qKPP8I8BMC31pJ
177jjvvuVregvGAevLF5cfzr47zIIOLx/povr6XwQuhlf44cWyBoYbIY6vEdXpR13qw4BNc3wYtL
sL2xOynhOLWXVsfW0TbZCMOyEgl3XJeBF8ffrAqOdBhUFmC8R7i57pGDWxnmAwizZQnMtntwZom8
4oRAjBjWy04gg5+Y2u1BQz4ZnkObYyt/pz4ZnsgggAKhbNq0Y5UbkiCSSnCfLiMkP8CZDCv1b0JN
TgSgFEt4Ca+XBirxBqJlzxvXIZag/zIRrV3/AII6+m7GcqU2z282Tan5JRbs89X9xL2FRJ1J+2Zb
IlLtXzgMbY1Gc3GBIUb/pX1aTYPSua/RuzgwYMXqvQUqAwrJQnZ6VPRoNLAyfyOQwKpd8Udr10Nt
L6dkaeUx/a8AUO3ZTmiygg75C2vBmMuY8PNoxYOHr7OUOTQmrIIE3grCfUwVYyLjHr7leI2DhNGA
17ubSYBuTJYQptvaPuXKEegqVPnM/RuIEKL92aHUxVgNayRBq33ZuRD3A0Yr1qHpNr2uADcno6XY
CRuoiI+R283toVfh6ra/4bJQii0mNY88aroLtYhebB0oaNJQ1iAasNMx/T8l57ZFZksJpEO4Tq7Q
sysON6JH+UNZUdxk7+2AinSiOk7t9ZBwvKw8Yv4ydjrYCC4f+jklQJyXwCRBR1DDQpKXXTNRFzQQ
q/eqyRrZh3atnCuQ2acyUHDj14uHFLSuy5Jb59I3MQZEQdazBw7ATKVrJF3Mk0H4U50Vn1XakbXY
5G85w9cE+mHDlpHF3A8jkWJiWI0TANK5EhAAnV5E29uJ2dmh36cqqNyBtH7/sFW1mibtBLyuIh+F
2brEoj3DwhyDlhmYi/xaMYxr583uD5iXAfznb5BB6iVTgyjqaHkVoedYi5n6y3qobEr6VIURTY1G
Ok2KE0vVz+MsvkR8xTCWGDuRh308RL/yPqGzbqVT6mOmsmIYDmiBtTwYBD7mq6P+5UvV4geXR4F4
67q1xP5TFYKgMCNK4PSNDr7HEAEDe7axb6Z6K+EHrcSh9vpZ6uuBW+b+7hF2FOXuXQ+p+HrTxttI
HCdNP3L5YJ5laaKhFvFCBEDqhXdkPngCa/IdPbSp2OO8o6D+9ob9OBJXEaMg3/rZ1vJgax/RK6Wv
WviTJEuERXwfKU1N1vuVhxcSetS7SXKcwi/Exi7PApgPmHBx0JEI14GnFX6S5zOjdAtDVteAb/j+
XgQzsXxwFm3pkUcs4aoXdJbrMXmky5zIvrr10rXGO0LB8RkXMir3qQoIT7U4UFnRXWERB0M7IsWR
YH3zcRpcO2n7hPy/wYGxE7tWTdlOCLWnPG7lrV0gvjCl8gAU6xf+SfBTq2trz5KbalQju7yELiYY
vM+1aJeGYp1Z9nSCuegU5fbJrYgbSLvuPmDXAy8yavi0+K4BzkAIVF7XH+ieHb99R0bx7gEFtFcC
ywSllKW9tJryBLyWIHej0uTxQSLLAPjtkvlR4YMHRkUYeNCKw1hS5Nj0dG6XqcFn6dyJWD33YBIb
pjh+UwmkMdNgfOLWVoEbxWECdHCV9knmLPv7iXVTQe0K5E5koLL4ndjd3TEh3WetMAsiwxEZIUYw
lwUbY58/Xol3YjUzPz3bzdUKbTSKDoiOdaehG6Uh0nAYZFOVDDFp6+5JkFSb0AsXzcpbH1+WQa91
vpCdgiLKCfspI6pIVXxUv4unNXz03s1utdbBKO0hMe1wYHq3/KA9PD6U9GIcAIoHyb1Pqz/iMYqf
zgqetWVV7e6R8cF0PTSo11BBASxkcVeEi382KohiEWi3L4+Jz0bQe3fc1hYhQWDy7lX+NJz9Q34f
Awaz9Bq6YofQzXm+iZeNhTh2XE4bhJYtS96sMnrCxaBEHgdnQ5arhGNyMZtypoN/gayxQjfOZcAb
eMb0KB/9wsiRQMuQf7SPKMp8Z3lijd2MWhCRrMvsPwDlIjCCAFPFWWNeRXsWjtZRqy71HHuoV7Gx
uYm2mj6cWXdriwKzeJdSuHbxFCw9s6CPSnRuEKxcpXOSTusdneqPjjvy8tFpAVN5TlGFYLffE4jF
hhYzzO2IuAW4nWtfU2/ZqN0zn1dPGwwQdNoQFlZxVQKLU2+4Mxf74cTsBJZvqNkGMzTQjXho1y1o
ioryo0l/8qpJxDVLsjkNppA0Ta+7iKoYbLg3JkSgVUJRrRYa7IWMX/MD279NISEVosMMqII5VE7Y
/r96DK4xiaVIOuQQo9jusAlhhuXGnuS4MEc9D3FrTDMC3Uz96fQor4MgOVS3QpLM8LW5jEr714qD
ZKdUhCGJXRJO/7LjXpvMhU8uifEXTEiIIIcU+tyoOsxhVMlLzEZHbgKOpDhax3yPfy+/LTosC6Kl
33GdSLAGX63nvVVlSrTixVgyiyd6HEZ/2zN7BnGZHRkLnyiG295D62xWe5THQDMYG7n41Y8BHRrO
o4wiCbQvscqPsOdqNLDg37eCqXgB+o7YCAwVa8Jp/bCGUrgF4CdtmkLBdemkE42L+swLc2AFqWI1
98Aqm4Xg0Q7gCZ5vLwAFhOy6rYOlooSkGcCWrNVqTKeIMC80aXbX1GPAGg1QvvSdwIo7FfTiPQFK
jCBEw0GgUR6ODxbqYSWZwz3ANrupXZo1DZ5qbVfWdwjbeHV6NuvOAcn6XAxqY4lKZm8isc9eu+Ll
ouENzUbpGMd5KawCBJpVm0kIiiG+SaTJtp7G9JXYQmSTEuekKcVPFJIehfFSfIEeqfKrQUcK5SS3
VRzPqfQkSxvKZt0Id076bnX2RTR8rubu0Z/teiZ8zjefGzmFS2JgPr31mFsmv2Ke0eLK87niL+ZH
QtEtZgCJPCCaleG3fjXJTgww+ziTiaVX6MIm+LnxaT1nM/FtA6mSZHtmMbJd63n+l444P2ZCcP8U
uBKQ/4YuOrxOrKET9KeKNyeipPlyy/l6Im26FiSlZnjCdYdPq/584IlpQCiXkt6B2yq1FVl9P31P
4VupEcVgBLjsQz10ROKCJEzZQ2p0vdThYvyAHrruAkemWt+kuuUhnI3ERvP0cKxVRg0tJjMFFHc0
TmO67azr4NRN8qC7qYP/3MCLPwEdg4BYiChSWz1DZSf9cza/faG9kzW5ma4qq0v9RMc9KRLxgTsu
KZxuyVPym/rKwyH/DViVBTQzdhQ23/7TjJfxY3HFZFyQRSal/gHj+2hfBcYrLTcXJYw/0KlDt7wH
fiszD5x6wHa9PXqT47S1lO4VaBFXfdZd4LTsrj90qFVBPKxihf2gQCKQbPE0h6MYpDe4bzPuR1m2
F9ZJqSzRM583JgLIG7azC4wAcSmZeXb88MvLDnZtws2A9f23wsmn/rWL7BuAC4Z/qwEN0x2AEJOI
KmTzXKIf+kQi1JALcyjz9h3LGv9LZENLnQ4F6kM8M+k+W/V9IP98gAY45+wzzGNDLhNVXyY8H+J3
q6BoBFrK6y8mTFrPR+JzV7P7NtnieurUWYsHzmX1twXgXUdcYodXSu5eeiFPM2l1OhrXRbPGED/V
dyRbC/E4iKe8mVVoNtrwGlQdObHwukqAwJ7f8woyZ3Y5q86/NXE8vI+RZquWI4RROUU5Mfrd3847
yQiZFdD8KUHPno12ezREK+pMpKBZkPQTdQzS09avAfJTwiri3nJs06uyOJS3W2msYEWBuDYzjMdL
kzmeyhqlRZtpfi1yyTzWeyM0e+A1TkpY+fUZ+5KQn35JL/gioLeFuQVWiV+Ox5MXpMr1Bx+GgwnA
JM4PB9bYFGt+tqMzd3A4fgPsvj+BbAHAlbbncvKA4fndfWEkb2Q6SCsXDOI7S1oAgSTlXV1gTesi
PHKJkvgu8aGAcUjJdAJk7u6y8TCvSmfcm8pWJ+mzyVZWys8CiTxX8N6L5DFZaBMFT6VxWGTjEzV9
IhGpIU2GmBogSRBcprVWM1NRkgUzKW9aMBg/e5TWSQBT8ofL0X6U99X12EED+t+l2dn0KOjAIAFg
lscbV48YnLmclL5kDj2TZtTwFEFLpkqwiX+N8DxyWZkaB4gU1ANK3dC7U7FstoSPy85v1kdCqvp0
CtVGjfYE64zB1lq7RSNuijfpBDM9FWGIr4mYJL0mfOCxHYmCFL4DcoeHGy0+69SDAARPaFSOdRNn
R3Sg+vEEDOKcadjxXmQyEBH3f4WVYUgUew5k8p/SHYJkOe2jYvNpmJUgeqI4PWk7f5f+MZV7LQnI
2biifwhqk0j6vbnMoY7JvrgAstI7U4J1E7bbpcugj+xeG+vM8/9RA39r8aOwiOZeCqQhLeOYR/nu
Ft6qTUgijBhiuEGmaqescuuxXoORgk0NV+QgrwUfRX34zGW7IyPDyD3hkEaa6CGapYfgDBqmO3DN
DPJx2SX9P06OLk0WJQTnEQY74fUowOh9b9tS4EfmBxXhn5KfYjI/qpqVcfjkqnZxLLO+6nbZVXch
nycgnaBv1J1mdFKP3XZ/eSH0AT/y9Kg7eODcXvDxIBNWZxa/duBHFPFf2cdFo8+l+sQQBF6dqQS/
4VodHb1CeIe0sb7zooeq/f7tLe1RC7wjsQb3wGLN2kg3O1K63+F+OxpsA9Am/yTT+s9++XAM0LXD
GaKS/lM8yB1+lyBaR0CeGTqQd4Gvyr0fMUL9lxA3cPEcfY2fRRYJGv4lzH7C5h2PgPJMltbNhBLb
hbch91O2IoeYQea8HYaJWhm/DrcYMKoQwoHHPoOjQwLx4PUhZy+bNfYTUMLRghqRB0HBUNF9i43h
4g02BcajZqOM1Gb5i9fRWl8H8kv/jLxbhQ++LchZh+VwDxFfp6oc4AuaYGXAni9tWaROf2Yb5mr1
s6hXQ0noCCS9mn2HbDbmA3RbWZB1QZJ2ceLJJogWk1wzEEJlqhLRemjOnvBQTIEtXjuw9C8fNDdq
1E+2al3rGTngXfbdPBfsQqzrJTQwWZYO+tPqM7nlXFSE76ZMnjDnbatU7Kb90uelbuHh/KYWek8F
Yqa+8CT7Ru2CBrhTknJ6IBpeFakzwEviea0aMVHaH61CFlOh5IE9WI6SRheQP99m3DnLVkDUggmo
QQGPkYHooHPHd5YkahoqGoKbEakJTOqI+dfI4tNuFZeHH8evvR+9A3S6Jv262/cwA0BbSwu9t12b
0JBvmSzeIXLdvCU/phsxczZ44o7CG1YVyinp3ifnsEfz0h8JQibRbYrsv1qWCtshxWjY481tV0n8
b+/+SZ/Da3J0uiq9Un57YpH9wlQl8hw2BIx+Axm+sKPJSg+uUDDTiSbiYB7t8xIiHMYpKrrV87JL
nAQBQNhK8BiioDEm/6K5y59CgSO2BhVis2Ecm7hDGws26waqBuDXdFFCRoQfQS6pBab+D1DHfNJb
imUp9Fz2I16ih4OoEvc6Q/79JTjhyJirTvDtnZcn7bUBS3VIzu/wqJGhMdNBJs1bmqU8WqOCa0DH
97Lf1eCrgWAGwha3h69OidPAi2aod5YCQos0vcJ3avSkQVOi+q2C8m4i3YHiNw4xg2hNL/Hiqsso
KBk9XTVdhNh6cj0pK2ny0DU4o3G9Tc5t/3guTzKcwhzrLztJdkSAWWu0xSfvkbUUs014rq977l9h
sbpLOm5VLVgaZZMKrfK7irCWJPtFrU6VL/btC2UykTLs/dN2279ydlicOeTy7ItlaDqte3uCJFwl
eb/NUgLNtfqyK1I8cCk0XYFNGCKiGLgttkLmWaNGdqDGZtbiUXcE69AD3IKaL25ubVM00gfn9h8+
xFzMWefCcFGTKTJZLxiYt2K6x337mEp0RYdcDrfuNsVR3+ROHWKnQhTQM0OmlGhWajOovZsO6bI6
AZfyAY5UnaqgvpiufSJZ4WXE8GZL7TYSVPMXBjtRkl52VnnMUCyPk6FrVBbwSjUNToVvb6/ja2UZ
pDRWPcueR4s+gXkF1yE/Cyfy6spnCfaZWUTiM0IREEkq3uNX/9W4v/eff/6M/N5Oj86QqJKbxnsy
PHUKuaTw9Fm4LQubT560RoH/eicDeWXp+kqsWxsw/Nsxy9xd8U9xuuzzgTSYje5t9JI4lBlZHvBr
A9HA9P9vwyCxlJoN/+jrh6Gl9SXx3j+gnw4g3Y6vqiPiriZlpx4bom8rVt681/OX4qxmZCxsZcgX
b/PtnkOT1a7lZX9mF3Pi26P0heySS+n2HAARw1HSAni4jUj7d5rURaivTY5NSZk5NeIM+76EknB8
XI/4nmoaLPHU3reMVga7WUYazr0/dMn9waq0poJtpY/Mty3l8N8lTfe4Pj9ZPGUbJuOEJGmCJ79b
Y8VvCFW8JKC6NP04ZV0SdGWedarMcjRlL/kAxLsi3uIj0hLHuFjtpPx8BwH8+Rp2zwrVHdV1JbC6
qJV9lDlO/vWH6S8dtlF7Vox9dsSnZvFWKArin4SH0VySYcKMgXdU0WhV/cGefmwRrmeJROl9E1Yz
+EtZwCyH5P4iNcHfofyyw/WTcZE7rwwFPNfYAN1f6T3UzalMVORRAO3/6FtqJCQeXbbB2bXZyLZ3
Ak2n/2k5AEwlLIYlWlpoSncORC85qnetlHG0NYHEnRmBbRHqr7YbGBi+q9cdcWQjJnnYtTeGRbs2
0Lbg/0NbXx0T5q/xIPEvbt1rJacJiAKZr+LgdCy0cJF8U4G1X2iMVf3TcfHBgFbm07RwTcqtmW6C
X5uyZ2Ptc61yDZUOcHuOp4O5i2Hia91RNdIcKb4o0h8Rg+tgVnaB0iECJgwvUSTV+BcOOsrMwDng
bYp4t0CEB9k6g8m/Vg9PbyHsbVAn+FnD27HtoE2xsGzZxaMuv451j8tbemO4sA2yEfHkb8MoGIzK
DvFMvXSjsssqSPmQuo/QxwOl7/XnzwUuvwkn1F0WdYOgXP6YVWT1dRYNNtvx5gghFEuXqNArX/nJ
NRJv/WvELaZFipP6/j5+YvdCWTq+qu3K3WFss82HaIB0PgOSiPvy3vd5dJcqco3NNNQ1/RaNN8ji
xtvzu2hSfMdzRdY+61TMF214JjhIhPNgkzFP+dwWQUc2DJtH9OFgzVSS/j+pTkiYHeGGJkkFeBA/
fFpmkNCl5GvsRftZvOtZ+sBksowgv9w+76qOkkbhLAMPwYkAJMmqzM1xdDgJ1Ql0PcfAVQTbfDHn
njlKzd1t9l0GpZx25vWs5qQrk2OwxviJxzmRXFHi+WzVCUYUPF4WyrOCrIR4UzusOSH8SwLGYL1I
KjUV+LdVEmhUpulcI/GRm+io7jPGeUKNXThCbrpKzi454lMNeLgAxyZ3ANvfC6yrUfF6MZMe0L0F
FCP+n+9hmM1vhqERoNkWYKbh3cRdLG53CInGd2Oc+wuXucylbs+1TddbXGmsa+maP81V0QpTkDG/
O/KxpqHOkgNlEcWcqKeqHQorCg/uZ1WU0pCkyHcnyaow4LBJ2/DwwsRYdNYsC7ob5DSxhaonnTmR
U9aHG7IuzQIRqG7iQq/73AcVxIFBzGtNeUqEEhXXdkL+WQM1cSkVrDFEKBhWRPPZtaUEEe68QzMl
m8UFn8oqxusufIzCGfwWSyEWPzDYcfT2t4xDyMKY+DN9eAD/9bITcqrdUeXUqY8BNqZgwNX7AqDl
BYwcWR+WlvJOEGREUyOXBTY0x+VsSUZTZdwq3AM4/dd5Ug1OLrAmbvvA/ui8unJ4KIlJf+AKbDSj
NWVFGjPzFQ9NMjHu1DjJkIeXVNrUVMZGPaFHFOFONKkLC8ouh0q0vWeUHvTL0WWYqY4GWe03a569
taf/H9d3TKEa7GjgrHQ+MNvP16pZ657wlgBGCr2YagXS5dqBYEITsCm1uQ8Hsq8XEdherv1BUCwt
3816KD2d+6s1zDEe2Vhf40eoewz86UZf9WtKlE2TCKfNbOyRvdVZlop2+tU1Y4KjcoCLodEaz4v+
S8XYNi1Bo190CCTThn+A8/VliyMDOeNiHaS9FMpviFvr5cNuYyEtg+/HyVsuK5ycwyU/uHrCXAkR
G9Lx+NmSgLEz850XxQDTeI2aApFqEeUn1qGGrO58YLMHxXCxOgLhehQgtCSgML4D0iocEH/S7IwR
qBZOczjFQwgz999BY+p5Kmof7k+YK1gqS43bL7O58F3a8kLmyUEHMp+tMhaN4JMJgGbH+AmIhc38
eHJoPnI7PYpX0LNW5Mz6eUc0+VM+EY0YDwW2m4KPSmC6EjtAQuCox3F5ozB4bNLlwIJiKVOoa32W
+TGEfefLnHt9fWtrcQOYYSJFY4w3fwbxxT+r25+WmIjo+KjpvIulyz0S3OB3g1gNOg2J3ZPGwvxd
/pSqjRPwagdY18VvcoaJ/1fXfjqgLlhVca/eOq8YW8oUMJILC2RIJ8aWHcSCMBO4e7kHhY80kP6N
t0MkU48rK/jouRUI2QzTgrznmnEB5JMGXAiLlSNeFMvxUEZQDHdHb5j3AblEpCW3c8C58FOLfpl4
JXCKCEc/D87kgraR/gF2lmL2B9e7x955//uJhuxr2+Ttq0b/PLXys3fXImlmmX1bPg9tgvVjQkxl
qOWFZeagZdHAWlYg+CRyAfHOYWYtziU/rNYdC48mefvDWZuBRKCQSJnR5YLN7KWI4sP6uRy1BS6w
AqDfakz/JggZjG5Ry/JzCptTI0/ZBQohucA1Ei87lxG25CqEnSewSCb73lLhWZA62JqeIiobnlYB
f/tStvuYG2Ln6a6aLhSwgIW2AFOeLNmgxZ7orAUlMik2DEG29H2FrvDNMwNQA8YbUpJiuX9hhTi7
MF98Vu/cP6fSXNvVKpZBK3IXHjVuY+Hdwf1NQHhaIDWKexTDUiye7mi4pPWJmfTJDcmJM+K6alF7
SYn+n7cvxj398v6j+BVxxjMd34btKw3uq8KHixXMHIcgi/jVa9CVavz7kAQ73MXwajLFGJz0WJS3
okoDIsPHSjZ0zkCg8KxOx8d3m7+Yv+7mKpjvsXzAjb0PZTF2fKjvBtr0SlNRBh5OHdu6X7hkvf78
dLm+4wbne9Z2bNzAPXz+yyWHc7CUvMWmXAoE0pdYZbepdWrGxJsWGne8H03+GbbGih6lVOoyIORB
Cmvw9JDoan90h0K7II9MvVxaOOnzi6tWZYBn2FdD1zwnT+VfO3XnoYrY2zPQwhvEdAzF8b9MuRoX
VjfMRmzvBJ913PqTDdR2+G0KpUkrf8i92q3DbJjactoshdefv57wRCIJex1GkvJaEsUAew3gaAua
RWUZgc5BgrZD5aWugX6PdgQ4Ccmxe907cu+SDizubSN4A1us0DB1vliA/RX8IfzqS/ivxpk/t5gu
vphnPUIw/om70ai65Whzqu7LZ+lU7OXQAH1MEGTii44dnTRhX00ivVsmk+a89x9TYi2RChvwr6r2
kVgP77Y3Jr/wlGa+3RCvOt7UUlBvu0BKfJKsb5v1x0oGhv3QbxKosyfz52bJRpKGkA1B0bH6s/6U
LYYrHWrHJXh+vzU//UBHbt5aaTz5J4YAGvbr2Hja6eWmyktr18tN1XfbFOaFAZlfOU906yl0nLZ+
JrElL5s7GYgbHcyTp94aXVzNNNwDZ3ccEldrVs1cP11GaUJIfTsREiOjNE5YEY2VV2TVtm939Qt2
CBSpRqt/PURf3iEI3Bg2vZv4g5fzfqLJZ7kyujjFvfFv7SBQ0rHNuFcrMsOX6+I7aQaz59Btv53l
I7o6HjGuQRcE5570UXn7uzB3nmSTz9RAj5Ua1WX25G5NhDHanxRAwy2/weq1rd8MjLalLxF5/rVM
sCAdbIzlS1gUY6xBNverk+eANYbkoFPfIyhid4LvAq4RigMTQx7nJmrg5/7buZo6WEJoMmQp+3pi
12uhjsnWx9orT4S2IpM83aX1er0Uo5bxl60hSHpLgSWQln+oAZiThWdsWWdl/mhlv8NsHouQVf/Y
ajo0ZMIeghJe+//Z7Ez9IPZd8H6nTALED1y0ngZRMeyd+e8nYdEnkF0WpWuKEQ9GM7l6bM9TAxGy
cjvRuzsUDNf7bi/uu/PxUQrSnZxyPJuU3VsO3KS2ove+166qiy7s57JaRK0YJk0cZtEe2nRf6H/J
tj4MFIqgVNC5awIoYUnxTJfxzbsLqh3st6hXgsm1/6+Usvu/Kk21a/NqNkxTGTehNSPXxmTrrxEW
Zx/+tywEWDYuK/jWIyYIDqbsiiwLjjeqW2HKSqIHT5+ktvrkjdKvJHbkheSeAqUsv+oYugyxBf0h
PARp5Ea1nDYnkEtuDetv+D/kUF8QpiYnxyYYmU2pDcFFhZrqh8up1okjD5Tw/MPPuyNxBU5Z2e/K
oQjCzTANrpVU71yugzYdoWCfN+pWmFzsH3vtD6V4iwE2EHYjChf+QiiMNAVF+6WOeYWc++v404/G
K4ea8MFRJj2PYYWwGzdKmER1DexzwL/3HFy6pU9B5CSMas0HmPZPobJ7qszRsw+lTfnIhysuRMfO
OTk31f+TFnSthwfusi9wUpp9wgURabGTwUwgyknl6+b0FeDzmvPB7Ik0wQQYAEpj+MBXTyoG5/RD
6+yV4WqWaMNba4O0osMzoN+ZW0/tlYa5EXZwYwWQH7tQBXXPTeF+U7uVyQYVfvYBMnAByJCrRQRb
WskckoyWuimwgUhUyqTEVJwzWsv5MXC5w5t7P5V8p9EZ/maxy60h74A1IPhauch74psH0kki2jSn
OqCKJlRcVy1xiPfse89czwhZ9J7kEQkIfFSLERh6x+acLeGB+E0OGhwznBk7fPcVOubskrWCq3JR
A+33LQpjw8T2/wPyDO6IaqZpYeM1Kqf4RC79vE6tKhakDDqoHNwiE1v4/sgyIJgsd4batJVJbPqT
IjVxfcYEflb4Ufb++Hv6dqlAynLUrkFKYqnnd07x6unR9+CUtrqlOAs2Bm6DB9nSRLmDciKPGoFt
UgNcUg2DtAlvAirOFQAfjJkuUirs5yLjKJQA9NirM2r7vGrWNPQRJ6IpdMV7eMVy4IJAQZ2Le6F2
59mGzjgIMZM6bdyMEX14I63M9ZvHMhIcV9q3vkfot2+zoIhPwN6H9u63gIhMdf4pFJJCnFknz38Y
8ndyK2+K+xygl9iH4+YX76piXkJDUg1WXx9HEhivkeUl1sglItog8T7GJZoxt8VvTzaY5eXQsO6K
Gp9eLOWBxN3PSl5D28ahV+FwSpZnEg5qOPLulFdRfyvroTofTNWrhDFP7uCUJF6vzTBSxhNvVnsV
Ru1/ieQaV9EIrl+nGfBKavWbga63Z09+lE6AItQ3du3PuDH90IitToD9HGLzMxz22DET6y2PbmYp
bSY1gf9fvo2gqv6FkOdQm3VjcUBpv3lJ8OByvJKk78MuKfA4Hqw2oRjY/JLOssF2vZwJCwPgazAf
6FtNBqLnFkiLeDImqWi5kTDTHSOiN9QvmQBVwnPcMeKF7yMnADL24FwuOkqGb6B7ERuEgxhnVjZ4
HzNARUJ8HrzccFM9EeEm3eBzPb/m1NRX/ECSv3GwolTqGcrc+irgOzrMa8o8GvyOZNsvtX9KpXYO
jUAOqmHHMZwzAAoWEATuoeSvWpJC7nwA4dP1av4cLhsBayp2RUB1uFX9bVm/UF6ksXgDybagPCJa
Nwt5tnQg1k5hybLwIsct3ZtPITEBgm5PkNJ4tM/hqwNrMvK6BVRWOfcELebPTysm2U29F8Uu3qFE
yVWy+VZi0au4M2x4vfg2szCxEGRcCULg1SKTHxrx1Z3VFn7xS4BHkfMtYNE7FOPaE0+U53r5hWLy
mmr3K9/nlkU5wNodxZDKjdVR8ADqv/NTWgK6FE4d8MdkA983jEbV9OCnYk6I+vUW/YQzjDJNUeu6
JxSHfOxA5JnHvIwSVmNI6n9LxFmE3O8zBB/hGLJMZqKG10UtKvVmN/f6Wp4SOWvsHe/xn9Mp3tIy
niw3JmkGf/IoQ650K7duh5nM7oirI+F7gAHGVoyhVNcbzwxkwl+96XS76BrBNe0jAY3SuVJJHdzp
8BaCMOpcXLF+SjYACpvg8XA1Mz36FqNIuoy9Z8uYdHM9iXG3BXLJsej+Lue9LiIWFYwK3h7jKouA
uMngPRdLwgclHK9a8/moTYXEkduXJZRakhm2/EuhyrPnXpZ4lTVSu/wCyRtnkqrnmA2c0xa+GZVn
cPUk4bwBAmJM+ynb9xejbHRTLGRqT5M+PysvFOWd/he89Foa8grZzklgtTAzL9ndDLFEXlY2dsFO
7uLhQdCGnzc0E2GXGxJyUnt1/9NTRBfN5V0U/ZXhN9pqR0XSFiMBH7dnqM+ABJ2jQeHbFOoVXLBY
r2dyruf99ZSsF0DmGcDjTT8YC6Q9rSyPJ4pzSohXFssTyJedE7zYNONMSVzxDE1KbV5ikERARcIw
QAtyPyOQ/sMnXq2nRgH1hlUSGFtemWknr7tPhdqkvDHToQyE7J7X5JfCztCQuiE8UrhHbwCDfsDF
Lj3H0cn/8aWL7TmCQhHPz/8aaezx3EzBcDiqPdkQCWs4r4tEeTVBovFqbKuztXo3VDx3RfIDI6WC
9qvN2JUcq1zkqFkDPx5nvqbONdjPynRACDxZOgsPpVSeJHuzOiLhN9VlwW0Qmq7uU+qKy1NniQxF
0Xy9UP92D6poHi/4nbyNNbmeM6vuEQ4WSeA1TpibuUY2vsp4tMZl96tNkt05BWU3exoW/tXd69Um
PNbNYU7wDImsE3+35H0k0sWSjSTKnwhGwVc6PAmRhSlg8wazhB5xD1Z1IJKiKfEjMvU+Oq27yjdH
SokZprxY0KoOf0pimoopXv8T0q19PKl23WfGJgV4zkFsmUy9x3L5o0vFmt2A5eeB8/CxW0jHcUxF
9fe0TKmaHKmNds93YgGU2B4qkmUYbLkf+b4PWTKK3qGif5vcQvSs/xsXN1aDCYccd0jYEvxFS4oo
wU8Ssv6s4oGkcj71SY1CEVG+PQV24LKhYgC1kJSX3WQPvK+ZBSJ9NaQvl9i9pGGTaMy+D2vM9vYY
i/XvThTK7IiDZErXItR2MoUxkLFbCo7S92qZi0jDR9k10SZWu7hcnjFjAr5GtILLIeMdZzdqwpyw
NX29W8bmfSKcJNs1OmwaALV1HCUo2pEgj4tdR8K6r07zUbi/Ort/MpT5fEp1hBZWc13Ls/xHcOxo
i3cq8ErmU2460EUZudgmkS/nD97+lEV0lbHtEmZPvvm930mtBkqVonJ6+4/eibnkjzhyOqg8k3bH
FVaQV8MljH2Zt2D+Hf3KIpMKcnRntKx5nZFFHVIV+nxj+FhNNp0kHTCscjXYdiyiNbw0nna7MyGV
Q0LGHNXe0qSt8mCKdL+QFJcnorpVhXm28ILzxmVHLs+7BQROS60VLwKHTs8Qmv5AfMeL1jt4w6/y
+/7BiKG9gtl0TnrZgjm9ZMJkXRwCms9C1Usd8kE5NIagWFk1dX5x6j8HTjp8TWQpXQTpXAoojUJQ
5PFb4bez0+5Q7zUV2jNFSLzQSl7kFcYyO4f2yjHiQcGN6B1HkD8WmgATUl0uDMYCEO7dAe4uDGg5
kvl54E5uhYh5tdzB58aVz87Q0NGOM0yEia1feEtSulX6L8aUVhForIggVuroDpnHjl+F/Zzxq9Bj
H7j/OVJZM0ittOPSs6gmz5mxMmDUG+RECn/cuxoKCKcIgons6uRD63xdBYHHzzvfsczAwZxUd4bF
eDSNrIP9QZakV7M6puowndYm9wpt3Bcv17XD7NL4H/N+MiGq7q0DY2LSdjIt2nm5jpbyQ6Rx/YSV
kFoN4Q5gmuJ1LODzMCAO93etlr/Ufq+daoBM5d0UktbRVYzF4GIsRS2NNUwHE6zH886zA0KIXi9s
/pHfyF4rL6IjYUYjCO8SzSr4Jgdb23peEQ31q6jgKkR8oYrZaZzgQN48GoJjfopEInrkmIo97eyO
qan2L7ORIuulE75ZdyV3CwzjfmPNFMgYHQofBSW0iX2eXZr06tziSJxQAx3j9HUNXwuKSrwyOhjo
I+1X/vveASNu185ODcybbaGZOPLFQ8NuTYZutfGgvLkq6HrOouZJtgkdTERXcF2Jury6HJvg1QHJ
lOVq2YeZbGuBeue6fyct+uxizAVGIDpMyiqyAfdRjA8+A2ghHEr68A+QCMVvvSmi9Tv/3EIdJtcI
fArCE1jJ0aTcEHB6hEOEgYZxmaT95Cjn84J0mIqJ+Ele9B6vZxp5DNyhn+oqOiTm+c9plSKcbvQr
1AQ94BIXNnk288rjDWrkdcSyubdgABOz87HuNaB85nllU8qAkvPyoJm5oW4WKa2E6qGo1JS6rzui
FmZicZlJnBL7NIt9LuHORtmFAwW6JsZMmRPVqEVZJuEc76atNw+1xCbXjr2dGwjjmYvl3a9QLu6j
N3URenT1xA2elGhX23QY2jIp9HrNhlvPInaT7TnUudWs7CafWo06R11MUonH63eoNvW9uSv0lXll
hIcGPJDc17+vifelYLkhCckGXESzMEfq2MYG8rp1ANNfdRmmVrDv6M/4YdsuM73JwSSgn6qx+BnM
7h7vabxjhuYMmP7PNBb2775lTgWMMdMrkR4VhJiwfC2HrLRofIGODiqxELxVgj/9CKDthfNMW/KC
6CRfCdZOXnkumrTp2S27N0C8x/CC755Hc0Ow7H/iW6ehLWOG16/1ymSQYLzpLhLsb/iHqayAftPD
Oiaq1DUcKTS3pGKN6YcsQL3AnlTgg3EO9L6VAz6u1bMqhM7IEO38gDNrqBfK52xNRcf1+fqjO2Vw
9zB+65c1jnWcUY16H8q+GzpLTCyJD1gULKMg13XsGR4hLwtYR2n1VQN8BWjhfAiM8mv4Ll+jSa5K
jKkS0q6AFsgHpBmXvLV0RuE2r0EAUm8tJ/KhfeVWIdo2kxtBsZgze/hThOwK40e3FEiYi+mkFplp
zSfIKprTQs+Ae9jYkJTkgF2suWToTOFtl9rkHPATxT5uUMRJkO5JFo1FczLc6hrAjkZq2bZeh1oM
n1q4Mk90X5b2J1rT0t1o2+xBWuOeoHIDFC/XcTPLxo+d3y5V7LDyPSZY/yzUD9zYwwzCDRAGwFyv
4Tyr+GvubE28mO9SHJmKoJW1ng7fARnF7e9NJBE8p87+v2kao44b4lgvWs/U9X5lwzZa78RsjkHK
/0Qrm+EkOmeUiqMH0E2MGY9Q79LSsQFG1U1ZP5X2feJLFZMQvaDNuodDSggCQPNb7vUczWcehv82
hoqa6DVAsJ4q4MgVGqOUqx+W008oWFkcm/wzp8f3LfJdlrSjauhB0Ny5J5jgkVBIt2zRfAmzQUi2
jzMTJniv/wcPDESgEy1u2dqGF7/sFto6jGuhArz8/otv64LOzgacuce08lj9nMKd69vEZGSnxUIN
wLucWg+fIWm1FNcC2b4y9tnbnH+fIs3gse+jLNs1Tn+NIqi8crloT8SYRFttapI56lr/2GLGb/WS
7iOVo31v02wCajBHqKho0yvdeqRaKO3Me3bjzA8OhlkjJ+XmHUBlv+oUsdCNC7dKvI2p56x7I3C8
AhjY0AJiUr4+rUzaW/7//ZWWwlP6ow6BvwrkwV+OR7WxJLmL/+nHN2AZonwYTiRIjqz0w4ex13G+
YPNVGYxlhX3XSAd14LBHXV7XCm7xxy3IARX8OaIUojLaVgYvbcMpaVbAnaL0FomwywHLO0mMMOzB
U7ZnN8A3vJ2Now2dVjTcB23fwSFOTkQgdi4ZkAoxMbrI/qsXBptF7GXXQ+pXuqcc7w10P0ijmRsE
sfVqD9Uxl/kFjVP9eZbzcplOXOvobzBXZtVF22Xbhkw4OpaMCwRrIcg6jn7ZcBG4KN1MPW8G00aD
ozHXUXlx3/A4gpx8PzYDlSIOECjosf1KLKJQZ3nCwZ4nhkquWYBQLufABS3ghj+dZZqmC5yXM+/3
n9etLyTVa0K1emJk6Dqk/SPahzHKGM3tzq2A98y0EvvpswmPl7kDOOnX5j6rQhF9G9lxvz2MOdaO
DRyMvJUf2iMByzHWYWiCb/ioSLSNHuifnTsZWTW7tOv8cKkfuGgrzGzKX/3ehHaN3PFFemEzpJpF
nahvJw50YZu6kDr6vXm9iHWqAYF8M5CYyGoPLJEnrChCECC/Hndd83HXrBpb61cMKNMnVpSer+22
/kjLdzb4OFKQqv9Yal5hwQEY2F9Us7CAmA1wIzEwL+UOQsfvViM3S/3QT8Sv0GXY6D8s31rAhaG2
g59zorVusYhey3nUZHSJqB9rXYry3Ju7chxOmLny+EXxnhpvbyOBnbYmYShHwU4Cjcp1jDvMMiS0
97oDrmtIkf4sS5ke+kg7GCARpEGndAv6Qbb+z4/kL8QL8IeX83/ykvj/QcrfJkQtAQ7ytKGm/QLI
gizvgNMYhhEumnUxTYACEjFoW8mByMm+i21ECI8cfu7CmElocbMheYvZxz7GlDK10SwF3bkWYWWp
AaqrGnQwT4N5p4okZ1bhj/Qrl5YAHeBQry5KVaqC4JBEgMgamiUWg+lEhWI+VDRI4n9MoozIyBAW
VEokN1K5sldH0mLRj11ayhft1pCYNvUo5iEA54dEg2DL20samrcsNNmUu38EvHHbrf03VnWs+xdQ
pYqUXO34X8ifiLMbwyhTMIivPerfsqaSLaeveZuHf2JGTGI1SVYKTULxMxOruyw9mN8IsbTvZkRX
E4272iVm6PcVzoOBVWmJUh5lv5FSEBWreOcx86GK49loY3HP4A2B7CbM4bFKHe175sE/FceYZR0G
aU6iqYFoQNIcmV+JH9VkI95KvDpHjb43SVGoG7ANqoOavDG3g1jjmB6hFtTkCDt4e3sqqakZeHLx
m74uE1IyGcQ79YOZ/M5uKZYR8gVFmzZd7WTkoRIbYADBfvW5bW4hrG49tBEEgzRvKta+sGnM2k45
nrUzfjXXyVH3SrbgDVt8OhK61XlcL07J/CvAE1mEk9m02MA0c76t0kIDLx4MZDIMYfKxjWegYVfR
p1WlbgjV3BTJYBuG8ujdarzkCrQ6W+ju3n68v5YR2FhwAyG8jJd1doMhsTGXkSFeIqKDqujPDqDN
HXf6guXvTT50X06LK8X4xZIGHQ2Tg4jkaX/Nqe8YbSUCmTYMGlYVhIEPsRL2JjMw+59Kc2xzcy16
V8DLYa/VPiiG8kcpet1VhMjkyoKQkA1nyGHTHzL9mlG5oWpIyb3iTHoI6AW8iS5kWEx2+ZGmHwF5
EF1NdIDOFR7d1dlESxJklXG7aADu5ESb4gRoUOXcGMlgO1rBu+vlD+rcrI58D3Ro3LJ3iDhQy+qj
a4J/gJtS+Xaf0/JORTD4mV7q5YzZUYvxj9SzARnRNprX4wG5C3HvfL6bA1rA5V0VikqSlwy7svSs
PstinHlZSJJZFNo+ildM/LY7JvtqxPCed4nTVhPegwMXXhWdMTY5y9mh2Um/J90u/T/j2aYJa+v1
uREUqB9O85RaAhGgA2nXr4D7wIhiPStcFoHn/LAPHTpMNDqEg+nfkHndtPyju2J0Ch6lhvLLL21b
O+2HIs4Q90kGKXqrxUyDVxZCwyBoeOlmjslnEtdHMVDs7CsTh7NYnQP+L9HhrZNbaK0cMf1ujByU
g/Z4Wij0TiU+jypKS9InRq/qbaPcQSwp0OrSuZl/3CisDWAcQlsXTVIKGiWPUgTj5vdit0dhPTQW
zKct0QWBqHnOIzN6X5bykbLGo5qQHkLjihaObj5Vc0eQOBtn+GnPLiLbhM8Aa7ORtYoYMR0MVrTi
idWP+ZD/QjvFEJdTMHlwHrUiI87u2lZ55zFpwd+t0sHwmpPWrdrjVWDqYoYau9BjM/exDyH10hmC
pHWZFSftFWqOWUoYeMZBAD1B7cQ8iT7FgUueXfmzD30A+y7Ag4AXS6X1WCyrF+dcnLqxOH4cwRWC
mc8FRtMhp/cIqwIZ0R6WHmKurRAEf7qCOhjRB07yBzlyQl02Nj8tqRQ/YXLg+OKL4ej7v1iZ4mCT
tu1cZtV2nJ534No4zW2sDJ8MApkVhl+gOhA/SSdVjTGWSe9NJdT4larzsWKpg/9CYu+cKkVqD4tM
b+cV1UwjauTWA1HXRF8vj4UyNPg8RSQxe4tO/ro6boRZRfBKCoA+7tQLOfRdFwck4qaEZA0TU3Lj
fMpLs66uofG0OVuorp+q/6Um3sOwMfL+B7ytfu2w19PrNR5LcBxr9uvwAYT/6SQGm1uzwYvgz5A0
il9Ip+o39hV5/Edhuh2lIsHHKP0He01rH7qbUu724LSgeUZkXSpRNnNeZKfllrFReWCmNB8au4Yt
EPvjgy6PP540W1TDWlnoJkMCbcdr425UnPgU2C1yrvK3IHbB5DPV23e8tX6s1/oe2jmADXd1yT6j
TNUHoKvL1ARyvlgl6h2gA3/t5vNk36xCajjvilaDzE9mAxwGjnvk7LU6akacNymJtRN19tGtdNcP
UsvooMiNNWYd9N8Ua5iYaPB9Dzb9rZ16wQAl7x1MsfZQKcUvc6nyq8/Y8Hg6XCiq/u/rNESyGXXn
lYUM3er+bxNqcdaLIGDmCdPKHvvD7TO6j3mt4AEGBATGJpg4hBVB7NOWRXw894IXEWpHyfITsXU8
w40GVOWc1z4iX3rN4GLR7CPeJD7mep/7DwN1gt/c+DHv7Stx9LWMN/GU8MGX7d1iF/wDNgfLHtIP
N7fchoJyy9wjgIuy06eqWSfYAEfPkJ0OEFx2WDvmGym5IX8OmeSBe2kub/Qgf3fiWrf9mrOilIOa
e5skgwj/3GFAATjvvaDp+v/zusn8dQrJoaNOYJIl1+JFsSfrRQdkDV2PZhHu3JzKggyz5g1quV3J
obqyfvxX0gbUyTcQXOYVkZJUaDS0fnPVzszfMT+TzJGCOyvUSbRFtsMvqNWybiK1AE+mziOkE+iE
7XrWgi0gPDQLcFjlwNNYpW5nq7NRT6476SKw5YUWEwzw+EzHFln3/KJUR9+kbEvOtL5sArrx9J4F
r9xqHqMpo4hzuk3zYy9rVvk46FpRv0eDJ/s5rpDlGPGNVRHIUtZMhDW/4BxVmhsalVs/Vg3Xh74m
13/NoYCSGF2fhf/H+M9tlBCW9xnjmTknea1OKTMRU0dHpYJsF2ZTVpxTav5i+XbIz+39wnRZLlSn
ZP8689LtThy7hTMN/oUud5nczlYjnU+lvQ+DpF8H/sO0IFLrPqy2SpuL0/0urBrkXKdZIPaU39bl
TKVP3g1Ck6xil7Mu2Ni/XAeup4XOoxsfe1f8V4nwQ2/cY90UNMOLiloTl6iQc46SFfmG3ob6N9u/
baSBW0I1RiCKTgRrel0D7WfJbaIyp4i4vNaQSuvJYYM7lFwFYLcvkNYrtGVKjsgj+XEGN9SZ6fIN
/PEARCHaRv8zoC+ZMCeo0WMjvGRiWlqCaSmUPqRuhs5Yq/pD6bN9sGeORo5pLg/gEV18IywcqgDc
BKHA8zob1Ad5scqBTI4C4PXk6oz9ugi7bQ8nKWk5MjqvRoTruC0863tDMmXM67f3Ou00ClTw+RkG
OEfewHHY1qHH4Z/s+vFuxZP+jVvrqXl4PzMZRZwRskyt3V84OIiV9MpKLQxIZLh4nemLpxsv/ZnX
cvb//H7zAZTnK0pHnIF3QK1MWy/CvmLqXhSUX1yvIiHnb67QKnUu+YBj+JqyAo6YJDOXgXJYJ/ki
Sy+eqQUveClJy3XugySQVQ5FSDORaQWN7/nmkeSFBvtJmpFrFjayyIowcg5TfaLnxb/XohN0QNv/
pk9Z/oKiYl693Q0lxd/s5s5gV7DNfj6zhIyvLC88bVNk1YceI33tD28ma4DFIItT51DKdgwvaUXK
d9gXHp6M0S4Cf3x3FBBR24mynVJfZU/4f03lG0x9yYGbgd4501Ipzr2ZnmkRCU6cYnG8T/Y4qWvc
zYY6fKcY9oaC2/nlqgV9tL+i+I5qsoiDd3G7T3VMzZx8cOgvjr2ISqJtO6h9aDLg+QfbXC4xdbOE
rKEDxLAIgPB+fIfK5NWoH0hQXtccckpj7rII1dbvRFtBUpnTP8xqV2tuylFwqh3DZvwnAtyn5Jqw
BPdSXNh8r+eca7hoAXbA3M22XCmjlQPydr22bIXpZ3zQSjjRE4GQB3MlYQseC+dqBjl40/nYCVAO
cHw6lh0gJXNgWrY6IcEMqGbP9iJpkFLafyTnMgfY0bMZsn9CeE1K0/8RKIuhnQOeNcrLJgX0V6AL
Ux6OML4V5ofVJTtY4ihJCnDpwRmuQqivb9Ojh9s2r9P8QX+G9qNoEvAfkwH2YF26zto4y5cT7Df5
Livwb3xJdkgCPhGvb3r7dqNGsWDXp28A0Wd6/WeMVPNNnV51548onugsA1KDI0Un4JZmJpar4UxK
Uj06G446Ay4ozhyndMzV75ZlwNQ+e2pLAeo4tAYwsPGMGFlFSJNQ7J+fIZ2+5fnSoDCDKNKo/CRI
QLUxpeuDG2QM1pLpgtPO7ZlLdPVR8GggFgAQdn9k2MWw1kOGy21cusBuzKS3ClErucMha0TsIKnW
I8nmGzWXkuu5xL4RD94srvvztOnAvcZOgrsIOkDb0TRU40se73E41dvX69WUcKiAN8cLH/ZnEk5c
u4Vo8HvX3lKabMTJ2OAS50IhBAd5FDGQ8vuBx0hFYtn8VhDk2COIdBAWVEGyMe9wAqQjjrFzqXFo
nwY+W6/turGPrXvBWnHCqNex0gIMrpvq7NlKSgpIVoYaR0VTDNMT14ITYA6hs9iuBiEAkQqpCTeL
ryqIy2iwcHnsWWlPd9Fx+GyJXlOstQJHmoKUFtbuRZ2ipGy3jtVQUiGri3PusRFY2rmzk/k63m3x
JfZeZjuePP7JQaJPxU8y0ryESkfjlt69fjQrVED/yjcM791B/BMws77UEZm7LRtgdBDJru945nLS
gFmtml5oIgIer5dHlpMGvs4xibVw3i+STBdyrdMqh0gvKQdycJeWT1XqJZkOSIta/yhUySAj1Hnb
a2ZdoPECS8TFNaM4v6eJ+900F6jg+2dl/ZLtLnZOKh4KJGmwrfhRhyRhkpG0LgO0JK0iRQK2Q9qG
RSr8MxhojrbLoSsjI6jqloubEg/D5sEXJ2zpDm4ND7LQRjQaUN5vAiRahQrUgajmkIgnO0IHzPRn
PTGWziKDL6ab5BImDBmGLo0XxPRQ2CeLqhP4eFn8mp3Nh98fVlLaYuhsIKAZT38ZUo1cD4qYHuzJ
WBkKbbhmojAjvKea6RcK1DHZC1QaPK3U3TkdYl3JI6326a7LzeazZ+6F9KWgoxUVFXd0u8SBW7la
SvjSvvpAPWUhDs0crovGWMBwOnrPjmvamFgFiFEgPtGeo4/HsM7sYhWtmch2GPL4NXRgQkRLGBEX
9Wj8j1BF7eAL78Emw1+GrYG9iyzu+CHPPwmXkCjr5WhMTf+atgp7nCHQIXPW2oqQ2tLWuySNddLf
yA7u2lKMHCrrVDPT48kwpYUvNDrzAjSRLcMjrJdqgM2tCO7tsb14BPma08FkGgKWA5FNj4qjf84P
Kmt05KeiZC6wdz/QJ8JA60IoKhGlIdpXMfbdBenUFTFbnJd0QbHpXdoRGNduT5vrJ9kvQUsfL2V8
aOS31A27BYB+ESn1+YHTBoOjSU1lxMvePZA2594SKu43lYwgAqoSGjDY00GqGoJwl2LPAQfOgmWR
NW9mTicLzfnbUfhnq/7YwJjlPzuPxvHagjqSBHfHOTxp4l+KXoxWB5bRWQ2+ZHcLT7N7ZJ8aUUkZ
NyQ98N57iV6c1mwbKptl5SEoSmgJ6wQwcMVRQ1blZV9fpluHUmMRTO3PFlAz3Rl1DgT/NXBOO+EK
9YK2Pp6od7S6QkVOhQFTsf9S6TZe1sf0p3EpmOdJxuvyW3BVIxT1OqYppgK6i3mCIPC52KwyzCav
w91phk+Sw8j0hSrNlXZEu7H03YKEVumMz8zrVnMUSDRmHSme7ads4GRpROUhtFGzbi4wRVcnC8oE
KETkI/C5qcXQ+tfSvADHkRvtNfi1o5HmF0rQ7uJiIMhfciWQOsbeV5teokT2BTGj/IUnglQvfZc7
fR+aviPgNhOoE4BLj0HC8m2oDFhvSMQI0F9Wyb6A1fG0jZmvY4TaeSsVG1O8+NXThxtD3jJ2Vza5
IAd+RuKFYmnTJo+WFjnWJNZGq2HmlqRP5/+T7RIfIiqrHgTYSpklk8kYDoalNlCoTigSslbFNmUU
jkq0eMBsvrvUdos2B5RSiBtnRLuZsXAhNcynYxm5CGDYl5X1NaG5rb3oODUPLB1SEx4e5EpBzAbN
wVcaT2bYe5Dcf6GORevzva8mSskA6r7vBzIrzGKCM7q5xof87NxzUFe61tTa/qDR7FmFEde/zRzx
GvokjPg07naumrUPp01VxlLLT3SpuL8Ik3Tur1DFskGvQVEcIzNaY3E/n4Aipne4/jaC11e3xun1
HpzLWz9qvs1Ey5yGP/90SDCkztGsHBlgp2w5lXhjez9jVqHECv/xELX9/0OlYFg1XLxmBtC9TRZM
JXYYETNNeaZaAV1rzPCevhFwmLqPMD1DEjdx7eaxsIkNB/1TOS2cyhr3lpyEekf/u8r98Rpurg/R
YdOIaDjzd/HX2VXRlqMmbcUL+d3BznFvgddv+wPuDKVvNz9NatLUGlDKBQmWp6+872lvC1dBh/re
ojWrp78XFlgZwvrLFLil0HQe1OlZDXpHWUQNPbua9Mn3rKNxmUzeTrGqhg1H0ob7ZhiwBlA+FELH
RO0CLR2DhnnxFDuolNX7CYzW6QO2Jnix9ZKJ0e4zcrMVC5K+x0x1vwnVQ2LoXtc18wUMztT0sk3+
TI5Xaq1N0oAFvel4GoTIo+k3OAoWGdCVcrfIM1CZqiSjl/G0xZ6HfxQqllbIhQV0NdB+i+Yd6yes
A7I9TCcx3ozRcXRcXrMwF1UvQKJ/4TSFkec5ZZhSpE8Uk/FMXy0Ac4uPtiQuSkP50L0ASsp/XSaA
K8s7u5FIJTwiJz9sa3inFiy2vovTY2+nOHrNCCr/ND/fSooeaYYyMiVzTMXmRPOnDiqHmtDfpihw
TCHj6ENgnRNtEY3zXjhPjUZu1QUJDrTwGTjNseAYWcHhLwD7yrg4BMhntzwmY0FDNIwIoWcqCBGa
eLOVgVvVMPlJLJ0Rn0nyBKw8cQiANfiJk0FkICoCYFBcEhoaVQlbP57Ugj2S/d4na4JlyCeSdvGS
zYGrCR4bHcOqfKQrEfJ6AOm/HSJBCxu4AAkusbG7LnqHXea/Qf66brTyBOOaRsxB9Kx2MbIECj01
FlUhxkmAFxKVfNTODBJc2Lb34+SbQHV/M6ZzYweSm9O0FSmWytrpJQepcpFExQ5rqQHI/ieqixc3
K1mEOBXCeF8QYvvZ51h/V0TsOmcgT6yY0LiUzdz0SaBzNMVoqnm+clQWB3og7rsVNREj4TaK34pI
yOOCzSGzxY4DsMNhEJzBPdyZ4du/sRCr1oOnTXAEl1Zh8WKGKSMYp4MrJmpatrK8eN5LFEi/yLFH
L1ziKmlLDd8dF0IsxOGzGQ7WUeWOlz1r0TW7q8Y3YSh+JLWJTTGLgXe3hv5cwcACglOFdS9Xhiiy
hzXJ+SVntCxnmaHfBWDo9ZsIilheReIB8x+9Kn62WVzZQzzezA2VQgzTqJlrxTaQ+qX85f78DC16
WxBut8gZbIldvDfBOV6lbazu80zkeLhsY7CzmP75P53n69OynQ96fVbIUP6QmCxWlTceL3nl3A0y
WVl2bGPhyG4b+vMRtQ7KFy7I9QNxDUX0j72DXOAMbZxhb7eIPpBEYBOTAGHbnytPD3ucWRZP+HPv
ofJ02XjCcZoIbj2UKGD2YBhh/I20VMZ4wqLQ1ASb3uaraLSMiptH4uRacesg63IHb+3zh8QcXusr
h+2eMN2Yir8qHsvsG4rMpf9UDCnDC42c0ZjfHXj9K29LWj1kvROnkKYOTExPJzpZSP0cps2ioD1u
HRr7kSkomVSDxZfuSNMgEeVO+WgYdm99VZ2dY9Yp+yOt9sOaV77HDGa6hc6us/oPM6iMhL4AaeDY
LcJLifLbB5xud4FJe5Vd6NadlWQptphNwZoJ5GMBnw1CpRar9riSTtvTKiqSy5QATMP/TOddUvYk
TcphgZ8naE9XyzcuKmkZHEHUSWWcmeK6YkPcTk19WpfoCf1WHyPcGKg5acAh437yYtdRs+IaxcFP
PyWitmma8Bq+LjuDjOHQqSay1blB1TYr1xmAvxE10TC1sQhgr02BbtkRcQtQnwn1WEZIFUqwC44S
1wsjCuj3HqYVqtJEtwh7+V7WzkfyOIJEwEuq3XNfO+QI9U+vuJx6xXycDI8BpJ9SO21Jv7mR6B7d
CGsIGHx/esmAJb80R3t5PWxyEk5zlnVLWUCqbs+bm1kHvkkR6r0R1NPRaToK3Mj7nYyCY6lTYcEq
j3AP0zzYYZVvLBu4V/04gry6ySBXRpro2EfscpsGnEo9RMzf1Jn+ypQpKW9l9okADutzTZ36x4h/
7Hf6/uRu+lyd+RQnOGqI/422CxGL8nxvSecOGFwVdCfAo9vsvJIZaam4IX2zuFK6862ySg4CY2gO
kC3yHRbIjfcSEz4Vv7c9sN9jDXaUMhysTMuC0iCQdcZiS/eUtI0tTx3+AHjp/3eTb1pBXhTfEzeA
FJ7wq6NcBivtZYMdXaguNkRAI+HizAcjlzdBMQ8u4WjBPNkvmQ6FVkr31cza2esH1bXJTHxa/QM0
oOPMWZVIs6iHurUijQqwdFjL2bRVYuk7oDvBAQ13NZciMFZmHWup3k4HqpZW/4J7yArdRgiH3Rlg
FDIXZMz4JufP98UH1sLeYMgitZT0n5pKA8XgLpC5AHhZvac5RbsEW9H1qcaP87omn1OI6JRWQ0Bu
sF0+KQRCrumRLPx3Oo4Spzyabf7SSVxSrbIF7vzRYb3HgFEqBRIQfWlwTlbni91YUI4VlGg645K3
eKCMVxOCxZxvX40FPGeb4MbbpzoqZrMEZ1TPePqih+4gruxbmH04eXu5BXt6+Y92Ez2z7xplqIPJ
hqdnkYsl//kKFjXZr2mptXLQ6gOhxxtsMDgGi//uq9zFWrlVeHLFqnLenQg4RKEi/1nqxT/KV/7o
+sjztrpy9cCdnevVsd0/RwXStjj9w/su++9ToMCQatNZYH9fs+BSMFGc9c7DAV0q3y0JmeueKFlL
FU8wzB9015Y1Q6Zwm19th3lOYAIKvFFtQygj2eNN/zFlaB+2W/XfYP2mTRu18bL3Y55QXEEc3cx7
ntnZqObla4r+R0Dnb3nGUKF1DFmnmv1zDbSH/TidHA7rkXG6AaC6GDzkyc/8ENzcRiUBGaQxydkz
FYgRypJXtDL+vFFZHlNm/qgG3Es4qCGel0MYKKGdgh0LXp6ki5Vicuh7lr4JFhpUhHCRIrqWRxSX
V78IYUGmhICEAaYUrwpReYxtdmkaioRKuWyImgyTBgkQsKdWuzieZJkZG0l7s8/AEyGd4xBLjkdP
8DtJ+4MA2lniefrIMmZhd66prKLrN3tZ0FKM+qOQSOpSsBK1XZgdEnLcQGD2PDUvliK1E8WNKZlw
NIH/W2vJvEkJ8WKNlL4LoSdcUjb0SA6u/8esDsc02tYKzlDAVhmfpEBTWwqswfkr6jml50O/7ozA
93VYCMBvTzOZcfcvNYtuV/on6Dy3MTUK0i19ds1jC3qLs/75MD37f7uH5XRpuRWX9rhQTnEwQOeX
3UQ/7GvRVgZyM6jRqeSTArNUZqPRd616lmFICbWou9mZlCmHH2/vzikW0Mo6CivdYwV8K45gicXE
ncLxZUMIGCGJJicdIW1fNHm5l/EayFe5Qk0Sb7MKqUqQ8FQa1FOZgEpkEfo59RYNN7WB3eUvfMnz
dvm1mwQ2ld8/kKJPESHZ7Q+NkUQ6fufpkV9iSQmgsraezR6YWgTO1FshAfmoueRgOacTejsUyEYM
p1pxMl0pmTOMYUyPBvgIPzkxl2OnOYBA/Wl+znolw2oW7UOpjyByBXm9Tpc5xTCLDBz+kSCud727
5E88d4wYIqAnoCueYQa8jBC6fFKfzIB6BQC4Jy6uRUJ33CUKkOCpx4UHsymRUwnwyxF15/WvL92I
i/8u6Rck8X5QiYmbZGpJeKHY7Zhr04Gb4KUIz2K9aommvLyxYEFZ0sVjw2MIS+xNDpIEnIEIZsjS
GInXu3sZXS9bKYHGKxbHj9UnxAgE9RnOOVUIOmMb7TBKolBEaeZjpGO16veXv8YhyLXCQZxw+/BV
9NWMue5O3Hu9d64b78gASgj3uYq860rnm0/9Af73cCIZKNkDYiCfd/7DFmVX2V4krlPktovDyw/N
SbEHaes1fihZqXg6F6l4LenOSMFDDd8z5qZZP1vNmItAKP6ob6v3WErVbIoM4NtrxD+9zOGT1x8X
9OMtzebdAoLlxDMFBCsB5RN6jQYxP666flzr9DGBX2pvn9tNJiduZZoRVT5LfGWYhn4an2GhdoJb
REBen5tevbu+GebvGYF7O5TRbs7QB2JDySMopCZKVVykPH/wM4JiOdrpT9YGodRFNfftEcQ=
`pragma protect end_protected
