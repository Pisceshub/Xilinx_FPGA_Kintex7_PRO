`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
KknvL6SYSb5dRFuWP4AJqBhO3b64YXO1jXJrKEg0Z3ikGAO3obMtU40YwJiJW7ipQ08/Y8WRYNWh
nV2LdqH0dA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QLUbVPatcj7IWeOM7GaVpOxxKXKrfEAPdOAPmfRnpcapAKHnvWUhcysRYZ/rY/73FKWInR8HJilV
JFgxROZVCNWQ1zJhGgmKt04WHahOu9miHsfm8H7yNJ6k3TsDqjbc8beG5UCVgF6x/gDB8LRb2Vlo
OYeUOl3UjHyll8Sbd9I=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4fDulW+j2qCXqz735RjXksliYlPtal97cQEPC5accAQtxDw7TbdSqrHOiG5KctOIuaRzvRMOO5x
8R7f4K2bkMvIUjiiFP5Xw/fjJySLFuOiZoiNxxNdz5n6QQgBWYDepruKbEU7yj9zlmf0zEFmWZo2
ShS1WpLwP3B9Mcm5hJ+0GZ0wSeVmrvJEKp8kqO3uW6EVpKbiSMmBugVkGUzz9ZrIbzEZlELi+wJ/
HVgQM4hNwGKaRhAKNMJGLkgs6Mi/pI+CqjdrjRYK0X20OxPYi7+y3i6gUy//rkWJVRVSqqxJt07h
XfBm/2egXCeHNQMVyg/cuW80bFPZUcKb/tb28A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eEHF/HRqboErONr15dWGPiKIhHmEp89NzpKM1HVNOPxPMAhm5Q7SHcs30Gyp606YzPvXAWOwIhp6
yShxWJQDMNzjx8XLNdk6Hk4q1OFOlxJvftzg6IwFePhX6CX5M/h6gWDjhSncOnYuNt1s46FrBJGA
DJZ7AbtD39aEQbpRrtRqPKdh74/RGoSXOsksuOHq//+3LZGY5WN1wdVNJTew5IKMLtb98TYlHOO4
w28CobD4NywkdWMYWBeN1weCfLySyzftQavfk/dRUoBAG4mBbSm67pDUnjTuzD/BMIiEezbjKgGt
v5JKng8K28aaFylCDbrjWbQ4f0E0MG89P9bqcQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LBodvKMdQLsL3NITg6iyfn6uEr0nsFsSECbcpJ0VM9GPtNyhu1PCIqop74QUK0jX7gNod2kXTA0j
UPAVU1VbFsW+W9odvoIvVhgiIvptX2ncKxVnQVrYamDTZTPdFxs85ZcmhfukKF1ctZJMx5QHtsT8
/fgDo9EnaiAwUK6EH1vPn8nlJtMakUlaKARMU1hnWHBUkjruM2J062f3fYCx1Fc0yI51VXZXtNw2
A35SpeR68WKPmXnaWtRfYcT55OhdStBuASxbBHMItu7IQi56vUWP8LJm5L8r7e0VPvAGmJGTHM8m
DRb2QSYwaQDB32Ac/WNT/HueDTeVlvRT+cXLnQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RTdH2QVRkLMNeDjWHM39MNQI9JpZeMEnnaFqgJIEgBuj3R1/oXRV+h+0yVRQ+SMug8jz9no0jCSS
W3wRM89ooYAXiOYt8RwiQibqZKat+R7T7m3thhmgMEI8uoi9fGuXrcwO/YAOvNwNOuRc5iytwydq
EbyW4aM2m+CrXKFlD7s=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hNd+z0nXH9GYvgjnhDJoJvhFhK8AT6oUoCmTuJoXrdeSPSICu0d2AmfE/9zKTVob1byyZNQ+dZJb
Ma+7SxXV1+3xFvececBxzrOjVMq4geH8T4yeo12KR/tsEogGtiBVtNuwOoiOTxmMqj4v1JDOa2o8
G9PU/lTBUSoEzibdcIpQyhvP7Mdz6AOWlVWthHuCNvffk52oBkFkYg/wxqRli9uZ+ljnrd6rXIeN
pcjEkI9ALbBEAZnGGMY3do4kdn+d4UrzbiC/0FwIrw+uZYeWK2+A1bCZ3JcBMczd2lYYJYQOACWj
1dr/Sij9Dnl2NTdY6Acp6dQAwn2oASr3Hs8Onw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 44400)
`pragma protect data_block
F4D6nIAHG9w7CzDjTOGl45rj1wrMCCZxpk/PW3zCRBHortjn3GKkhEhSOKF1o+is9PbYawqiQGXB
iBpvYxLmwMM93kU6zXlXi7eR4gCEzblbk223GV5+hBrY4vfS4cmRQFvhTtdtgAnRMqKIeUwZLiWd
o9O7E1ho9DFNkr06v0qw+JJ8FFfUjo+w4Y1AnAXAOSHK4ie1KJYwo7yEI0pqkXvOEoBW9CVhQoFm
nU6wPQm+0fupvziyEwJxGR2sihkzHx/FowIgLcijdT6RFZDbLAIRA52MH0Ix7pmY/37vWjvxX0uH
NpYqQ2MsqP9udJuSy5syRLCtQSmtw9+jBiUDoRgU+VZHtysswupdKsO7AFLC+nCxFl/J3Ir76P96
V5xAvTaUkKy9/kC4L7JaovCliuH4/uLdYV59/OYAZpWYzDACFTDkNjxUOuZ2qYaoMCcpo+XKReRx
s6fFmnSUbHVLz0CASh2Xd2rrwBZ/20NUp+4rIES8N70crHr9b8LEIvnW/I3DPu2qc3tJVxtpzLbH
Xiukpx6Ow8p7vZmxxi7h1dQm7NqJaY33P8luqp+ca0uZQULv8fTmffzfDYfqK16QeO1GQpCQKKCC
nXpHbXynXcHt2K2fyzG/vrWbsSgOAh+p3Ub6lGr5CMdCAm0T/NKdEgU1ysdKoPg1WP0aobK97QsH
CdjjqJcZm/q8lupEG6VLSF0LnPxa6lLHtgFSLz1HlJU13g0WgmGP5fjBr6KHnHvmbFDynAWpI74S
TYU6JxA3supbtnTTgSCE+1vnt8HJTaq6nyvh5VwiqVuLa754OVHw0gBAFOlb55/ycm3K7eQbPI7P
I2l0SILYsS2pPiQzrSboMg8ytXSvW7ugdF8ir6G26WhQ62HK5UACb2NuzprEvjFobNwOZU6diN8o
4TdEl6CvgQMoYjkRYLNP5zyumGWBtU2XxyIA7gqzCJEycIuh7ueWBoo3tKNG9/g17v/V1TZSb9bo
2f2urKRpzgAveJEbcUNhRfRs7wWg1Gc+UL4aeR2u9AAFZBLglKiQ6cEq9OMoewSER+5uprhZ0Zh/
ODsjfcY5J3pk1jk+ObJbJmOtB9fm/yORn8PhQ9pQtsh6EjXiizEgVUjTejKfHw7xdjBiqnGCNP6G
/jGoP5wrh/7d2TZ2hKsDU/aY7mrfCMEOu125tWVmxWTwDZD8qU4emsDnpzq/oELP06DX1chpkiGE
jYnQTPawLfzYC44NWY4nyZEd2OLhEZ4igV+i19e8pGkWcK5tPbR1fCc7VTjqvOL4GioPoLnOhV/g
WEYRALm7+wQUZUG79HJqdO0aj806VZStsbyl8PtEmr1AHzzrdvDP0GGjUcNlQaZAhUInZoQ4uUcG
sIQkOW7YZkRz2K6lI/GOQ6G1kZUBG0PTSPcRGBMPwPldRwLgoUuIzjMHoMzeTy8lAbn1jN6Inffv
HeYLkT3kdseot/3Rue5HzVQSqnz0eGnaZUgBawRFSEBQCJpgQ+gUxh/k560wtLA8rjasyxhYZBgB
9CzwAML0eDGPco0fb/pAZr5TwXdE6ALbi2EfMimtlZyp9oE8ws+QSvAwNsn4SDtHbLCvYK5i50Em
W/KVKQfwHz2rFsZM1sMIyorx01V+mBXWrSjR1+wRxnuZrazMpcaXQk8drfVq42eGwAAk7QgSimsW
1Xe3gw7Nca+nuHSTMiUiISfiEGJtR9ZliIfx4GXD+vJhPFy0YAsh8Dvn9Eci+RevP/BAII4eM7uE
nv4BZVUmxpD90d8nttVpPxn0UqLLICIkPPXPDgz8+p3ImRFNQDm5dxf2qY2DKdbrYWGiIg81tT/l
1s26fxWZSdXN1KggyG+0yrWG94RQwLss9Eradv/bHaLxgeQ9/O9ByWeNny6ngGpQjLO7Q2BG6q+u
8y9QbONJN9KHG+FtP2Dd43yz0Ims7tqvFqkzuBDo9LoQN4tT82jtojK2M5Bb03Oeckzrqrkdlxt7
gW+QqJOQI21SX4kAkEc7Y3m4uHuvpRQ6DEdOXeFAx6Cn6N2NrdneSsMFi0pctSxz08XMdpS550Ri
2C8BmAMJuXr6zt5oHffGX8j/6/4Oys200apHnHQrQcIHj2OeZ4+cno2cuw99hOuBD1kHv86ccfAW
JWxm8KqnjRJTo0lxWwmA/W+/2DIOaqEE0hMUM2qHu0GnjWjJ7jfwZnhLoDIpxQ2fZxgYQTCbzDQI
2FY0Dtzgz6pxxqXOC4dCEVziKzwJP9ywskQkvS2dXauls8L+HFhZjoWa7vjedx/zPrr8pAOa5pvr
Kg1ziUUWajJIbdLH0cakENFs08OlRW/IkcPKRhsuIvuaIidjQWvv5EwKj61S6Y0eiPverqKZ3E6p
cO5Vmk6VlNBlw2HzN3FIj/0LOoB2mfFpEPF2Bv5okjKHDIPWj+xzIiSS/lquAdyebwx6bdv4JRx+
m6WpOhZ5tFQkkgCZOv6cZtWrOz1NtmAJSHEtJGybC0ZhUl5/ee5498h7PyWissGXK9Qj+3F3sE2Q
yMGezSilxXbVQq/ki59wqJKA1G3wQ5MqOlCQi/JwmVKUCWMkAlyB2jh6lmK1O7AEJ85866AEFnNT
0oSTtiC5a/MjpRomBP6j2pSyB39g9e50tqdZ8b3LiMSNrZg6NZk7zKSC/8s7GiwIC5KMy6IFksYB
X8XTE27X+8LwuOomyX2ILwXBm8uaVhKliLNuSFNf9q4unq3b5TM+ioWrdQRmUra+HUxgG7ZdoorQ
ooAYxTIblkAOcdTAcfFpmMeR/d45zXOySTKVsLQcmzrPwdiufpipzLIOMw/jIHAe1hqR0jnQY/La
MSTtxQnw9EyO2gCaoT0mfUZyVRb2n0CSx/quEUUWY7tK8wxzRFeRTVva1Qdfph+FEey5SkneeA8W
2fN+rAWj2pB6+LQaZY7I6sqPPDoMkHi68o9Tl8VdRW8W+mQpcrg2ZxGIvMWLTImewP2ISPAv0Lkf
Liuws27EIAV7z9E+U0I644KyI5eNHhYrAO85MQlz7/hjtokntZtBUuPy68j8bdaW1g5/MPdl6pTR
F+MxMu4WcwC2wLz+sBtFsjJX5AbKWbSlQT/23PVLOHbYWcsgyEZID/O+oNkIVwkPgmpfcgN4E+EY
abbONiMZ2i7SOXvGZoTSyCUVMETGnyAgEDbEqKB8P+H2WfBQKhFBSbrviCnmZshS8iEn+5O99I1v
KXPWxLqyFov3V62E0/atS7XEDtkbb3xtB8o9xv/tLJQxvyaCu/x8C++0LHgoFpZYbJ9cJAJ2A9h4
keHIWz+B7wvwCO+COyw4+wJWrGEK4+eQkYJeOHjvLVWYyXMLv9KiUyCMpDkxdEc9VokWldWKuyQi
52X217mhIL3TN5RV+nYDlheaZZ7Y6FO9QJOHayAOlFHdPzCGWi01TvqVhENDroTdGpveGAPdYFj+
eaayA6vcL9glCheRqTut6z3/Q3WYqEvsjh8hpymfWKXdjvw+8Vap+xuRhkiJMzqcTDpknkR8bwBL
fBahhDfAgehrO87iQuJE9q91sY8dX4mbyIyh/yjPcFBslqT3bRwX0t6fgQ4+GpkqPdpxdkKAXjkm
wIafCe6V+opEnjTXOdbYFsuc8JnRqZGejIeHVSNl4w3v7J46ffkzkJtmP3F0GHxHhscZUgGknUid
27OYcI70DnAk3Xzh9jIh6nefSIpDOV6DlellJ6BC81BTJz2SoS0gj3UNsuRWdKsUC+dXG6/NNbgN
OsUdDU9vsg2hMjcQ16D6t6aA0GWTbWsRTJgJGgp2+zM3eJEdI4uHH54iq1SElxpkUH74aObct2DR
uqcsZvj8XkqdJhR1+r9zrhWhLDJhBuy/CxB9uu3Q1RyGHXZHnWyrnBCjzRHTg50sIZvfVVCFxVfW
eLgSiP5QbUoQVVuDgBXj2V5zcPSxLn/Or1k9gmFxlHhg4qwMQm1FvEyTZfDxp8CKWHt2lcbtCnX7
7yAx3qFsPlhqgkHj3flzBVSeEVN0U2TOo32camhxk16A3a5eLjzLH15SGFIhRQXdbdGMCyPzqFRT
kZSB+KfWdAtpdz6RHg3CH6J5eu4bSvf2Mw+EpltU7+EVpWBkrrJpTYWD3jrlQytiY5M8u4795Hxy
0M66cAAbNQEEleKaaME6GARBLPLxBmt+jrdgnXn99+/T8HuJtZ7mIjtyYpPRliJNFUGxGkUI8gXB
/F4wlxOvhPBnL3RO1B+aH1tJom5vdvWK/BU45tD99+9wQS1md0xxq2J5rhRyFL+89hKspgdYFnc2
80ZGidf29agr9imrKBGACtCcIPOE+pR+VQHr2f59xk7i1r4LSDLrbDXNaZpE9EGgApc7OdFkcXeR
xOo38rXgScdZbhFzmq7t42U9FKyML4NWDECVlsoEzfj/PISq5WGh25Anr0VC/Z1sdz6KDmIeuRxc
q8qtxMbkH6YGviwizV41YIKJagxLhKGKVTPeWXUQcKACvl0xk4WO9R6SyCRtc4LaYvwgubzDaHgA
/4iGNLCqH/JvgI9m4uP2ghrzHZJGNurFIQCIZqWEmov+Df6jECfiOzxxHcD1JAPgONsKrtDzkbiE
VElon+5EGPyrFAuEOiSEzlSbfh8fCyQm1EOsv9wFpw2SVKGgFrBHleKLYczKruEPEycc/xgct5A9
5+kJLLK4XWCVQTlJGgReCTOfspfrFbq+1/40ux220c7MhlV3AsS9+zS6CBoK1cZcF4/20H+3ApZo
Fa0Y1+czokVwu1nGm3yv/0SytvqZIV1qW+Qa5pCzZwe/5O1qmUHoD3O62lp9D6kRYwR3XBSuFAhI
Idscb7guGztn7QCQ675TwUj6BL6k/mKGaotnH1t5Y65eraQk0DPgm/xbFjzuQLbTIF+4Bh352tJv
MLea+kP/qOZr4E8VedkmvcqQ6pDEVxC0LgbVZRdecjNJV8mBL+T7vUjEO3/OHbi8Fi/nLHeymgtD
V8albC2c7AO+GDf2wxsdb2+Fo7VN9cMJhePHuhCLklgkNCgN41FQ6oNyHvES8Khj0Gyl46wcGXuL
rd5Ke2sEsU/kThmibS5QSKEEl9TDWSfZkdcw61QUEe0CHUeHaxW+GqCd3Edj3Y/UxmuKHe8G/HGm
aSjxzhRooPD7FO4tRN+AxAbhpP6/iVaPj8i3hs2y1dmFT337aPsOk6XUX7COu4wacwKWrc66WdlA
+lR/gWLm/KyOaQzp8bOCXxgS7dy5q1KnL8zn9uq+Abr8tNUuVVNxw7ALz3GfvcqSxLgKhANKodmq
kD8bxDxVPcgruSoZW2ySn3VNB/XJ6wy2/cEjZksQC4aLukpKIXuGdz4/8bX93gDYN6rm4NUFWh8J
Fl6bZEIVnwS+ZxWodNLtSNoG4UW0s1DgGmGO0fNAORkZIvea3wjxOZsBUnX94pmesMhJ298d3m5H
YMi0aZ7uLYBKlPaVgjDYuEhvW3RV8lZCQwp1xEua2oKnx6V5KQ8RTgX3lIqjVxCWOWuI+CLhoTme
Tq+irHKLWSCp/kTBQNRjDi6A9eyCv7HvtM2Q1k+r1sDrcBGw2HeWXRGWmEtWUoUj/t7M5ytWDIuX
+2SDOyW5wpOd8NoHi9ZlAKlasPbe3cYOql92S/QydyGgR7nUkuuiJp0Qxgzes5XepjNk/xc6wMEU
aXM5eBK5fKyC4/ZLCXTBn5elxE1N6bwKnv4hNtbPngRCEXc5sW5tem6fcIL1ZTF1EgfbJpVacCpz
gUwU4x1XgPgqL/PMnIjOoeq2Ozf0pPaLwTYIR/+FnhPWF+KmxSl9drW3WGyoZTzk4TKI91bmQYpN
DvM0xewa2WS1ULb7SePk0eUFmNcbFV5uCv6L4uRPCkxb7ouxnRNcZesUc2vUPiK/YgNNFOydg4Ue
xnWdVfO4E155x/HAMknJ0PoC5xt+/QkpLWMEfeXLtHetyB6AmjnM56XJFt1jIOhW/+avMwo8o9LL
33lUMHNSjmE7SJH/saQqSSWHWiNT+UcALMHV/XCUNfZ42rj+lg0NRkCUgqUDMMDqV+nlLRhDs8FV
tx49MyZZy8613MeVX0I4yPIF4b6c9Xub/TXsgbk2XZotctGBUllhvy3eqZrK9/dyJcC98pvHs/Yu
2plK2enrP7AVOuRYgn8Vdt+U9/rDE9j7ZaPAU3apZgwXKqr9fnHoXGFu1INuN0Pmj9s+ZBQNJfSf
sPjG6I56dQQjBofyZnC1cn8V2bv39GOnPMqKiSaPC4ypDzK25qW8YVMLsk5X0MePQ8MD1nlYH1iB
Vko7eIbu5DqWFs5gVKl/DFFzpx876RxN/WXYD932+bkHKYMUcubtXGVdkwdWr5T16CflDtRr/dsS
BdlOq4tpVR3u0FDjIWopahs5nBlgZDn6kn9OT1tKV1ZqHgJ5mK++GhgbdnL/4cWwuR6Zk0d/8h6Q
2ndphTw7AG5Zq2JCJVV7A1qvYoCtBbTkgKe0A5Sus9mn4K0euuFmp7qczofY2Knqra9Ysr1gjCmt
P2KJqZHT4hkpZ91vcN5BE2+VbpC5WWRHBWSayhKz16+m7/bdR+RgqDFfsA0Zh6JLFqFvxS7F9bGM
dPg1zYus6R9cZ7zFicCBIvh9ndKUEDgnibUBaALN5tDmRB/5+mSapWeL7tQq2tkiCMrk19jQomkn
il60bpXtliZXLI9iMaOWmANIP3V5E9yegILvW8xrtGCjfXOi6NaWmfI6+/P5BaWbh7Mflvj0FLDD
xNmMpTNn5qItrfgFfonh6htBroiZKs41O6hpnSbTNUaNkHyH3nsroS1wZy8C51FwpLRTcjiapDQe
iXAHpYUxPueSOUyhmm0LGICYXZNx85X7fpy262od9xE8DgUP17AUQag0rJSSr9Ob1MpNu6R2Zm5c
6sNv8PYMueINnZb+2ENOE+vF1ekrsPavnb+MANE+MLoBT3SFYekWuSeaH4gDjMvUcQX6vlpZeTPq
KjYdrL+66xUj6Zv6I/ZQfoWqZxzyUtOkvnC+F7orCE0mp49bNwqw1qFmpb8GgSwa/naSQvwSp94H
oVqPbrpWWr2vjgHs8aso0i2R5iHdXAkV55pauJ2wMBnF6omi5k53/OfDIZ6mxa3hOZHj8K6xmZOI
eZC3h15Kgve5tpp4TPQaUFnLfaYXLu+zZ4q3dC04z2vojfnSDagwErEMKdkVNeit8B/CjjOtOQmo
NMUxXu2VIKEWr5GhMz01WrGap59FIwN0kUZZ3DMFIb1kUy4ODsDjDvH2RQ1t/XXSNswaBrFX/4i4
DCW4HGw9+T5qYLO9EFYdJZbdCJjpn3nC5e+HAcQi++YQq7T7UejcbTpHaZHxeXORU7XgGxmVFNlM
E0Lu1EBS6SFWyZWPMlu+08f8jKEhqsLTj6ksg5YoF85IRk1Gg8sRkc8u7un3m3gOi1XL40a5GnQ8
mlr3fDH002hMhBopSunyStX+3/N3vQTTYZatsk8+S3GNxPtUNKAq3oZ2NJS7u2Mwjb7h7V4Prmka
3M6wicuA7fGlj2nINmvPa3CfdlhCxxZ4mN+1U2FOOQykdeDYe0IpgOXK7V0gVAeKSBdO89KdaP+b
pCu3/iYTIwpVf5xsAUUYVkbCmjGJo38lmHbgkO/7t4avoF4BORN3Fje7/FDZcVbtEqC79WgS8iXW
J7EGFxhFm6eLAIDQa6xLd3KO4HGS7z4L5rEKewDJRBJuydYBdFoAMcWZfytLe2+nD1L43EAufJLM
FfZizEat2iNYQa7tU472uy+HbdNc7R7dZr6P5NIWDgub6LqCBfQHFu9jF7beJrmdHLy52bPphFJI
lNKHfZIVgSyj+tSiadovKp3xth8tqxAQt0cmSitt216lubktDhltCvtwowD5QMnPwnkXkXVJN2o3
F/gpVwitF+Ma0IK+sxpbjZxVRo5H4p8dcwDFoMnTuW5A9r/s1d9/qvGu/KNuRXiB0vORNEIrR5m4
JouEiQKU6tmUE0JXhZFnQ1iWEsyn1blviKgnEJosuXT2PRpHuRmNCaQKCEoAAjQRFyOGIiBaQdc6
0a4rtjBaIo52r1wm2iX0TN+CPWvcdzzpaT8biVclVv2vwRqrcQpQk2XYhb9CUoNIw1cT32tA3lp+
ODLom51ydOheuYnmZHH137oVbeygXcSTiUHNaXIDtq6fwX/3Q5aiHmTa7OLZ/utY6XZtT5aix66m
dihB2UZeB1lO2Pb0Y3JxC/VHIly6E5mcIe/cb88OR7gYqOKUez22eJwntnEMj6EN+x8gMEG755k5
fp0OL5mnen0dakxov8QMfon2JT25LhomTDEQl9GcyQa0d8GkuoxR7Ep4aG97jtWFdwBN70ZqDrpq
xniIpBaTl6HQAS3X2DL4MbFHtBm7doru2HmBk2TA8PTIe+PV5WpS5XBTMSq0r8LuyQ3ZfaUlikik
YVyfIPqC7s9HORf4F68h5zL9Px338a5tHoqd3nG27Tp7oxSMafYrKGsM8Cz5XsEVrHlzyX3nOOFX
giY3LGwfU2iZajnJDdVs1bUJY3LYOVsrUlqdnSXTyjE//174nmpB6vSF9KltSmOtjFTLOb9Cbo1R
vGW0Ew68tWYj2k3CZ+g0/iEpzhHVhvOhjbi4ekYBzJuvayW+6ZipgOKBfZ3CzqLGSI2ivERnkW3I
nPz/duCp3CMsWpXCoBV7+Z7liyFD/eKf2WrgZnWLtEnQFk8cRXlMQPTG9vlLSN+5hx4NrCWEJPH/
cvLy7HOaYZWn7mq0ahr9jTvpxIV78wwpg2sWmI1xRomP6v4QfqCxtu1qo0f/rOAeqVpR6sJjRZs5
3c3Hqdr4e/CGUdSH4xSJnSVDlgO5jCZMzajtFTpTVIK3iM3D5ZHmxow+Lwt72RmdmL3JC0F2iny1
TSvGfrGjDok2toiZqGiZO2l2akxrWC1Xfc1ChqpNXO0x4+JyDXh4u+HFY5thjQZTiaTe0QWuJZtf
kMY6KjWHM3b+I5uvWacT6SMWLTtr9atHllL/RczuyuqDFeHzEFU9ewoltzLibw7uh0Ks6HsXrxfq
15pAxvsWj+q3GdCUwGlEbK7s8xrgRAxnPsrC/BTe+I+vtOFuWuDNtJpehEH1a+bXANkpWPxX0OSP
vxHN6/pjj3ANL9UCLYsi9hCwpOFky89GuDodzLpIE1nMOOw3TaG2nCqbT4utqwo8ts/PpKoqwQuC
4GHEzs0d41183M90eilf33gYLgRiB0ee1pLmVd1LAlCr3IKMhgWba9bGAzgNwjnTkedmExychqs/
02miEMBJaZJOvq2UN5y+f2CGG0kdTUBxC4MSt4dnw04dNR4uZH7vce0jGOHu/aAF1Mp8ijDL3RZs
+3Qw6+h/M/72aV11SnLCbWwr0Q7zRgFBo88laOuHmNiqb7Z6xIdqa9f6ZcfKAjSQG6V1jmbh3i4m
QgR1YWwK35WISJFvWzjKf8RuOOi9EhViDUM/plywppasijBqduChlWWMPuYe2LW0KOjVZCweiFhX
juBZ6Ch09Wr+cp3I7h11pgjsYyV/UMxHiFh3ktM0AaW2Y0irhjWghoznYrIMpB4of5A0JxRei5qr
h2FsFYqdHLqiOGrLf07sQ2DMbRL5i2ioSLAnCIJIlUtEAiBLa1XgnuOtelpyz8fGTCzE9bk/OSer
wpIH9TWSMxQsZsAP9VDznKXT0l9eZH0K2xfSQb6GvqCBjbtjwPcOkiLHMGd/JsmgulmxVh4Z6rks
whXs29BQfGiJWsm3vGkXYm1tLz+Ji0obFa8SwyXaP5FB/3WVZGYF3z4PwlQHdQ6xJPYhC8zONRml
OzsNWbRjTmPlESEGZJcbYpTGqXIL3QIWScdQXtYWXrHpsPwQl450JaaGQyF7b4aD/a6w+zsyYjdh
3jUi/ltRSIEW2gaVa7q0tffDascHtqwXUXsReqij2PYV3tLbIejR0A86/FgUmy/ihDe2+Hc5Wf7o
xHk73etIPZEtQbWY2Jo2l3i3OO9D7d5zZ33J0W9h9V8Bo68HjyxIAGYNvy0EhweHAJvOAKPJdDr4
u9tcqhd4mCUk3zpUY8HXrSMumkEXvzpLcykqcVSXXz4hAFxFqXcX3bEu1hdOx6AYGJeo4Sm9u7Qq
PWhTELEmJh+6cbj/9BirBcdVWg2xs0AkGyRJL4C/GrAGG4j49PzfeDnBeJzGujWGOp9DUITUkuf4
g2CfAkssIh/UGWjG44Y4BHAeMnlBv+xyBq7vySLEfe40fO7l8HV4bsA4RBmA9aZ9sgPseKWIQfRJ
4USCIjQmzD8/Doz27Az/voHUxrKM/Dv1x9d+6J+zDpQrxX29Yq8eIZNQ2z79FD4rtdLR6izrSv4v
7VtleIwBfuyc7n1Rcy5maWYOOyooUtK9cuJY3Y7LnSg0znw4sCNU5214sf/dEZI5+M27SLDPWAMZ
FRE+sA1uqzFHnnPGN6Zxy2DAxVLu0C+QCRaoe0JcgH45oQrvlg1OgpTJhjmnHnZF+qGLNcwXgVc7
8459aOiX4SD+L1iY33VdJmbCp7Wth/V+14WXlYMMxtsShFzGE3zSxNHUEkfU+Hg/vwMivElbORph
cJY14Ut+FizxDoUer/XFaviR71KGsQapHt2zJJDlla8BVzTdH6d1GeLtDXB5j/+SHIpY4oBqi2iY
4mfFpsfdWfQpUIly2/6NT/f+G719OQ4BzdSyP6kSV92Ens+qNW9shgfF3gV1bstQ+g5iQyVBIzYN
5Jy74vTvYW1oI/A9uvN4BulJdjWENUWWT6NCjZwsAvlHXR2ZN+JetDJzvWxZN8zhCPW1y3CU6Agk
8E0bUR95Ighz3BsXz5k1phzDJulu/2UrH7ist9x0D9x/sasm0kodXCB35RX423Cd7JWxw1u5Dv5Z
cXDUt616xKS2xAosj0qIlSRxAZK3xsOqESoewyj6l12QEbElBvRmDzNA/6cTt4/03g16GMp+PC5R
ngY1ONLenH1exURL1ag/Z1epUITUX6aj1WZ+/k2mHxCpzvWZMr5jC5yVJ205UaosxwsgXvnvpAY+
dgkJ92udPycD4D0WBv4RwdQfTFl5vTAsdDnFAlbH/TrzStxLzhXCxDliZHT6/VE7VR96rbFG+pWm
kDzVX8bgHHl2LhRXFypBRDEDdSo7OaGjMhTmvdGAgUUU8H+p7WC/1HmEEtqeDWNkAVsj7girf9nT
ptyt38Zz+/xex/uHZldga9v13goB3gti5URJ1DeGU5BOwUGNkfRnucqzIp4Obw1z6FswLJTO02KY
jYVYwIrmhSOP611yVXSzmbeB5Wf1dn7wxUOrWZJka6iHg3JLkaBtRtiufW+z8szXi14+e+XEA84m
zGvhEOSDfgzdxo5Ltm2jirdbM5qZR0KDu4fiLrAfais7HHhkj3KZhSU+GkR1Gbg2UVbmLfVFAtl4
V4Hot4qU7JwqEf0TlQ+Mifu8hfEsXCDi7FKA6KmANEVo0uQF9TshERHorM1ooakVO4O9KSU8wgym
bt70hPGGw/wejohnrGEKrRoiq7RbxE0B9gd1iS1qqbMUOIKbB29Kw40vldHk/YPTlBwZtbs5ThOu
s8wyEdKnva6MQ2cGWEdk+eIu2hLG+twlaQizTkaBBbbA5m82bIuMWYCV4s3Dlvh4id/1gDqjFS41
7+UZ37xL6SDABvP9iqrBXp+xpNKEoxjarv5NdIZRit7YkSJ2V+xrDTxzT/Hte98xJm9vLjFm6oky
085c3+zpyGoIbawSgfufITeFKShB0fMZU1C/AzeqfF98ZbGkIsoOOPcLIDVrXmWrX7Y9DsCvgaNt
7S6jzvsjpnCtuR+mnaEXaTliqbnGd/5Rsq75h12cZhJdVH3IfMF97jNATfosbqOTz3GZYtjOoq2y
PX4hDp/hVXOqqWOZNG36vHxLz6T2tpsj5M4peFhCejjkOMjyAI/MhMit2oIjavG0EpDlQpuzD3ee
6gLWGNKSOWOp11aQoyx+GB8NY8HHxHXITZqU3WjOrwye9WZBMt9KTqTQChXWgJDelAFmgdr2OtED
RaHkfVRdL6onkvd0QusgEC4KXJi8J2qBOYnNPQcuA19wJ3Hx6p0p+zAxMlYKCJGs4fRtbR4BmfCP
rKDYX131xfAs7e/+ZovfF+TFbe0w3vFDSJA3ahxp8qcp64zh7jnEs+/nvrPYAofONFUlqqzLU9ge
+WSmA0GDRtFvgWBnqRl/D/ZDSck1U7hqRJzqf0jNMw24AKUrfsdyJZGw2xoQx3tpPTtVArVagyi2
E0wPglXNzasqh8ByXTa6vjHIuxRWh6bZMeouwdp8IBtWNYrP8GL5P9BSk7wMU6MNoTXA6G7n7AHx
Z0zWra19U5WWmiw3JHMXEZomwf1gJmZhT9cK4syWqwLepGYG6U5Zrn0xWg4aIZDoCfMJgIkbVwVv
+nY3+gJ0RAqEuQg2T7Ik264u7r3w2opGIHMidvufjjYxvl6jKjjsdYUiPjH2Di3xzz5lbUKVE3ez
OJ+GpAE6qK5b+vHi2DKrEnCM0Ih0hbvZNvaEfIT3eT+Nwr37PFvp14E8n1bS8p8zPU1UUBctwq8y
cAdmOqcZIerugPR7UPvBHGDB3kDwHDfdEU3e103qYqhOjJXRwDC+vKY12LKMQaGSbkiygfO2Al2c
W7/0q2Pa/tFAmopIHptSYeY9HRgJUruEKGZvZ1PJOvGZAWqVHkcw4r3GztqFmEsmxDH+ydjCK5Vq
KkGKAChqEzWULYaVfjXvqkhw29o5JQbmTbs8BCzy/XA9rdpDyzpE3tc77H06ZMPz8jnKRSHBC1Jb
9DAXXizQUTKdZtNxAvWC7MuyCl9FGXjEUsdVrHG6Z/yjFpoyK41RgtJc50qSkXODqwgpU6xXm7M5
y7tmI73b/LAKL/oERN+maeuyZ/bFgeZtzHo8RAB6G6SMWtO3/hs+NwA7MiesfFdGPrV4vAGpc72Z
m9E0P7boyaCyzeYItivNEzYdp7CeAjLr0VU9dVXemcDI8JeuGG6YtOWnmIszHRbx46UYGjmeFRpn
Xg5Qtw+tulDBdbUN2NK689010FduBoaYG4EWmQegYRvmZPwaCKuQ254bkJNS8vYCsf9jBMcU2qVr
Efeu/sSmQZBvHD5cpDrX7dLTWUyIQnSIWDzxQlyZLSwALZVeUwxeA8YqWnroPmWnL2/E7UiLqswy
pqRqfKT3AveGCw5vJ+8667NsKxuDmkPZlN6gu3sqbZSRjS1JyqYDiWg8urwwrzs+H4UGVP5G81AT
Sc88CDr/n80+Ox3snT3xOCU2s8WSHPkSAAeUCCT24kioXbXqxj2o8PBgzg8JzutIg33uSUK3M518
Ql/D4xwv488b32m+3nTmmTFy0IWAUFHL97aqov/qX5OdkV7HfHAAEtGsdABuuDt2IJ3OsF4BdteQ
2cCRVFP8l7mIhh4Mk2gH66NfQuvUpvJmL2TpcPNL87gLHVXYwA/i1zJ/HASWIHq2148tYo87iSFb
GgOWa8g6BgiOIZl5EP7xRP+wSGJBib3sFlEn4Nct8r6gi+OG8buhLi3Xft7ymlpMsgUCq+MipGj/
JjqV3g8H+SO07MBqchvIk0NcMXTrlOi+7ij5FI7ALgnrbgfJo09/rvMkQfZvOFQumCBo9UQH78bV
UfeSUwdjgz9pHKJPEhRAD9yraIXeMXeUEEaOrFOjQHXvWneXL14bkakbGV1NRpoYVTeqRNKCJi/f
mYGQABOxtdgjV3LF7JsAvur2HPd7M8Zex8AR85L5vVh8UBdiKtQBhzoILgKEFpeQ3rsQ/fl1IWoU
D05c/uv4nYYQYv86VqPHbILgaz5B0iN8Ewd69SCwSFhD5hwB0B5BxSO6s1jFWtSwCWTorRUdHKHF
X0C1eV+svvQfhBHY/n1ez26kzmXjWRxjK/Ow3FaI+1Z7o1WPSYjkZW3ybt7wK3A2IJJOtRh2sPIY
mYkZyuOyJzrnQ5m98J95L5Gb8+NyBCKkfgwkHDvOKsEHiJilYXCvFctPaQzchYDxm3dW/8/7Yqe3
fYXz8Phdl8drdS87MeKX5NkuqfirnuXmSwj3bq49URcJF0tSdvRHfcy9eibFjmwyBaJSYs+pUcjr
JEPY8DCy9yz8i3pxBfEYIuWiQeM9RsSWsN+aDTo1MiCkZyTAmlQe41F+JORrNqOvQLneZPH0C+g9
RGM8ehqxr0khhnJpxQrkXlT/fh4hjdOCfluPyke1ZaPfvVU3V/Hpcb66maVIZglS4TmiJqhsL0mj
h/erDbPoK/v8aQY8y8LH1/vprQE1sc3IpIBq1emmSy4CgBVMsf1752rdTZdI4AKyxJfKGgrDFHn8
/gJRCPX8DTDhUgSzQS/s1BDy8VGfz0ahWpoIiIP/n9g+49OD9s5dVJ6rZEz4kKzIX2O60o52Vnq7
f3YAXw2gYDgFmvM6rJ/wvr3FuARNg2tkYvcx3a131TSXWL++4D+6Vrl/N/puWGEMtiTDJ4G51mEv
WPvXJ/XEP9w4EASsUoMvOprfwwEVTqUNTAniQY+CZAavAW4rAHUPzFwXAQm97CLgWhZcTSW0h0b9
lkaEpaplUB6i43ldHN3sZ4d1AL0impgtN1CmOrK7Yydt7Je69lQbU7ZhqNdReCEybi0/oz5SnBuk
TssZ3iJMSImy4b9I8kl3EKD5dvjD3AJ06GFKQVRqAynN0P/P5rRmifxtfxntztR9NXYlNfyfsDfT
Ej0jqMBWV028vUn3qrg+JzrCc/z9ZssgMY4B4U1p+jiC3A+Y41axFYa+5HPFf82yiQzpW3FfYgrJ
VuZ7jci+8yyl8TFizdXOb2N5bcB6gDd9vcOOKm8yaUzJjozmHzfnMYkbM0L32TUnHciClK+RPvCV
daKB4mu8i99f3EWr+u4PteiXZLRGDq7NeX5NjRHH0VFJeoPYnnmn07Qp+HlsNpMmt+lN44t/Cf7W
DwxZb8OSoWjNrYWjmREv2pp/UZ/T7VLSreUcsLlnFkzXmX+/tcOAzFGrt5MbZwGchbsLMMQUPe7H
pJgzg8MCU/awH0XEmsGj7CLsee2yuhJ3+3RfLOBzbTIKhpeqmq56i6xdBYNMdbi04F8BYH2DNNJU
jWMGUw+npDGDOfsz2PP57mAU2/JGCVvRXesGFWXlCwHL28OY06CrM56/8EMlZspZDapeTnvN6NTw
3NmM56p5E/4FB9N70SEUnj4y13UlB867IIDeQXB+J6+RlGky87VZN0qsivuKu7VGxKwqkIXHXP6a
qJMrTzvTdAdj1QqeFsZ/JVKw9cWKxAoCeseNEKnCJIFWNvEnV5zGxD0IBWa/VH1wvkFaXHbdU0Ca
Jzh8VwPFjujlRo6yW6JvWER0turqIhKg0BrnaIFqh7GuhsykqGiOm5xvm5kT2ybHXkICs7mQbTUb
SsVWCQgBFAX1OilIDPCzVqLgppzMJvg7bDYAQaudqbykdITPDC+Wz4ILvI7vcjIWMCC/pDYeBbPt
Pv1wTVHCyRdKIUKQf5ZnKf5GCzFVNjoQAJ8dqdGJGAVM67AR3IDU2PUb4fMg2j5EdQzUR1Vs5jFN
rJ3vk7baw8rBuL0r7zqxlxPDTMkFRm37ks8e2d72H9NPav4DvmLSeFWdhrkYI94EaGOHSGtg5bGP
eVj58RAyo2hiMcfA5RvynYlGGf+rO1OzIYK/5eWtZZdaT3ieKZAr6Wwl1cdL+XXbfs11/026kpmV
ErScNc2W0WiUhpwuVKuH22h3PeU94F9ESEcZWKTGLhxe/IdG65VrwUiqFNOHN81rsngBueXXJfCX
xNO17YqeIUXhUvF7C0Ej2lxdffesT2rdiEMfscrfI6l2Z7ihWyCsY6KIqv735DdYZKGaxH+85UMD
axr1DqK8wq3SbyH7IDoDXtOFN3N2utkiaXbt+QRTxuFCL3RlTlIwEQAAIOyNWXt65y1616Pw6KCy
qjuAYo2sUG3+SB8sFMTVdZ/kDr+VODf+Hqfw7azx+QvfXb5NcWNsCeWStlyMIoMO7baCSWh7oayz
LNkuRDyQveoo/o25EG7igWH4CH0TmRMCuUHik57eMSxGxSN6xSTkkA4xGrOtE6LEB/BXUd93s33V
TauaLb0li5YSfNQTpmwVO87CyOgWOcv7WivjL4jrSzxWsxdrvY0zWpztgKE3/+GI+gJBjcE2KikQ
wh1JI6CPs0+EDfjvkxQvNpx/FHfse/dJZX5BSXO/Tz4br08zN12JN3jrQrKQTvyXmRtaz6jkGUV3
ZqopYp2xwYMpKACFqtNKWe7rv3VZAcCWzzcXCGGPlwGFE9JVrOze36WL1l9EreWOnTm0o/05i0cU
pHpEuA5RiGX92Swe6SylRaFU31lmOeVBPTYazsB0JPaKHHCz3VI8DGJV4Rhwu1LSSDnK25X1Fepu
MyPLcuM4OIm1EDP8yiO99v1G09dZGwQAhr0ah0p2LqNWEvd45YSZ3IIvUYgOAcTKSO+KZxmSwCgL
YKymVpZQ6bCn5uTL83s7wJ6zr35F/EP33VuslWc/HaPkYcThmUUPfNtgUQL+6iM+W8KEDDtj/4m0
ZJzWQKgI5vmLK/HAcVrcBhDJfgRaINscVNmPV1/qYyqf+NIv7YsBY+mWXUJFitPYocbF43ix7pDl
fQL7qxA6lkRCOZd96FM2jdsVWqMj8cbPCOsige1PUwhIzqFe3wLHOFOXmKEbN1VAf2QC2hCb0UUr
kt/kTZCNiJ26sQjiQkuwE7SQoPGv/gpvU6wmeTupy6Xteo8/ac5DTRowjCHPlxquaz1WUDryXpa6
VJpIRnnhsjZpse0c80VRF7vL+1iMI1cuDHh0NKfd7wrMW85kRuchg5uJgCS4wI58bm1Harpb7ECs
SXQM0aoBADzO96fIXqEk+ICawsT4Qt4NiScsGTyZ2pIgBULlKyPxgZ5XXcOfGTrjk/XoKdZHxgaB
KJ5tcWIK6X3RFtyjXDoVuMrAF8Q06Kc3hu8L7cK8/nGmBPwWJ+jgPXK60eQSmUZm7oIa4Y37orw6
z3/NpipOHiCHiQL7LJzCbXHOc93HQIV1xUFfF6J2e5kIRSikK3GCOx4iJbdg2c3txZ1I14g/JNkE
qH+uU78pGofFmZe0ua0e2aoUHmt+JJXY6nQCjgYQXFHqUyqUKjGA52VL1PBJXXwWT8uoAbgdYikk
OaZuyH0PbjqVXbbDo4w/iKNlykYiu52W3CvPYjpje/qbj7AK6r8nBxw/ql48A534Y5rUTxUzSzGS
YvUQY3QebcxDXXt9qaJwltm2YheqeHSwh4g6BJLkBQ7+1fJjujO2kP24a6VR4MIuyY+cxXSYsQUq
ocVxt4FImwehZ3W2PFyj5DYgxrEdPglZi8/b13wRf42y92J5xkZmFfI3lxImBt2xbXeOyz2ctfGg
676Xb3U3/RAy/ZZL5fzShFAr8Cd2XPsLlaAmyLf/VpEIJM05uVPBVZ7bORRYCQHBg6o3MbQP603G
P6oIzzQrS+lJc/8ls/H/ome7Hmtipy8Z8ITrqjiGaZzbxpbdLCLp3dQVO7BoyZudS6ExKC4JtmSm
HjQpWu+6nb7GMjWouIsXch4Vfb5VsFwRh5tW6vW7J675FsK+mPIfRPJnIQ6/6nt3/LNKJ5/aqjTd
/ZP8lSxjBcBGQeSPRpaSkFllN77vLXbnZcbSRhtboJVpjgY6Hw2uel5u1SWByjKFh/JTOaNWIBYY
bdziNVo4ekgLg9dNyjSZtvfiq912a4+uAGByfk4VanrM27uURW5FNtbCJ7C3Azb6w85ZWmHou1js
8zx7YDOCDG2vtGiFszL7XMWlHT+Da0lYF1uUSXp1mzMFgogoxWP/MBQkMaMK/SEoiWd9Q1RtZw19
cq0hq0yar17CVWELg7dGwSXv+RSbHk61hEGVPwFKv6kK2x5h73WRiWYq6nuypFAqtcbcQpXVKRQY
ZAYp667MYIkCUBtzq7nA1ju5PU89QKYEctAramgOT94Ty+t9VLpKbSm6hWCSDw1as3gEmTqpSyam
mBZC3nVc683uawePoRxuCNuQc0+d3bc7xwjHHuVQHG8dD3tKKE5fRHRYzVRxrU1HxhvTf0JITc3Q
6PvKCF9fTR+IBA9OpJKyU1eLqXg/vHlqLORJSR3UCndMf/IO7zQzYhE2xoYOyY1CIyeYkwgiOzan
OQvD5RPeFTrRJ03SBlVPtDiaE11ovE2ZT7ca+YJuzztdKFWSoYU0M3sjuFvir9RXCrgJCabY83ea
9mu4N2TQ/CFsO85yMEmghBX+oQxnro9wp7ZOzXfSBdk6lso1QGo15bP2z/bWtjVSZryv4mD6PwI1
XhMVUyZjlcGh3cq+1A8bRf1jgvoQlfObSb0TQagyirRGxoAX6FpEr+CX64wIEEn0ugK28nzJAFL2
uv0vUHeSTFXlDUwetMdww76vcNuLI6CULu9tA3x/GnhHdC9ucPO6t1ZHZ77OK3RpRdXsMOOEU2WK
rhrCiRroMpnpYKEsiIfnwZV2LXE4OiXI/Jsm47tH3KUrPg1vBsfDIsq3IX2Mf7rGug20fxqKrIyj
wK5d9F255Y/YSKvBlv5nzENHo4ZegODcq5MfRN6z+HTxi5zFRl+T6ykwgX9PGBtBepk2HfrwrA/0
5FT3Um3pgVCzsdolzGKhhwn6MUuwUkGgvw3HuRTJGef9DGuc0YvPaoZngSbc4dPv+oW9oOv2OrSN
dRPhZt7+uxrqr6dsxFlbe8jJ2JraBZxMscmaMZ3u/OVz3FOB7+5ToIks6pukCbgvpU9QlpgJAq5Y
I4VzjNogXjKHAmO9uIjWHAmLkCaRz7kE3vHiWDeiu6WmRNu8sS0wqTek90ILIpljtw5co5U5mbM7
33g/wRy17XrpNCWdXGsik7UDMotVGt1fYtHido/eGAXBxNoS/lZRxfA/rVJ0wc/NHWEWi8P5hJ8d
Q+OzoXKA72GCMunkZvaSNhvdPx8HoC538sM1BNO7EfOiROwHe8UWS7sytvB/l1d9BXafTUaSfL/b
1czlu6aZEwVFq7PhYlZ7HibEgKuFYtwJ8RudrQieodwRevgIb8IyQW7vDu/o71AR2OuSnyPcE+Lr
uV7PoDXh1/80AgD22INcwmXoW1dz0WqWB3O8cb8pUcBQMnWRXrzF2O0n/hca9pUdpNJ74lF2NpHA
nKZTe9k7ohn7OEbwMRFAff+SVwJfIFsOBApE/BCLqGIkaJv/cR4+4+cJD2vV5nlZiSd+GEErRET5
kQ1oR8FXuNnMuk1NohVIzrzcmnepkVmCxZPv3TZIuHVx5WMalF9+v3XNwcgo09n1T+1vsPPFo59Z
a68Ye++JEjXKEys0LSr7YKcdWTjC/wUvyKivMWb7dq3pIC0g/uZrKc6dtLg3BWnqcce7cH7I1TQ4
0hMcirz4KCLLovQnlviDB3/+avgqlrDGylJI6xsdzjdtOwEepe5NlauFIPX61FefzHWHu/lVwxxV
LxkG2zBorISHJ4tjMcTea0eeYFiY74RmasUe0efreLoGR33qcN5AO0jYart72Ak6AgwkSHtIcY9h
0SnoXulD+WLlzD7RxXu2yjMm4GInxxD5VuRhKOHaytaMNsopiyNnGVKg2rwrZbCAfoNgPJfSkMIX
yUBPkJijTs58YxmR04OFqfOpOH6XLi8oAIQ9Ei2Q+u66rAdT56GRHhyfMNsq7mNs9uYb1wDbIeJn
ywpzaES9bWUVYfQgeLR761vrVhzbAXY+9MB/Hkv4XInjs/pzB3N9Kjb/ETt3cLd37n2aC8w8yeAk
/gm5D882r3ZTcABbajyCXEw8QVXhaPE3JJBjSdv5KkSVZmM8ZqFvIzjB92tQedvg1IJ9SKt4ZPk+
qWz6eNm5ijzRX0P3o928iUNJkjWINp9rIGBi1Mv1swC+CMABfkfUwpbNxpmOUag9lWlN5UnJ1Ztn
aTSkwb0AoaV93aadqxD0Ym8wmgkBp3qoAOFMmEqQ64bqeV13rS0BNpC3oDsOyyQmjYaQeJWGFTZ5
IiSBCzBbcv2HbLSUmcZRmqEb4G2bO8sTx3OZJZQ4YbBZTdzSw+iYkU/J1mZFG1dc0ldmhi9Inmln
7BCxFh+uV+ywrAZ8SAbgvHXXWHL7TPbeHe/GEqdW8C40i9DMAh64QC80cy9yV3VTBfF9NptwISKY
FUz5MPNAh8PKUf4+4fT4x2QCKE6KM/ZnemAkL9/FUG38KQJ81N0ZtPgOuDBxipnsalOGWoeGwqT/
6uLBo1iZD4oEbyxHEbG/nWel3Uf19ZDqzojWCI++x+xW7ggtrUe8y3sk1Wmt9WCwVhEXkdot4hHK
T/De3NRHJ2/lowyqL/JD+sgWgNOwSJphGnKqP5TKdvKkyCSeIgbhA04IleHkyhPP4JPLqxgMd1x1
bllMWZ9QISjnKhIHl5ooR7OuwAzF8T++9uyJLQmd+HWXd2IFFHjU4lQZ3091ZHMPzssjCrtlRlfW
WkOBAAmSVUf8ngrOnFmrOrqo5TXRDaNCiagkZFErr4VES6D9rL871PQrm2W2uYtAb5OlPml15hGT
BTsItnMDPBr9+Dvomtha9Fgqo/t9BtF9re5Tkwk8ARi810VeUiaZ7G+nSSE6sMhQD2cRs5brWm/h
ftRWKcHJlFxosoTcWZUQ9II1BGc1sUbLF6bgrG6W6zs+vYox0bDfIjE/NIeTnUn3hZdQAmCIRE0P
t3BOKCgT2yi3nV9TfFRcIYGV/sXGy3cnOVTM3Z3SopqGvp/yA8cuFQm68OaQONZzAgWLAa6+++tf
hKiu0wTyxotN3lCltbNm8OL5h/F+dbTYTjYdnLtBItEXv451F9jc310/bC2l0Xp9DpP5fmi+3tJO
QlutFfBHoV5u6ELe5EOKRfGkahoO/7QmMUX7t26BvLmY7tCfmKFkmv+Q5nWLk3cVJsdDd3EaopWK
//se4zzI8uz0NBUCQJk8cQWYPAlzFW7+G1G/1Y2lPQ75d+lUUCY9tKkGU/zn3RmSRNr4aLqrJrDF
MSgSXbNYQvi4h5naqk/SI8v2jh7PuKaELAqRQhdsO/izAzGxLznIsBhnV0L9NaJ5iUSk+Vbi+GtY
52FMXesfTh+sw0ZHvJ/2Jk9CNJ5DHlz8wBqaKdNiVtjooLrEvqCxy2ioL0NkZPV/QrxnPLWnAVCm
Zb4KsJ6TWBeMEh4aTDjKMcHF3QWjbW2iTRpOdrA6j52pd/H+H3BRPQ2zblMA74seF0WZEnnNgFwF
eaHgXo7FtZKaSCjhgAkoQJoLZTxbQdLUmuET9gGFjc1E/KafBPkzhyZdDW+ZPaVg2XcVeECl5ve6
HYB1pCKHTGmLA20x4Igei4kwgH/XR/PhzkAaoHkcoILIWOxrChFN6/q1ovkRggB8RUqAvsnGQ0EK
7TAyD8e7qlRZCJZ401nw5pypuo/AwRg0JFUU4RRqIL349YfJzoTTp01cXE1vWKXRk4qcqfKhqWtQ
fjbszAIT5WyPwyb+izcU/CqkJZKvQ88Cry6s3eN9gUIQW34MtWs1dW66NouBOV8atG1AbIBPlPug
hGAziMSJ1Qtb+O6g9zqsYAoCuvgtTGceJ/aQ2zPtpnn+f2xfzGBVTq11CaGxkSw+E1cpDR0LV0Sg
HtEV+f9s3Z3Sc3oYxQNVEFbIzUAmIgz/buwJQFKBjRst6+6KpHgvB/JZdbhlnEwB2vud57tUyIsB
onDL26wSMe7GgGK9DzH3DW/r+2IWBHYFwVUKxdysgoE7kwtX+DzAhkSTC1xdTq2oUri08cPHKfQf
yut4GuMS1oxPp+PDejH+Ooz3QnKr4vQd4LiIj0mi+6rRrkvotl8/AJ74b3j69GCyZJF7Pr5KcelT
k91fiMXB28a6hD3jASFCf5nB0YlSzwzdknkyqNtY+LQsg6yjgdGcSLenk6sw8mfX+oy1OZPf4ldB
PgAn0I2PA5PPJChOxoWbqsGXikokqOhSDyyfxDvYCf9ab/qyPnEjU1gSLM5XRDeUXdj8tRqvOYT0
hUQDcuoT0JD/93ufp7dMrWnWVtdkT+tyHv0L77b2n6WWsjQYFasMsx630x+jsZEcsWLBmgC6SBtK
elOcihhI+CA6qv27Zb3EumVpdPvS5ogK9tnMy+gGJE3Bj8XtFa53xbrvHSt7dcxlooOsDpDlGbem
VxrASaojcJpDfGf8ueMTr/GlWiFSLJbZ1YitbhUxLYgQMkiX/INJ+5nf2ffIMpHxqd9yo4/+2pxa
FR0TEpX7SFd8qm4SkLhveUpWVTZswuBbnH3r+mngTkG6w61jU8ktl12AxRrurp2+9eFitKMvTXAX
aOl0kp6YOZGH/cUMTNMTkEmnIZ7EmKdX91ILUXBE1lQmaB6HHqom7rm8ZFU8lfVGk5ALdhXion/N
z+Tu5Xk9xUrDgwOdyGnqrAlyHnavlq+8FVXGGrLnQa6gpqCiDpvI8ja6hBriS2A+mPWZ4MXOUR80
aaSmX+c9OP438I81yowXgxiHOZANRr9d00PXyVQhKy5bTN0tw49UNGEB7vW2FxMLDHHjmh3E3+M7
FqimWZfdemz6A4jSAcYcwI0KM1pGYqIFCoiyNeODstvwLJuupJti1uKO4r1IbCtidmy7BlAuHJsU
fj6m8BLTZjWNTEjnXX++sC52sFu7SNJc6nkiylHhlXpAtDo1ulsJmo+xWhoPpSBr6H3iXjxrSR91
ZI9GUE9TUPCvQs0W1kR6izvuKcRLyhxyXZGnNrh+XQXSWjBo4DnUDrnfwsSQQOuzmltNke3JHtMh
aWumBmcubLJlqhCvfJMymR0CohnDxEXC/BSchzuYatJHTu8O51tgJHgn2t4L/yUm0OC6T1W6q3AK
2rRQdFqeSpxspwrjaxaPZR4z3SnG13TtjOe1BmEX4dWAZzNmARC6UFZDSdFEqNQ9Y3kVphhXkP2J
r8VUw3+bZ+Ect10mOUG1k0PNosM2TTJO9gEuxhkIuW1ZU5b3XzdKfWWEpYYfk3dj3tm3KWRj0qdP
s43M0AiEDGpLzomWgjROzZfMYhAUpDdcV8W/ajfTxcOd50EjTidIauxyb84+F112sCxJJM9NcotZ
JEIZYXu6Z329k7PkwgLG4XjRTzo/U4bQ75GBmdJ3JYX9OikAWb1DRn6GyO17XcqtfUjdxjNWPr5n
DXipmpJeJRPrmadekdCtBnzkMWqYl3FIyomb0XNe19jeZyxcBpZZyw98AENGhocZzMpc5GiFJ60G
3vF0SNaHkt/S3Dz8TCH0BvD5px5AEn/El/SJt3IRHY8AsAG7t0sTMYRw5Azj3Vz/vHF2L+0rETeJ
V5WNEzEgHQdJiiI1wBoFjZjhfy54lYAN/K8MX9cspubFH0VH6BbbLp7yCQrPl8m7ZA95sMWXoj2c
62+81dPkWNu6m6rVeRyTdkpgaVsmejtcEnSDKEoitt9QuN9yJCRzfC3hI20BT/znETqDSMNJfk9K
3RI7qA3iMCOc02DWgcRC3FwuAQbMASN3CfiTDmmqcPI53URk0e6Cst9pLOtMdU2pKqhCV8jvcf2r
kHo4l9z1mvae0S7A6+pqjsk+egsEPOCXwSkptaVam7Wyqm4AL3ktXohQgEVXcnEbHAHF0VYxwotx
AYNmhLY3bBHsdoA39Da++Gfx08CCrN7hQyvv+rVZJ87I9LrHk3Xsy1r/q1eFDKFLPqpvW3mO+8ST
As/LI/BboC95me+ywNbgsQ+7pM0iGzXhU60xt9qMUwPTEz5PB0fpXDHKbkTjkM6xjCNTqU//BWYn
p35+Ja6USzK9YODMgqbaN6aePKRqtyj7FduLzXpsLxWTnpvSTxOUMGdbciSaYZAWwCKYVCO20mcZ
jYjsTtiZPiNtUOZ5aoSDMORWkVyWb1nwGnLO73ij6lEqXJNcKCDCp2SSnd804TpefL5dPKi5zTRy
J8S51JE3hoYKNUC/7mzi7nR4yWe2QKdZt0HO1NHspDG6m7mouDzzYIn/nWpGf7wRSihiiK80fMN0
e36Q++24Aw5bMRno0yR26Q2phvsR5Dk9Pw66vJbf7EzJQbL7yKD76JYmGEO0yRO79Dk7BgLsyoIs
nWLmOyfXJLWGvLDCS+ATRYGddtZjEwDWz/sePsNUNTyrDlNb7fJBxaDGlKsbZS7NxTQyNrIsF/Hi
Enmd6oZimcaNWdWRutjr0nh7WYV63C7VhQXRXg/JYBWpTgjLk4PF/1KzwVB0pJswuAu+5cp2uRZU
G/oDe05tluYjqQQJCh8Qj8ARNRICotFSqTJ5HKotkI8Cu7MnzyMsVLOVDFFwqHaVuh3P2+HAqDxM
+tmE8kC/nKQ/pcnhABjNCJvJ9vCm1T2S9lZPH2kP87iapj5kcCVHc0a7VswqMIjCSPtbTvIpS2S5
yuNIrkwoiwns/CP4H6Lf8zwf4lRqwic0Uj8WIHM9sFmqkDD6wRj2nZ7m5mLQGjtlN3ZsXRhj/+b+
RGQ84diXtFD0aQ49bvjgPMk2vAEFETQfqzXKbiY14o0xEXfVOAfbL4XS2rS0z6KWQPxWPmErO+C/
OYNozLTSghOU8ovEkc4FIYCZk6+mQE0zsMPHORuOESqtBrNtXyL+SA6yWEwIdOvd+QS/heKZROmC
8FJliT5ZwqfGmSBxzV40RhCys3eg0ZTb9rxjtE2V6R7LqDfkVkcoNR0u4Kg+uNkJtIntqMyG5fbK
rvN32jmMoKGlwpjTdsKxzgC+QEz4GXzLUyhEF/HzqgchYRTjPf8+N4S8SiMVzJdnFF4gvIKUeyQq
Em6pJctfdrPcBeMZnZxjvKbBXXQQLbj6sBtTS6zgULm/6zJjBzpnTBKNJaahjX9RY5qhkoc2hdbG
1tz9CpXFoBHAd3Z1BOhw3GI6uJ6mZgwXkh3MIpwGFfA4vG6Y2n5ju6REPDSk3GuF849NR69yAmxE
DQ5IThSQmGbiFPrF/evU8+RDvR++QCZH0kQ/dXICbpIe6lutbFUZgYZffJfiSIG9JDKvaTW14QEo
3G0VhkAIuw3ApbOESDptIXOP9yBAKhxjA6t2DAzXDnUUN5YeWm6biO7omn5WwmCFNM5DhVBdRqR9
Ejq3H4TkpnikJloQgn7mnfIfvoBzE5jIu7p/34ekma5MqeUJwjXzYXEeQxyI+bQrndwZZsLIYrAg
vKBrqHp/TJkW9vG3plySsoSdKSr/chwzGOvMMvpSbIpVeR8Ts0K+ajebHFFcUoNPHEcJnLekxRv7
l0s0oVXj3C/E/WGMiy8ks86YzyANLRsVP547lgP9E28XVrt1+wMdNvnlyRlftwh3wdv8dpzAi8TJ
CCHgCY787pXkEypmqsiINEQHJsOYQnCECNpKWsIOnVTih1vpNRG8V71v/jSyJa+jQd7538cpkgIS
RLiXU64LoP2MzWaghLTHqtJj9uwN5PQuHsNiV9/66wyrIrTTAmeS2jJqlnXI5sszBC420cp+Ebh3
GFHVzlkJ+Iz1+tfvpbRyOgQwo3xX2qWM+hXegVvwTrSeIK9uYk9SzbyL2VY0kfQL+IjwKEw6jaXD
/+ItHWrwrNeH/3r9jtz/cYi+flpdWQKSQgywmxZ5SlZfaKm6Q0F7YzvOiKoENFwmj8W81FG0tc94
crLhd11pFAYQepQJ5KcRDsUwYMBLgu/ES4g1dnvx30UZa9rWpH9Q1zNE3j4tYtP/ws6yFFcD36jT
4C7qMaHaHnS+KRDU3bXL79ZY84HUZCoQ3dWTngoqkhW74HKeOFNPtT3Efh8LMGwAbF7c9GlxNmAX
yQ1lDRAjScdSFPvHqEhqADlNUox4V7eqqAODw1JT/hOiMnjKsDerNnjZNHbMXq4TnHzwbffNGtnO
aUtBT5TL0+0tm6kdXkYXmgYKwrRsvF5MJD77vhgmxsWdh//KH00pKy3h3HdMcQiMk3qvZ0TALnmw
7qXB7JALzZkRjkSQeTDW3gcR1Sq0i9S7GWJniND+fh2DobbuDiaIQXrOb4E/uIvgyAH3Qn5km5wB
/3Q4yrxgT/amhgLF6xoalaLpEEiAWZvFdhEbPrtCSPd28G0XSgJzwspsD/C5U/RZB3D1hJTHOz4/
lLdrLtSmHFVw1CR7NgvuZ5MpP4lUNdiuR0xR2lGvG6Z+rLb97viXXI0RJ2H0I2R9aH85HiKCmSP7
Q07QM4WWamDI8fggRx1lBvtvsEcEeXxlZmi39opvMdew74VfoPaDCj1pcMtIh3bPqYrRAo77jzAP
WN8AHdsJHBFwSjeihDE830+NM+gNk2JJZZ9UJRblbJJ7xhVqSzJ35y2P7HXQuETJDiMjHUy2T9Uq
O+LFpjsiZM6IyP3J61mizvqTjvFTvCqBzxhIPPMV6WkwcMNPGonKAxtPIYSOBAcZSNSadJIc3VSc
XmiTV7I1GLGbZSu9u5+XPVvWTJWBgtIMlCyAmOuzhpKt9u8YaBWiQ3dAcKytOYpMajGF/GX91IDZ
RpTWSPiWz7FlkrKkO2d9bbfEIhyyqqzvTEEVFY9ZncGYWeivQYhRgA4lt6/pXk+SUD7BFDlMYuU6
9x07BmvdAUVfMqGrHYXeH9GlO3oZbOh1KrMrX9EkzlS4Vkr4r2ot7TmbgNuXuZ+65+/C9xYGMpzI
HxExI03g3vDQ54g8BexKciaLodPbVGMcEY3vecGTzGfJSgnH2wXTyVaEnlYsS1a51/AZzjdOgQNj
mxBVr0+yXM+K91w861WjmiIM1ydQym303xZbkspsUhI1MLysrt3nQL49dnCwABZwD4mAIHND6t7J
BCVwyaEwPs2RXhJYFSrqscaK46JGIDC5uOceDzfLynW6ItKjG5UxRM5lBVUqgrDUeaz6b3IEt+rq
7KmkTrJkzZervV0ATnKBmcBdPMSqbOdB9H6IWANndbEywepWvOziByFulHdG2uSSiKYnIM/AmgMA
wEuFrxlhOASrtO5iJgaVXDfSwtUr0Ad54CPg1xzEFLUgoi80pAu3uX1stENzmKf6/EjTxPgWP+Tm
XVFdApkHlGMgHlXAwO6LMBsOiud0Yp4l2HSBniGDfv3Ae89Fknfai/ykiF5Gkuv3VF3C98hf0cIx
dFzprgJs8Oyi8ta5JjsyuFVM5JM3Gr39gJIP9CNb8RTnJK3Y5fEt8C/R84gtx3RqFZLO0zyTs1ic
+tDnKCljx0snmOo9hS9rfCO49kBQpbuIjFTOGKAag1LHdCMBDeT4tMJMSx4xl5EheooT8HkGwnTg
WdnLtlChyNrgcV79ZGNxihHMnZakIXQOa2r1F+fvNjRYdc8D7Pu94q9SIZEnESrwlQdgc9uilC9A
oD4QNmAbeq0NyVzhTSUeo3W1vl6win106c3joShZrgUtJsZvXBoztO3XWMrIwzyHKu73VumD2AVG
URCon9JLYj8d8aJrYznKoJcVlaAWS2lzZ1mAC4/7SGwV/GDgdqOGiIkeWv26HyVtAN82/57YCTZj
UPjuOXA/CEkhplbg6jmtmh5VNNV1hvxwggcSyKjl6QdjfW85iQLabEkfthjn4Z0LnwGVmrqHMklc
ShYD7sqq1Bwri8mzDU5cdRhf8NrOtgCiAeeK2eaTeiWaGA/dV82/ULEPDu+AuRmsuqVNQ+wnAKnS
BDJYA502J/E+3xOHv9eLaGCnI/X3LLyPBm8a8n0qJLW1Mzo6u43apZOIjxSMjU0JL7LnEtpLDHI7
ILXTq5pj7vzHhQBWJav9PYa+HSuiLQHeNq+9jyzg9z6TqlBlBksN2+4IAfayTPRBGWyjnT2DD+O5
QB+ugVQXrm6HzDoG+mmjhiFSDNk8xuZfXI3UGaBiCUJrPcjSxPl0tOJibrreZZ1TX5zozJJ+yr62
M4phK0AVU3qMPkapDI5jm0X1gYjbRd4yJuO5bek11U6kRrMpvwWZsN+xuStT1h/Jfg3F4tfgy/3t
mjq4U0W13JghoKxFjOdkp5LNwDv6/KaqjeqSxuJUrW8+ls2JHOBtO617sV/0FU6OAsYsPwzF89JA
sK4k2SZIG8fRBVWZjcE/hxcIcqe4WB9n3eq/E0ue/t7oe+8ytqeM81Q3N1Yhsy5c8sO9McEB75zu
WYczzD0B+i4+a8ap+d6aCch41UPNe2XZRBpBlD+vF7Xogj/vAT9Noysp+xjGEfNeL8SiDqZd5nlV
9vGIPQojgFLkVt/H22PR1E8qGFqVSyTSUyGogBxggRqzhSJrfRCkoHpCVgbDMNMkV4qVXSGYGg0Z
SS5StPG21DWupp+MHj7U5NcBuiVSsPoegx8SuQCrFK1oFHM3eERAs44iCsGArXsCyxW3AfmimupB
1XlD3iqvrceYtusRWDEwQdbAYUpHftkm/2seW0pcgTIRyBQEewJMi6Lw5pk9rHVToQMVJ5GEzzD2
ekIOor4HdIdirMI7RS2HLWbOFb0VlgSJGNxRaJCTBJFItWwW2SpBXBncOzTHs7lzA4O9Fxib1qfk
f2tycLr+dPx/0ca4R/hKgHhhB+tEfD078S0zhbMsfCQbWVLUqTCEy6v+wOxi0bdoYS0WVT3iVaja
onYI93Gdfcq2vszNHzfbGN2yqA7v6dCrflZxHE0aaSq1/hHfWD6mzqPLy1cDFxwz7tZXc5XNTCTq
x6OWFXrzR4HHlUIwGmVd3QRKl2aJf0AhlftTOUXh/OSthrqGyDCExFpmni7sjxC/tDGMhgfIzDZ3
suhBXpzIaI9ReRmbGx3rUr+czOtZjsmomsUdeINnB4eVEJLm7iZDv/SeWS0rkETis5BtqSMHxWDk
m4eN1Pnu9w4B132LNQmL8VM7g93zD2K6PirEhf4s9KNkfihRcffD+tDTGufj9w3/c5yrCgDczofy
2FUDpfq+EJropKNGy1pEN+mcvLgVUWSkwaSzr3yMq1PKTF6rCT1IL/7AyccfsOGgXVkLUOrZmxf7
hlzcdArb+QAK42gBj74fyEdNS3KqETwj7qYuF1x8DdNlolOasoIU44uq3qcWFCLxuFWNH65YqKhs
eKYQYNLx14f3sN1uhuCac6ShPu5KQagPwTQkUis9K3EmvfDh8m+w90MbQVYgYh7rXy3GBkjoQBAv
pk5FSOp4Z54Do3vzTNriZ53ijp57+Zkiz5uli/AXymVA61jRqboY3sYUcOOCv2ZglXLp5Ruu4tcC
noY5lp01H52Kii3HoAfg/dYj+5JzcK2+LhOvyYspmcgsO63WHCqzYzPjMJLlHsyHbmfmLrFebLNm
EtrR9sfPfuQiuRSmp6inrx0WFUFh93fQC6SEdhTl0NSua/A7cRHvkwoN2TE9696B/vnKPAiXSst9
YOhrHEJz18aJlHuI9pbJ0lGBZNSn4YRTvWe9+aWbwk1OBCNq97YNZdS8NgH2XHVQogTdxmdk1v/v
cpht3dYsIVIwVJcCoajV9mfDx2+lMyu9ygHSrQlxpjY8NNPHvw4pvFa/K+/38QYVb38lJR4buCN1
SdN+tGBHX/AJSc+ZDRszjo9gYEKklv8t+e6DQpwEUySCMGCMyAtSF2FFnnR9TX/aowd98zde0xqm
yD/q7pI1uyX1hY2D5JSytvk3/3kpoe0OLFeGBFD3qFOO4LFIAHhGw9oS/azydwXYHUf3m1AeWlM3
uh/dHp8ltMbtuyR0uLaKqT1TRCHps+WNxv1w85HS/4sXXMB6TYRIYWWaDaAqgIJSsVjWbxrzjZqZ
VeRAP7kZCYUhXqoPC+K1zrB1ZEXlnOf0jluoTQL6W8jt+0tUUB907piT40Hs7Ct0RgvnorweSRsM
lFbQIJQ1wQuPfDpAh2wMq5SSgiRWKaSy9MM5EVEjDRQ6Xttikh8GqiwpwMqe4ffX2ZKogDNOzGBW
iLNYM+hA0epokrd1OUFGdT3VZ4Cd96Rmg+TemwKZp8cj8gISVR1gbjAbTKJN+V/49f2fZId7cOLt
o8l7nhCoBUzRzD2PlSbREeZt+p/PdcrNETij9LEKD0az9BPhVElQP12+yY/C4PfOUQo+NLh0Cy3e
yDvn3eqxl5BY7JaA2FXPXQSuzF94PTPoDrkx5lI8F+lLz8MeZ7EflTj5GQNb3ayITlaAweOCJrzM
6syU0cKn0jZXeiphCeDBolNSI5KIdE63PbjTK9YN/Y1DNpLJ3u8NyFHyxEpG5MkT7A0f+MBJvUDl
nPiLeellFd8Boek4fEG/EkNnyckUvbGtFhlpJAGQPF50XoSrYdzImtGbXKYxtm5BR7pc5I5po1Fi
7RVgzFm+PSrkpaIe72DaMJ+VM5YOzWDvoQCburEU2PYJgg9FvbT8f6c3Fnq8j5oVMTfCEPhoGu6W
4bLobwaS/NiL2VfsJ+58jnEk+pUnor2jVn4d/CVLkbpX8rO8INqAjpBooq/9qI+9OsAt/lruk+kJ
WAz+3F2sMqlPHfOIYfmWpMwaYcxRpEeBvzi/Py72RpVi/V4iq0cVHVpqD6Z7+UECKr/B/sxyck9Q
iLedznQ6axZ7B4HJM4+5D4jmQX8sFcRw37cJGFEKayl3Fu7PTl3ySBW0Meh1Njat7sK6msmECseX
W8KOMzc4oyfCR2wB6u+BREA6zBb0DE/8A6vEEtNjsl+GOochbnAeksKySqL3yCieA0yqi/ZarOyb
4/bQ7l0/ALiUIV3yP4YgJkAZqplEZSD/c1hwjhHi6KDReNzTPHWvV//BJXiGuU3VJf98khaRTZ8G
dfOjJIKehfOPiwB0FCx6P2LJkty3r8YeSgNrKNYY39jIQ/+h7sx+5j56h7KJKvTVtjuNPLhW/svN
iIphW9IoY9x0OSnPvIUzLpcAbtxadPztemy0p+pksUlJfhngIK/HfSy5hanYNCZtOhgtkA4KmwlY
mnfSB+1VLmL3oRPE6lb4W/y/SUnrC7rkj9Iu2krqTyXDYibCH72K/57vz+8L4exUe3wsSNQgsTlb
VzS/1SmTiC1LwRvJYsTA40HtUZ1eUuDQAi9rI4RaUARTGIrbynzTFzUNVF6VbkCZ3hKnBhEJg3NY
zfdPcqckQEiEHRjPQxpOsY3u5PcpJ1TO0Mq8caq1q0bCzWDtMW01x7z2w1sXPK6zpiO0x6kjW1n2
AvpD23jxkOUtT6QWaMlMmcaGQOeJjY6lydonSDeriQam11fRQ7wNhMvP1f+aPFpOZffJ34L2pm14
eDG1BC9PxXpKGlPc3DCDg7U0x7Ehw1wvk1PMuY1TTP2acGj5N/g2FFxfDGU6XpaVPQ8Os1poisj/
FglEUauSyFbXr3uvBi7/Bf1O4q/99YkgfEk5H6sR1As1y2gfUx7EJen6t5GWVWR/xFITYaAQcs69
ryerGc1M+r+hEDZvyeOd6Gax2VE4BlkXXvgdM5Z3EksmW7SFCivtm6wsnHCQUqa2FV7eYwtZVkrE
yq8gaTVLTFWuEMiNSNtGdHsEE4s/hRD0RewGdjfN8Sj5xoaoUiwxhTuU6nPhOwmvJkldCAYed4NB
x7of2kvYHI/oIubVA/JLATw4ySSf6mHxvpud/vhTKCnRHu6c74h7XWvo7KWpiiLaH6w3sJrNualL
Z4O2ZTEo7PxdbhrFmTmwV1iuNxOIj0o2fz4+oKgKJSpQfp2hKs1D0xa3J7U3utkJw1fecY0qxa4t
cZUdGm1zciByH0xM5bK4qBTWqAm/X3H2/6RfE0nheUyclEfh1ytE3TC5rnq/Gnjkn4KQZ6s6hMuW
rZnazPSUpQsV8IX03GxulZAsMjiXkeXSjyM2sFlDod1eRKj3Qm1KdNNRrna/LfVpNg2+PsjMon/t
FXSArJWJ5s9Pslt5VW8M4cPRI5Ky8XoU6+E2QgXjCvHZw62x+3qpGDb+fdiajfe+ZAAdaa8PDsvg
JMLAzJ2GAv2ST39J10kWwrW4+naQ1Y827eOoDJobfU02IIu/N9tNrEJtUPoxTFFEQPD0Y4SpT7EY
USo9HW8N2tkRzXgSrmBVCLQL/pc5++Da9ZewL4DEQ6WloLqFY8zKy+ClqnvkrJa3GiKUtC2N5/Kc
10HWLPyXFz+1LUjZof6nkMXyAe3j26St8XrJq+L8NOyNitJvUAP6Ip1JyEP1f0cR/hlbXTfaQZyP
oZr9Y38ayN81e3kKdxuo2vtsaJPnJ9yxgtCZ9HZ9WC3FcJKXcZ2VqFOnmYjgO84l7MZ7hHi3jh+D
DKJy+lhiys/mmI+x9vl0lvPLVLsbhgWKJg3i0tE2n9l5V50k4ZQkBYGRywkTxIzfkURZwwQM+x4H
EApc10kc4YTvdgJulto5AQMOJ0N0o+hw5Wm8WCJBxRhA0CCiGSKmBAdq5y82izB+HFuyTXnjAjR7
G4zTXztwVhUFWWo4OZ5SKY8rDvaoKcWXgcgIWi9srkAbaA4GPEfoM+TgwKFUwOerTRNcRAWf05EC
yDlimnr4JzN6sltH44LDXJmA3gJFpJvN2HMS9AP/QyISwrYkwTHI0j3wIskbqBfiYb2T+nO/uiNp
s1JmHTe9O62xxeqt0x9EWGGk3WCBrf/diY9fKt93cXyNP1/RmKhDZ/eXcqlCFj5xHJrRuecbe485
mTpu9dBIfelz8tXz9vdIH5emz4VwEz2ItJl4x8pwPX4aBGp+N9rL/3u5OO6CVHPQFhUVWPihBH7V
CcHU0Ml8Q4EEedfSj5j2AHwcsLwcqx1J0hWayLiprRnnd8Gc3xWOpuI2OJRoIkhNube4vKVV8xW0
aathsy7AIr3vIfARXxrlFL49ivAMLTKBYmc7m9CJZThd9J+v9na0DPtSE565fYPt0oxMZ0A+pyii
g9FfHWKoCLG1MO+7CFvdLSMwLYWUYEar962TTiWdBSKzEeF0abztNp1umFJENlwYuyQv9cLF0Fd1
malJSsD/8G0ZYvffKid/qAfK0MoGyRSN19sKra3/B+2hhDZ8ywxhVMXAIXpctJEZKgw2Y2g0lZE3
sIXQJSMqz25pxZhibPkzS3gaVpaWDCJV8RybR8DJcAhckKpJbdUJtVusVHJsjITkejz7f9CWXgLH
xT8eWo9Vlk3kxRV2PYMwP1fCoRXii8cfCiox1h7Hx4oVz3vPfBMwRmhT3z8/g4dXsItTJD0vg1ey
jyjOZhMRUhMXmbWV2McUoOBX21hapXXfsoUFDJ+txsbo7/dYxV23vzBtHCLjpLiOWX3lhriZD4Vo
6374BSuibQ/kotc8raViiiyw0rjQ+vZWS9/ZzYQuXXimsDtPOywWOMWWYOtUahlmtHODtIeRoN/L
5dHWgqSmzmuRtNUgn95daCUwSx2ovodSrxEonTyb7TMkBVKVYtNjTM9dtFR9wMiuXLRB9oz7nFtb
gEKV0LANXn0u+bcPtFmgTgYX3C9ZuQyQESEhrUmPrq55UgoYlulJi9rEnzhED0cLxy35ODwvdGoh
BAEQW/hwJfXZ5+EnDSgw8h7Gj1dv9KOgK+mRHBlNCToF+g4qfCmY76pyWxPZQI9veB5gDkvKpCaT
zzeH3O6kC9jNW8m8JCW6tmdQ0OVkpDApccOA3JxTHFhEwUkZqywLccYUaGD/AKrpoqRBvph6hZMa
LiceYb4t2W2BxD3KTKWWjvbup5Gb+ZOsTEh3RNhtJwhOiroXzpFTkr5NR6afeNC3dhsqL48VkDWq
yXbZE2WkrP+hh6B2Vhob/h4LboH1jhymPJt6zunOY4EhnHCW5K+3kU9FN9E023HQlXlQ3T3fqco6
0Mxt+MEpt/EnfS7oXiE0FZGX5Uv33ivnXaLn3judmfvigVz0qH4QiFfuYO7DChDrMC972e8KZ/Ox
ZMhjWJPqIpuMJ/aJ5i54dNj04yE8IQVG9TxziekErvPbuSg+obuG7o+xZR2XyiYBF0DDhjRzZNl8
VtvKMT2enlA/VrBdgpb1nG5/4yeEI47EJv0/nmXd52LC+GWmOrteYtyXSu3XA80jR/LUu+HDOT36
kgwrwPVU1zFVzoiqTtnUnwCh1kDNSSyKx9b67RpDSyQnoXRBZ4UT6zbNkl2OTEzkd8QeAxg+8KAt
54kfZeqXhq+fvNSKv+QSJ9Z1SvFuHZlWNOAo64sJeFVgbuOwJ/ubbAARf1S+YY/QEXATJp7V1EVc
oRG7mcuDiWNd+ggvicBxz2S+X8LPX415JU89OznZ+575MbDivrAD1qYDFyR35c8TgMQtadf8gDeI
c0+t/zfFkY074X2VJN2zv/N8kMqsrxyW/XnmxGidBW1oxb2C7aNT+ri//XIXq4idvm6HQHENNJl0
4GaoDTlbKzb5XpBKkQxaxs9jQT7psrr1xuRVako52KNB18D5AJOTiVDa5YNo8FUA9hoXhhIp42T0
f6a7BXhLcUlX27VwWOAKuRppVdEg2lJZOFz0/MGQK2Bj8tEyUdVT87l+Xgxvl95V4NaTZXZDFGkQ
SWtk1TwcQ/IeqbDgw9riep89y+7jRf1y6w39SW6NdCc7ZKAy8qcIuQR9t2nApRI/8gVaZdEHoxLQ
OGv93+AFWvUOcYES5wycwDPYZl/GE18CEBw2ryDUo6dmd3gaWIGSiR4POXQaVPJLz9bIl2mH8BVK
rYWvotbioi5riAkltJFTYSDwVLBdLyYp1gaH+DUe7HjH0Ltd26m38vYpoKdasbsPa1Crfv8SsQUX
QhBloIadcJllow1JiyDtg4hPTouC27bJEmoYuv4J9Gmrl9gYEwamxSGgNOBWHx6NgvUGnFe4BF5b
AL1uaCP2ehpu9KSsobtXjnGJRGsYQZujTkiFfVDOhQRoAa+oxWRJMzVo24HqisUx10NgUhZYLxHI
aoPo2QFBXIpFXnn7jxUZQNwcAUUOQJLSVmJ1ylRftIWLt4itW4c1nfT2iDwKljYQGKNwtb7+SmF7
8A16IpGrOs+/AcsmZqFO3NTb8+GL0/CZJfARf1N0/6N+1mTZDdmXuSmHX9czI7bKkP0oCFmrTg/Z
BdqSj/6nBLSf1zisC/S0vVeFmjN4y21Q8bN7/+qaWU1IGWPV2qu5oVotcd89rmSidG7N1N5tq4fJ
rrtKEZtIjJCrb4gilsGJ8osuXMW0Ia7NP6nGHkTADBWAivvvHrTYs+45V7eo3yjtSKXr8n7Dw3+X
mApOaDbI16SWRSrVv5H89DvPGXAR0tCene1NSoIrKMjTLENnixE527opXm3yZ5UTvKfEvJyscnYR
AqG8ABdPSAn4EgSIFWhh7Eff+kgOBFJj090yMfSJJlrxebFJRRLwyRehr5GDpEwi84ytdOCDASPO
nQDrFb9Q0EzT6t+zQDAajCtQZ+eRZJXgMvr4lDc5sHo8T3lOPIJ2k8WEol564mpg6kLzwV7VOXTS
sqsygnAckUgjcSTRl71VFETmf8HpNerWdOuw5fFb3BCAU1zlnfQI6Jy/00kk9S+7qDTIZR9J4QeL
+GfYhziqBN8CeC1jFuQFHECSg+mbsM39yLCK6cF4UOuF7waUwfCsQLGC899pEFtElQq5UqUyziXc
od7Om9awOjYvxh/xQnrvNQ86tuiI+r5wB1rJ1wX1I8dPeHmqXOaYYy18ij6Wh1J8wMHDM0dO37rl
o5hLbKNN6hDLQOX9wjramkojOY9fPoQTYt+N9fTpYliSjNn7una0VkaycZ4/Nkhmo90gYYbX3/v4
ErSs9GpHl9/OqwBw0ZejKT2mB0J8VPqTy1WhgJxkxgIPvg+yNkuKx/ZjG9U6dptHsz6ETGqGd6jl
X2xQH3NM6iOeRn2D2KslTfezSW02eonFdK37TXDe18sZygV1rURdYs3aXd3QPLo5+qfwTXeog60x
LiVUzfeU4mrv6wGx28UNlYcB0Awy8XkHyFFIKRSchGFAk6ly7+Hd8i1A4JCImUOwTGJ55lz6TXhY
CrLWWN+jJOzE4jGeipVZZv8dKmAJBJlhJ0Wt6crSQPrDJafYyoWHZtw2JxO0XT+2hJYdsefSpd3R
jeBaZMJvjQs+Mu54etxzwv/tWQ9HTtXduaYr0IlrZnmxjtcH8uVcFhp6XsHTW5B7gG5RcpJDi9KN
GLCwM9BwCD2siBUHs1VYhou90SkJ0h1sB/ahb4a+kSRO90u0nr7XPEi52jel6+qLv6y9qzKAC7+R
qcsI8+rjdPyb22ksBmvvQpBX2+ujUo9E+3+D+ZFjb4kRZXHRaliBg2poVaE2E3/AHCL/+8nlDGuk
2pgga9OKl3hXy1F3HXNLvsXN6BF7Qpfrgqc5gT1Gm63jt/nosjr1qlBUDY9CP8RgNCTvBKcV7mex
Xao4O1B43N8f3uhVFW1ujzBew9OPS5R7nWF2hsSYncZny2OXpIVCzBUQdkqWTu5D5VX5z1RL8l2r
KPd4jp+2/ksbSCfdGU/eKGeIwiyZVtlvkDcduizlN1gX1AHdVKsgcqCV4D22HWt+/qU8vF9qX3+K
NP3AXXLIKX9JHlpg9gP+4+FB7Bt+evpACxkmfU8DYj0JO4cuKPTdo5PRQ9A43IMgTaManrMcDX7l
l+pnDoYoazDa4rXPMcSyFQvaVUDJ2Safg0pF8Fs/rvDKbl6NvBAHXYlYGbVX8lFwIYBerseFc8gF
SkAUK25lQLLnvHbYu6JgGl6mR6AHb/vst08yE64dWHfL+EsYsXCr7/tpSuy6ewd9AOg9KyigRoeQ
RQ7YkB3PTBFwm5noIv0X/6zFW8T2xz/V5F/mVpJzwBdsjvgLBoZ7TdltJ7VZ1LVs6FnGHwsAsUpe
3xD2xWi46PzjsJ0WGupoySe08D3iC6372JJqSZlgULAj5a/Yy7GpnLw7LxB4ZNhME+O6qpQMnsOr
0uzBdRcR2YOtHA/rxjmBMy8x513jwMd7+WzKL5PP1ZdvVAvszCsKlRyXxL6abU1AyAN7pjq7EU4/
iYmsF+KNpOy37teF+xEN9mqknmDGzsrVxDj9I5FILDVeaJottQUBp5rLcNLMMYEgVMV20Kb2JEdx
DXeEFvBrRePhRh1ztLLv5pxgGRWb1DTLEQEADBiBpaKEhL5SfeUIhEqAKB0cflNyKP9VS6xVDYy5
It72irFGLSozTZ4rN8aoMUcMtGPUZLiK7hdWwnNF5HpHHFDsRSh3B0TBD1AfDN73PGjrHy9pMIWF
KeAT0fp7RmB1OcuLJfN26NpvgoqLqFKZSglaYcKkbzbB8jTZcTcIwasa9idA5742/ZeEPh3Jc27A
Fdy3WxANsfdybLANJEQzVrFLYzBl1slEOeszV52WRsq1exL+suUtWQyundNchmnBlGiUF2uqNb3d
aop/kMhhqr2xC714aXmCkMDfwxKMwViZvgNM4+wc/Te1zWjSkhpe8aofCyP7SzDPiM4qkt+XT7QL
Et1qwojP2euImzIITmjbmfTD+PdH69R37M/3gFfhjq1yZFPrZ6yqNuXZh2YGNK51v4l3YAbSB4pa
ssZQoPjCHcOy4TMLyfnKX5SeZhIOBqY+uw1qVrbiOg4Y0W/xiekngDLOvqugKAxkzWWR22M58+YE
9fgUFiWzdwjSYJye0gYV/fT1Gv5iZg06/igwd83mn57cWklYW1WdaPrbj736UBIZ4N56/FsTnBE6
MrLeXDhwYVCvL8qnbE76Q+Msj5wDkrhFUs+W3NO5IGtLgNQ8Q9vq8UQqZxHPIs6WV3L2Mruu82yP
qDd4Tnt9AyvpZ5/tvolik7hOXgPdFjuWHDaCu1Fhu+FdRDYxPZz7iZwYmE/2WJQzBmX2KYVJy9vs
tJciAjYQuzxdYwVn1JbUFn0Nz3I0Sr8RATcixeMWK9tjEMutODJXJ2Ygv+j9q6YGTsDTsGFvMtQ2
YDtsjqRndYDVx6ZRZQkpVvk3KWptRQzOCyDDWigpHQXrUeWuU+RLewTE43lkzQMHJS9CBpi6gXS3
YKcfu58dBBp7ap40bDNcaNDMkbtwZCdxtg5WAs6rdT5MHdj3/gNcWYF8R122LDPoSpyQDfkt+JWP
ynlpuCg3sAjoAGd+nENifpGH/gAMBNyIlHp6MKsNT/ZcsK6lfAJZUT25e3lNMhMfDTvLv+g8dlDn
cn60nJk572CNZHz1FrjAGgHOe/aUMTTQsahm9bHSpMUfoo50OOC756Wab74CbDxw83sQ+ZSVL5U7
0QSTvJPOmQCPptBRjIXQZeeb0oMWWVRCJ7BKmXzasSkBErQxgT76mCkQbwP19pgHU9I3iQcv/4PE
TOXzPvNesi4tmniyuIv5mVOJjSwAtq2RlQ/4j8TD1vrbbjBiN8X2zj6va6RHKz4Fk/TQQHqx6c24
eGo3KqXqgZ/XKitdNv09HlBnmQK6UL65X+b4lOS7g5UUCfBzJieMLB/uPpceXgY7LOF+qowzampl
hA4FvmIsAHo8tq++wqBN+btalZmSoN4OOSylEMxLlBH40+lBx1CW+qO4j+TluY0CX69zA94xXoWG
1JYglpvcQqK74wTL6Qc/wcdOpuvHMFWERzqAxaDzCw94L1+yAtceAFGN6LeJZyWv/vsHObEg0ZwG
rDgIwqYEkmSNhRhUIPyNzCQWtI9amNWd33Qt9QkgAsLn7DFreuDijGPHM5QklbxTjiPZb2TvS9AE
FNiTF9OV2AKtvW1fKkJVkEG8VyC+Y18MI4muayxNdLkSyBs3C6/xgoXAQ5EYPBtl/tDj1JMYKgA8
NL8ozgleTipaLSHDTz98ionXScEhUE4+0xnP7JP/nvQuLIZFyNZStG2nx4A166WdMLmBuarYPchE
t9WExyRPI1m5sJ0QKXOdsJ1OuoXjBpzamtMbxIP6JnfOvpU/PlVivid3SnRnojzUxMWIXmBW1XxF
22Zu4slfihpM2iTYlc0YEC1XhO6qK0e5f2kEZu3OW6TWFgC8lE9cLSCCTqHhsvUE9TowM6lOSFR5
NPj5VJsTth3DrpjSnI1TSoQDBZUmY/lhWjIgZqpr+6lkzHVf5bBT8778o+CvywJIyrsiIDrz6OQE
6WAuw1hz0nz1goCUEIu9NzSo3OY5yDNLKXhkFpUm+t2B8ZrG5SpTotaFK9oIk/UaY8I0pZ0gUEJy
ZAx9b3c5RA4zUHh85HhobdL6OLk6AdU+tBidZlKtvKMVUyOpPoncsDHi5Eb0kiDklV2zX74RDBs3
AIFM21GESNc/vLfZ33IOAj384o4uQttUBpfqSXXW0NVkZ2pd7ZFrCwb5zamGnYaW0TwwPeYpG4A+
JXiMbTXL8ahwrcMtVZRQ5L36O+HX11SbqymCxbW7nqJ3xkXvitBeMuGfbfFgyX3m7BcpakdU/Ihi
IQFQuYaw0crg1Nm+pos0E0JRKRPz9vavUV0eFi4PbgA7JMCNrgUtvI5Veojca0ko/gzSF7cT0xtj
Viazi1iJQtHShOhgN1MEGnS3u5qBl1GQoY+zQJspj7OVBct5IWu3O7Y9fKJoHa6EYdBixTAChqGu
y1LrKV/zCSDFqiIEQsI32Kr6S1K7y9tl+66u9Cvr1JyVJHj0gcld4ia+K4ZjSCcFgbbKZi5uInAq
v8qM7UicVOuJhlzkAU7sHqgB5nnr0y/wbJVTWl1J1eCW0XR5ctHanHd7AlwWIHc3Hbh7aepWXhlS
uQJMvMLHnRRz1mgc12M4lvxKGEB+Zucph5zArZABQT5Utii1OWF9FNK/ZqzWTdhT235buCUoVepe
Fzpkj5DdhD5+g3NvElngWhKBTxcbOHEm6yPTAoE1uy1i6x5xCpwi7gl0j6iYnEtXISntEMBHpWpW
UD4D5ZUelKqOmcbWxbkYceipBRDo1jG6nqNg5TeXWHzHWrHHkjrJSPXGFddaQlCF2RFojAstPzUK
7X71cf9iupcpL3SvMw7iOLsEcjgVDG8J0alQuztE6IfXDCIDeRJGbVFOL+zCnxeQefuws+teeuFY
vZ0Mxj2pttYSw3Jm+uk2BmoXigTlGYS/7uWp83OH7fNb7tVsZxolrgSdsT0XaPhLgWfn5qUfemGh
Us7IkuL13Ltq06T81O4YyqiMfHV6lR/xSxOc66aWZUG9vwbTftFVt/xLr8ABzWxy012tzQYWHPmS
frQ7t401zeI2N7rzXqxkGAgtbLupyTGxQQvY3VQsHA1isXFGC/j1aPOHxn2EwBygjr3WFeAfBClm
MRBpwCNnnv7h4HVe+0YNjxjcSS73iQnvcMrv9qAxfP3B+m54bFkMiYmfoa0xSfLd5ZnglqYQtKQv
RlxwzTU3PBHhm/qIdaqyrejndC9Zo+HfhP0EGA9Btbb+LUvY+wG02tQSOs+7ey171AT4WYGtJm7z
7DwX7tdPgTIaP3td0DH3b+AIhg5pf9+R2tk5GWaqbdQeHNLT2j3eCTIW2DU6Ik2BMG8/Hvx3iMy+
3A+nGkP8mHI9JnmZmQ4zpu7HApaxRSSVj1m+76f+VZyPF6AGDVw7YgmxH5+f9Qz7DLpMH6Zmbk7T
QiIEsyo8VZwO7jYCWkM2h9LqefeB+tbQXvIM7RN/0eUGh43dR0Xp7Sx8cL4XPTjX0y+X2IHUT7Vw
+mi9D3AnjdIVz2cDdK5FdnllFoM7BfUCb1X/+Cz7N3BGEwMFk/kAkqsZedpExmHS2NSQAl+XFoaG
pDjZLGtHnfl1gIIGiTXhDdswvfeWv63NnHvmtHTjf81j5ARxmfhO+pGktD7bLXj9XAV7ShsJUvRu
dvY0/helTfWqnhTeRtDTLQV3s1dFdlzVEMiMgk7Wu7X7qanOivGClMZlMyH15CjrszNWJi6mSE4/
s+Ekxw2gW0nfry58vN5FAPKb24ra5x+s0PblXA0plqzLHlcJNoqZtixnGdJY7kfReLtCxUqhiK+y
PouJV47cDZS1NvGJGBJ8a5q+g527mL+DPscq2BrBOVtXUXge5Rl+ZJfW0trQ8lS93Rvr8iPplIGO
AuooNNcuUslQakXFOUaNjQ2pSp0MFOgDwTEqEJigNUpFMGPn+gAIHoUQi730Cd8f1QaQUn6j4AGR
0kQrE5mmdc7o0fe1AbEbTpygsEWPNEyTl4KVYW5VXna4/eY2S/gF/jy0st6bdQNhuycN8WNUl0RB
jeSIZHefYJo6HUjrXWj5V9xmf074RRgUkH0nKemqP71h7X0IuZUX64ixcGuz7/uFWdRXiRyUbdWJ
Y9HbRYs/SzSGhpmlQpJxzbaav9yEbwJ5YFl9PtgnCVSU3sqX/Y9T1Vl5OdY79YYKVgR1d41c/7OB
clMveuPrbq6fy/NKiZ1AP8K23mGPERhVprI0AVdzyTeQ9Ojq/g8a6jwONCE5J+btBariwd0KLjIM
Mgm0MyYNJtBH3gF/xv7epkv+PdUS6HXLVO1ewEOb5fWeQskeDklS45reyRsBUdijjz6BBAnKLsoV
3m7EF1WgDbOPPR/XOMNLuCjJbii0TU3WCMsp65n/OI+36zxpfqAvmzSzV/Ktw96ZLXoOH3A36kyH
1Kl+z6z2WLYMBtk5BauZSF9MP9Kr8J70qi3l9BI3nFUez7GY1NhF/HivTEWvuvGxvfl/6HvAnOxY
tt9z/PrbUvO4o3pTHBdfMZWlAs7BSELw2iuqYKxTL3sSVQb4Tjeb8Jni4erpeaFgXRPAJFQpOFbN
Lln0ifGxKUTxMz7moQtzQX0b5AMZem4inSYggWvpF6oeWxqpV8jthl12czdEuOonVaAMTUEI0/UZ
cjw0pc/kQFVCJYgOuh4VtT/ZsEUiMnn6XZxLc5LrJpR8oN9B7t7V4o1iE+KhxRXoL4bPm4gEdFRk
d4rWR4dQ7hd+m+dvathxT2MPKmDecWemvS++sAHJJ70M5WA2LXf+juNyFO2TnHF6gzrrxjcXLo92
uVmPsBjpecTyuZgGHa3PQ2KEIxFedL9ogX4ck+OG2KTIk3nDc+2Resz0lR11oDbooW1mCRkKa0vh
XCKtZ/8QEekfwcX8E/XS6XkLm87bXfG8ULTgDSUQ5+5va3QHkpafJbNaH9h2DqyTlzHpQyXf8glh
ORCpwaF6BONnNGYuUwDwwbQkfYX6uk1pxHlNGtOD5VDDhfGkls8uzQfoaPRhgvpEzDUOp72V29Wx
MFOtC6+ED4TmMKDA+XrB7zvVrHRRz0dlA7ZxNB31DDPv5BCW8FR9ICIQJQ3xdJLDWeSASNQSskXH
jvmHiQQzr1BvkFHhlIGKQGllZWh+DCb/NRL/b0DmKjetrNpd3U8aYykUWLjjKkQ9fRI2yrshBerp
/BfGTb9Rcf3VBnLIrOmgoTe28os+qC1yaA5PHExyqo68gsRkpRsiLqlIi4VkLIaAdWh7S36HgURt
aJxpuRZqS6jDzd8Hy7PS71zrT8E/es9NHt3RIrIOaSI990Fvbpz1BQl/qQMju8gsvON7PxyvdV/b
HDNO5GZsHD+SxnQINXnwJJRef0bATeTutfkVJ2aQKB2cU/ZR4xt3ahSbNYrrpFWWKvBG/A7O0FEO
8B42tkH67R6w9XG0ZbaT6Mh3QiqU+OTokGuWQzhEMO0c0sXELzfP5srPoOWdXV6xTqJfbb5K4VEB
3bxjaJl0zYbEh0v1hUaWzVRrQPz3HG0UZNXnyMRMZAp063U86HTuKpRVUPn/qDavuwIVOrsLNPqY
srDhMX0u0nJ8z/tuN5w9+FJOSGf9qlbwdZf6IopmF9xWMGitpNse2OkDwKLkAJzZ5zT1QOkJOh4X
MSfi5Mo3luyd52pjRNDi150Vu4z1n3a2MA9uLFukR7HX5rJJb+r5Zuuxki6lVlRaUxpVBfGG14dZ
yAsTVo+M90OIv6ne2F9iXbPeBp9bm9xFwu+SKIHXkHEucRUyYBnHHeq4KAHHt7BmEsAI9LusnjBK
R/2rembbtz9pUyJmYqGTuaSGt7H5caTb/2baXsYNMj/OVJAI7bNwnw4yy5ZHDKwqYjw4PLqWCESL
M+ynEbJ7fCTX+LEfZnjXE6rG6YTVzZSBqhZa3eKjRb7ZogWeEbArGK1sneRcGLeZjyTcnHpb/RIt
ddAlYxg5bnVPjSM5ZgIOnxccQK2c1ZbwOKqegVaS8ZY655B7wuYiUQLtk8H4cZor5P8oczcWeIg/
Ed6JaBw17AV11QByJujCIzZTn+2OSF6VUqdDNk5AdkCZpxtyFH8vCFggYhTsm83aGFMl8QSoRDK5
zx5AzPiWZNRkKYOtENprcm4ETulp0hkATe6UWx6e1b7tq8hE/6cTPTCByj1eUwrlmqY377jVRl/w
W/x41KHs2M3sT8JXWHIei2+ptewLxkf7vO/GUivycgaev1FVuvzr3YXfCXpj3eTScixe1mVj8nXx
vJkO+19YZcbP8Jjbxa0lw16I7gYhh1OHubHmzon8xRr3C6MdiFh/RW1ef4GyPEtqVWo/qJNyBq76
E2sNOuP8dSY3cdcu15GhkWTU1R8ssYQmvkpc2BwSpqmgnTO9wZOsaF3Wv0rFp0b/ybSb0T2bjj0x
dREOJ7LU6l2JRu4Tw9Ci+KEg2T0qo19Q7e5KMYfOkq1PH3qM/hYKICZy+XW6btgnU3kc2IjioBTf
MIKl17gqf7TeywfNwNzjxmXoxURoBq+U7P2MQD9m9wF/Hpmktw2Agw++/6qidgwRz+jwQo3G4ny6
j9FAqptA/lfeouDgMmdbvpnaS0l3Kzgau4L71ShutjvYVO6QiMlZgtuWiaHAlxFaO3iwQLA1V2R7
9wF0SlgyPLn6Wxz3fUM4JamvpgXr8Co/oclGdZJAofPc0j9vQbOTYNT+eKaFvbS6k/wvYvjxVHSr
fDEoRzHtXxl3BA4A3Wl2m7v61fCiXmDTH33WWftxz8tH0+KBBFdd/J1Q/rNpbufsXT/FF1RpyNzj
ER5JE0kvH8jtoO0pfC/UDw7t6fEF/xaZiiPeFz5+klNmtDrHACd+OOWJEnbCT6VuPQJ7uGTSf/ZV
2rgiAgHsUv8LCWVJWCbG2ihOmAGH0vrbE15tgoQH+AHU+dukJ47xkDETgzWwNgIiEd7ltmFXLSTk
4DvohLq+F4/gOJ9kwKfqDbdKQN3sp16rxjs93anqq1JkfKcjjwFUfP4Obdm9of0jGSuWHmHqQeBA
3Bu9k7pg/qQ5+RwiJH2MCGx1IJZ1j+eNrO7NNJncS1DS/I2JmLZfrQea5OhrDwyvy5xsZTh1ZyH4
X6iqRl3Jzkh2pBLJo5lxVZjrCGd5J/KxJEHeXJxeabhiJE52rdTTFQQNhDwx4kcTMcHNB8qCCp3u
iKZYaVeOgnGwyBxFmzJoahGvs2g2ioSRGcXNpZGFQJWpHklODJA85lJBP0hsZ63jukPotC8quSyw
qpxOrVcJI4gEXrJXmzE8TW5u17Vty7lyJFKYf/0k6M5CSbu83H/H6JxappeTpviZ1l2DyHgJwFnc
JTgtyxFJ83vGiuDKRZwCKHLnjythQJ/Y8r/8ojBkCmbwaZmtW3Wv07eXDY+ZqkyXudF/mAqKBqzR
1TVqXjP06tL7sNaZWxTrf5PaFoDGAyG3slT0xeCimFl8gCREFU+9xgVDCoRNNmBc7nvLAs3uRnXW
nI9/HvqLw2pctalxnBME6ZtT8ee01P124iQk5Iq4hSar9Z83CxrewhLIsznHTUcqXM+wgIHGqwfx
wHtUCKiJvHXYzGdB0wEuiy2NGgzrj1RzEl9dfPRHOZYMVVer3mqR5ZSUbpsAjkWC/AH5B8kKsOyH
sPAO4VSxAbaGcM8OacGzeJlg2/eW3pgMdN5vQNZWUch3oEgxSBqbhVYS2IR7tLYuXDK47qprZYf/
Pb+4Mn6fbr1wmWjHPqLAfQAirZrnQtGl4+5ZEawWzfrobHBUFqVdsN8jyVgen0sLpaYHx3xsvsG+
F6ZaggguyaZjLo7c4d7EjDg8hyzdCRiCBHj7a2PLJ3cDxXFdV5sNJ2cUGTjMutka47YBNTtof9Ds
v9oLy4HjpouUy5HMiXDwXon9NMOlaCrRNtefLmwZfAARnuOdLnCVKxVxouNcII9vqP9DHH1rye/2
ZbUN5O8txMG0JcsThdmhrU/oS75FGUgmzUABrfU/m0s9pCqGwBFsFB5G2ALRe/vDayzZc2IW4l/d
2qt/QicYA/71o+nR5IG+TaIUU83Agk2iEEXkauUliFnLdREqEdfaesRo3DmTI0fnAvVPLZmF2WC+
jj9wBQdt662qANfRe7wHKuZ+88jFpuLPkmlH9ERCpvYrCp3DyJqrJuzSt9op2BlKSKU62OMwy4bX
hVqMxuGOFu8qde7LMHmO7qew6VwYuqvjYQqg8kfVAz1NlvEnMd2zR0Oi/9Q5yZ13CgPkOkvkKTA4
8dAnwqDkcuXGyX0VbCBFgwSmeDi4zee0LSPwEzxOhPlfQvyVw+o6sOviRnZNsEwVGFI8vxWRczlW
2HqFRHA7a5gnh89kH+9wvh55KdONp6bwRGhYgIPZ7miG2b3eqt5j76rrbYVMuPsz8p1gaVGKthDr
Lt83M6IBGQN2ADsyqae2lR7RZi5FviDQcjpPgRAbuuml0TKRyfgJJCxuWhiiSMyD1xMX7J5B9vse
gZyLojLpj/KkvgiIXHOvmrVTaaUgYkaxW52Z6TrqxI8Ptdq2Um1tjnd1mttY8FbTpyGTZoMvQlWF
XWhTXNQHlhU2aDbjqEJ5W4hPO+D/ToqBuHXIo9q1ZTb1YW9/FQPUrBuvMZKaQ4rfKpFg7bM5ETGM
bFuQRcKPu9/rURFRalsaf4We72TTr7Vz6CwpjM/7E9ab2rFPAy7Ft5XEtjOcw4vBMacj2yqUfOeX
fwxMScCMvkr8/TR8uHu1Bo2kE8tjWj3E0Qxas/8x61HQmajKJcz8qo9kV3dYksOTogqsnOVDtbAs
qv7uAPzyd7FuyhPHUrFFfcsMQuWWm+fOtrZwOQkRc/x2tUGnTclBWBuVVJC7XSzpKTuKZK+AeUyy
2wHBbeBpGqaexWZ5XS/PJb3VH8B4/s2NWAccGFDhwf8kTLQQtCCjcwIlJQUMUryEMcCm5K1p25VS
chgUKE34JID3R0FeUGXGvDb9lcq1hla6FTFiwCKIGj3MTnhw4c3bUmS8zDAG6Avmn0F+nu5wOyh/
qQ5QfSLLzC4FxAbZnwis5VRDSSp+DWKhtEVYEGhyxF5YMLsnkIorcfCqqJW09CHjmNfkir3RknEf
2nE8dJyI+57h3vb45WXCoP7UZd6AQjr4EfYmTEPm0BtGIWvxIqwAWvnpOZO788qSLer3XQn3osbb
AeaZkL+XNLgLoDHTIGpzxmnnJcxBjCgWF1DuzLOCUHlBgDn07IaSmFlTxB5i9zZ+K+4vjyKV/jjH
3XPKPY25bTPn2AQue+Wxgn0nOEhIl0JNr944JnMf3agRm3tSQyJKwLnBF53GWG3FxYgdK2xctLrQ
F1QVG2weql74k/r4gQCiiPaWXvTn1fs6YpiiGQF5pwh6fi2RbGoDe6yu1YBL8v8IVp3YiCWgfbZH
XzfyWLAwM25xEFIcKJQNVNRJ8U0MtUVxHDIDpjL65jLqvjoyXjG+ZwQv+MnNoeu3u96Wq0gJoEay
VDqH3TzbS03ND42m4T0pUhzY+hMHEsMM2NHK2zAlJusR/6+gPv4xWw8XDZ2H2jB3C8voe8dc2DEs
Y0nFoBC9igBIxEIbGT/54DelTbS0RYMbfnQwAomf1pVyFDgFyd8UnL++B5w+rgAlSwqrb15WWQvT
4npQWoUr53yMxjElTyOTcK49Fyvf/C5alZ1RTjn1AFMhlcuD/9ZenKPK9KF7GiZaMzOYFv9EkVV8
LX/1GBXLQ8W66TOlrl8Q4AQg56REFSe0EDCHy4M5by9ggA/z8+emvuDX4fE1UOi+fspQtRQZCOiX
iv4NMdQft3HNw9tBsil3hqg2z6L58TW0kGQMCPXQmLQ2lrJe7VBccfRjDbG2E3RYVVvhO74TD3Ej
PRHpTAOyci6crD/eNtHVmmKf+f8I9+lc+DrSly5qOM541nEYIIDrUAnG+jV9nPA9D4VA31XEivzh
PjBLpmDsOIWPs+qJ12fLPg4hI0+V0hc3VRQ/CaGMFS3nn8aegIhEgCXQBqvc7uuTSh8vqKwkPRHF
QBaxjWyU8s7kma2p37AdDI+U17+lXWJT/1ZcFBOz9lY/Lo7NZKMMkIiURbA6AUlutysZDvu5J2WU
buufuGpX7yR6M6l2jOT47a4r3ALlVMVqOeurOyu8jxfVL/yifa9cVhVroyd0zXad+HVBUm+iVJ81
RZmay7cdveutqTVe2+4yVGq5Uf2IRELz8l50+Z7LSYILn/z4wCsriZHkwOX6t6DsNz04ltykG4tv
1wieb6NwIdfmEWfOIJn+PpQeS6TC64f2SNvip12SPGGUUAKwgTjbQjAdp/oxr+gcjEREmQe2qiRY
YMjcPcxDO7DRM/Lt9aryWJ0ghrVBH1Lns9lpl7/wrI5VoL9IsKgLh2MYwlh7wfQuoV8GqWcmpvYj
GwxAo1XgMYn2zmM3rimpjNyCbihBFtUQ1TJuyUBN995ai2smYecblvzYxYArTwpw9Gk5M2iOFnVK
XNcm7j1/tytvTuc4GtHPCck9CtDnwhAmMeFk1yfPrPVh/feIkkfGrHhM84aD9unKulHSRYB72nv6
xSwPkRrJbfVqIzJ8gq/CROHkwDw7rk/v3D8MfmkQn7hHK1/Mm7hakojkUkvWeFnSBLLZaWGTuWbE
f1cCKpMe9aODzfCgvjzvsQ12AuA+Ng3mBOI1yKzskz82u7C5J3PQJ6WGU3O6GId3OAQcKnsosa+3
z32zBb6YhyUhFxSM+3/xuBwipCwwVmh9Y7CBdK3bjXCYQmUZyf58kotn+J5HGpGu/saCI/y7lZ1p
UjjkuRJUmxf4m1Npfod97p8p+q7JXknLuD9MupMNefw5oZRfqlGrKbD+UqjXuwfs0YfD1Q482NlK
UejcV/EKHexgRkcp4xdJy9S6yFwwJ11wikrYHdHQdT59LkplriO/GdDGzWhRk+qhw/axH4jyCUkA
CUA+WflUm8YRQ2ZRrGkvJbsgRd06+Y5vXkgn5BLGoYWF8P7Zrq+8/UoSJd/FpHBF8AEMZityT2DS
MDYlLhGAzS0W1L4X2XvZhpQmJQ1ITAuKXDgu+pPJceZDopFUJlpCruFDvN30DB6oVk5c4wEmVOnx
7UfBFT/1wyPrkA27CO/PXaGXtuH+Hv0W1lMBXO+q/7rf1aJLMhEvDM8Ra9TZH46Zk1RPGgXAie4y
AUGDduFcm8MT4oAuzUtSLosqd2WWq/fs+I+vwdQIT1q33BXCtgSneunWzBRAhpu4YULxZo/KwZ7K
ZIEMNr3byLK5iMKdDizhJsEQryH25wWlmDWegdbmpofttNVfUZgE1rZjHGVXam4DezfpfQT35/xQ
gRnLxKYykiN98xcqd7foXsRXlYvBOiTwvdFruYpmx/yjeGknNhQVqKjlIQi5VoImweCv5GYpPRlV
d4ATqWiyutRYvV3NHrpg9YYfuMOF1JLO4dWhsb6YSOvRXf5VVCUrOED2bHozVKDbcSAV5uI6ZZQg
WTvRz8T7MKIsuBbPrWxWgtzKv7NZ8xcXALXILoDK/La9qWxfV1fAZiV8r3T+pN0XLM/x564DGtsW
1a4MPJpbXVOvV8iZObzuwdiTpOqRhg2pjjYFO8r74YEqo1ADqh3nZd5jz1sBeBgSMQXw6MtZmpTD
+2NkWWZMI+Sv397SOJj1dt+xji2tpRbLYq1XQkpL6PW5FeV5PyYGIc6I12FiBuIwMpScxxMo9Xiv
I26XjugZ3h9VlTm9la1Z4QePmDh3X7j7TQ98W3Oeh0tz4gSwOj7m2eE5h64h21b2jIdpR1exTEnW
bBpGTFfv1pxOYhv3xBAlgvvU0dNJtMweoCQ0xXxx72OkD5jrEwKOwt686Gv4Xv58n6yv7+Vjh+J7
YZW/FkDUsAkzWjRNBh1Ci0/ytujm4BwKZuT5m2IfJ9qih0DFocR3bZg04ogodxR5m/EMNZsZKXts
WLouY0kIC0MAXHuG2USas+Aij1+aNTkqz1aLtw4hzsAcwhsgSUqDQpuZWKViFkZaK9tzK4pVrtW+
8awAXaFMffbsoMbK4H/UOb9WbwW5HsfLOvbJdP96SeogKzAU2FfwWfSv0xlPaLEJmACBXQX5CJAI
LC4PROa1rKPY29UnfUzn8epK2a9s/BqmR0501m511NWvemsA/D4WfIUsAp9U+OfN3nBLd7lmlsqL
uTho8vLp7ObFHtgQOsFpZaqXhE/YECJzJiTOOv1D4cjFq19zretewTNvmOpzwMpZ24dnjjCK9kY1
o8BvGEq8Zh8ZVWsEoY1jgGjTuESj1foyEsqoL7KOpvVHxRSr4g4Rkn8HSmCgrW8Bgr8lSxrhVLVp
cqiOTnzwy1pAi+5ro0SshSIz4IvTcT+0WYBmW9lQI5I7P3UUq83vALD4/E+UBTkttGVqyvY6AkPp
KuQomtwRkQ0fDb2dN27XJhM4MwgG4YOxABMspyJw9k3co+eOu1D/u4m+ss0CuCkSsNfSbDLJ3toY
XohJurNiE9XKllDkbgq2zBOwGdjSnMkDXX2dKf0H8YpdqJkB/+oYvK+/owojaJrbumKOqDREqm3n
2EkT+bzE2LbKe195+An8Qfoc13B81qjV4whGdQLjsYVmkYfIJ9PalgjzFaRQeTPqwehPTFse4sfC
FTNdtL/MLvv3MrAqGfmn1CegjTc9L0KS/ccX7CSPxkX4UlUTOlLSbU3y0EEShKqcfnNRUNXGw7p4
FA5f/Q1kIQF25Fie9SCyTBGwnTbOLKAnAT3q37exeBepMXUmgmv4leNqjpa6ncBj5Y3rOz85ZUGy
XBfJ8+jd2pRlisfuP4ySMZYzV+KMx+bLi5gThgRReSuytdMyV2GIQdE+lUXF0wnBzR/c1jmDYFJH
WWpkyO4mekMymfPp05RyA73OUWzHtd/R8jqtF82McU1c48YvcOhFtZXc/P5/KuP0RfyRWtWPofes
Iwq5ri7885PmIabcCUftz4838rszH+SH7PbezGScxnoaoeraeaGbwDgQuwy3xIQHPDUJHicO3L92
f6vN6Zsp1waoCnNr1bAZ68C1m3WmQ+V/yYXmEtUMY7FjAzazb1IHNIu25nJm18GGfIRlyTcSTtfV
prVtpsric3kUqkuP/qqxNWQgv9EVevhlty31UySLNtDMCOkTwQFjLGmDiMMQqO4/ruy/U9QUhsOH
lLmelbsJ1pta41QrpHvwmUbcRSof5Irl5P1LGtAeCcRphc/shKxR8OXMFY8+4Ar9gHQxfOk3lr+D
aTpdCPdZGA3qp3ze1GViS6nX0Y/ybVhlxyU4JE6X5t9EPMSi1TJp2rFUaNr3UOsDTX0rqHyZ2VXI
v28vezjwW/4BvYokRsjvCPQEHybNMIaGxxmb2VEIRcH64MkbpDElfIDZRMjv9h3OJztAG7kzNZyX
JK8hlKct9qOvNijGh4Bwg3h4YPZhN+QCx6CDyad3F4y4YZsMFqzjg0urOpYuM2uwqoZYmEgm7SJb
1qDVzqmWAg19PsmkwpZgF5rP+BEWR2bHy8SuBhfLxaxZnjw+R1pNbF7M/w2pdSj9kipIn8+Zva9l
8Lp44gJeAprlicfhDzqa6kr7C4ojB7Ipil+ODsRnTSuxPDUjRyJzHh0Vr+EEF+eYQdMUsJiOu0lG
9+pE3MRZ81wHXIQrOlqa2GtCU7FR4WIdE4yiSNsJEEKjDixoDj7Ezs/k8LCNg02Z/s8AGkvO8UHz
j1mxjhjKClLFXfOiuafJYq5fXucHJBoaFpPCJNAEb2SczSVMAnXolQiO+c8YpKS6yKZ0UrhfPEYy
KHsSwtRf4ZAFb+AFXvPwXwZTTCRduBllwArll/vRQXl8jZ5Ne0xKdM0DdpkbIE+OVJE/8iPH82vB
sxgxR9/IfsPVWttmzCTciu/KHkJf0+iZCo/S8yr1I80VrC+wa3G1xVwIQyDWVITFOjEknLS0HTuL
Js6tABraA6J5OS1cq23cPJCP2OsK1V4zOO7jVTQKNhziBybSMlRZWYoMn4lp6iCfrGSGoybRNdFV
X4pFkxaR9r2tUCvS9p69ZmdcFN7ylTnEE75+N8LcHHzCd3sCVIxyii1BjpBll8gYdS1S/Lq+ZuFf
+Bg7idvZvcGsgZETP3I+kwF9MIpVG1YTf+kK8FJh6NYy6JTs95A3oZNhtTqjpl3T2cPL630bbmBr
KUjFpKx27YXrDa9NOjv63ZzERJCrJz7MQwqzswlDaAnrqsEO1k7Xp0TM4iQGyYnHdT/OXR6Xuo1Z
YJnjEsNYWQqeQe6il+L97Cu92Pzyn1B2iW3gUp1qOa5CF8OhBRsXilx03PizcdBpIcYuJ0c1hCY0
reUgRAxefx4KokRk1oBeVh0jlj6gsmLB4zcxMSVqdZOs+dnK8Z0fXYRYVgsclilbBLaISu1iD2sv
ID1dMx2inRXGwe7w14AlaCr3ROLyKleorr5fQtMNODkuBC8EBfK2+zssWuj7BUx8IHpRsM6XvLiC
OmIL3/3WTIQhW1JV/PH+1NF0s3XnUW/JSpdcbHXCWDEGC6Nyr8svvHza5fUtKJI0T4cZxDeOHWfb
BpOROSOWa6atQxwp+//iWvRr18rqHaVeWQl5bz2HK/O0rNPrprJH3w243PfSeOt8HdIqUB0oSvDM
AvQmUbasFE95KrLo3x0LEQR3Dsvlho/0zFCSgJQd9lUhiaDH0tC6PbtzuUI5gKYNmb0T3yipASN9
BgrPU9R4+XzWwOJbe4hBgVdcNdrGZEZYuqQcONMGar6JhBNzntnWXq2v410Cs6blFLspH540nx7t
ZFYwdYiyz1znYAQFthQlx86Q+4kwLhD/e7daROz9EQyB6TZ6jxM+QEizkVJfQmCtNpj/yl53GO2J
qrmmg3JP1BKcPmygV/M0wL5ZQGq4r9hKONd5TUevvD7GT4ynVtXhNr8NLjPnR1/2t4xHSZS2FHNE
1uf1KHvi0DpBysuVZGv05jVKM5WgHhI//3r1n+O+tCJUN2zJmw8HocluyKeP0wgG1Es52GAJwg9S
t6fJPNz8MRf5WLlN1Qt1jx3T1uJdclUVlJayknlPYXGmXHu67EWxCt+Atk+2KF0JMzQ1m/XeSG5u
t05SUhJ0Ia6fc68z+IsVg6ixp6rgsiH621r2iqNGfcwA4jT5b9GkX4jzQ/gCIXy+dEKQXU5dJiV2
DbvSeGmYoICNrwNJFClz3XlkCTtIkkEpjjoGQ3B5vyEViETsZRByg5Le+aGRPlvtHcOqzNoRRtUt
0pEOUIk2X/o/0IYHrYVKS4hIHhEvsmWjTbf+8REB2GeIbgPIpqgeFE6nZCG5oAXQQLtXau4m9vHy
BCx378sDx24MMAord1R79QV3Aw6ZmNeTjbosAveWVQwm4WJSx3bokeS80S0yvfoTS3FimfyunXt8
aiuaIg6HcrwQD7rYOSuD0/QER+cl5c8gJzSRJQYnMPHwGW6I9IqdQIMIm79ol1xCtK7qtXRSQJEF
okqQid4zE2uUoIJgkaEpliJ/Gk7RTb7XLUF6TwNdS5jHUWMx8UlAKck/yH0KvGT7wiiCf9RaR5iR
ZvnT/pYqokQasKMXLxt54g/vb0gtw4gzrt7Tw0Dlc1TJ6uT5isvchf1oetfMYKJVidkxN3zyFlL4
EL3wJeNejpRMIym98L8bj/ssPk0vOVoGSVeaujMkQNvKfLalGcGhFjU02mu98zdZbCKRYt35c86e
xpv7VONpGCl5LuGxXqc2bC+BueljcFhwttNo4PzQZu1CaOkqkTFoo48laH5jYI/j8WqktmEJbAD8
FW6Rcdf4K2A2sZuBTBWjqYjtVL98xq79sQlkPVu6dwmbM4E0YoVleCD3f2Znlk73GMzBOr1WWoOr
BXV2FQy7oiuAs1WzpvvuKMROMTMuNut/eqykB6mfH4V0D73Tsfe9/b+/nJa4wlHbC6TXAREeootI
6tbX4VxmlfWzP+p/L/UR7UJnmCDyTQH4bdgl2a+GU33MyABAKXmUJsoNt4suJhKgp0j1DF6SDK3r
CuGrfXS9isZqqMRStL71/MXeoA5zQUR0B4pLrdiOA2KiPRUMYZ9TuzNl16s8x0nKKqpD91sQk4VO
Bj9NIZk9FfoxmQOyarSwBC0oaG8FGdwTtPdikJhDEY8YgnUuELR4zE4u0Ca8nH//J21Fl2n8GcPn
CWoBfuCvaI7nI6RDOQ6JOphffxbKzxIMfqn4LyEsoSxg7NMtpa3ovgcTx9NbzeZMlPRfN0r6vjux
yn5NezT7W1zETzyLsW8a3VbdpjC9xBfk99qhMyR/Cq+ZCfTrE22ANvRMwmMUhkxy5ypCBvjGxp3M
tDTjYNc7A51DgN8ri/Zl/7zOay2/CJ2HyJK5FUaY7kZ3+BAqGJuv/eVNoZylTkJgHKoT9etGF/Iu
pRJMKN35+FiRjoRYM57/drAR3r5wEE4ZAoHJCWIzsmw6JSNkwlwuKT5uXAVTnjxJ+vaqCho/uE5m
3PFrSuTafaC+GQ9aw59E5S7MXQxaZWVmp/sfnddP558U7IOmbe2/VAq8ecw0s7VmvxXL9oRViuvZ
vF13CGitmthwwPlaZS3pUJ9/pP5dc3J8E0BVQb312w/gWD/z4088QD900eQCjYKQS/F7tijeim20
sXcpOwDeNmkos/OXymb2Hqdr6rVSEzllb86OpBiY/qFCBHKGDgHR4tRf2ejAkhO2smwLDS7cI7XH
CnFELR1yQdZuNMXxgG7ZCVrofuMAiU+ZmU74tqbuWFrbMKZ0LhgKR+MidFuDl9UDMeeItjamTS4Y
nsWW/2qaZIMOfMTX21E7OaPLXuYo2vZDqdniM1S3j7sL4wTiDG5rnBcLWrFKzCbsPYUnpbfAh0GH
zmSBL5/iGn7WTmKZ2KlWiPWwW74BslfZd5syhiGdV5d3iK8j61hIhmEy1gJOLgFHWo4kDua7QdU4
Jf645zWmnTTUv1h1lI2KERklL/Qf38Uz6Dw9SegCoBwFobK3FJYcTLW5/922MYjzPH7tlAIjsGlS
9sPIRJIPYCr3lb6Ihzlb/ZS4jS7YkWYLwrxpIvQhb3sYw4z4emTw4E7nv6rCRXDUiiS/qCybkOBA
02gCOtza+o3WgAm2y6N0/5eCUjLVO4/zrILMjzXeKeuzs81JKjxDh2qCa3DGsg7K+KwUd17kcPd8
p/8Q5SXVgQdNLKl3j8N6gUYaiVmWeJdi78vfgHlr1kWo2IKbXRHEIvtfYy+03bz/vBS/diXUwL3C
q1NFNU5asE5xKB5/gfRRPAHQ4q9ZBREv0yhfuDkowLRWJp2yDPMtgarG5u+vm6bLHxKR08loQO08
H7B4KjpyavSMQEhSE7jXGABqOlMo6qcPSM0jLKCXkGEsp9+hq7RenIJWfUVicS8mBQT1Frw9cG56
C1j5K0KOkVSyM0L2wqrCPRD4byWy/qdAZ+Qy8GZRF7AYrOrCrh42hN4jFq2XtcNeuYAg7JPIapU5
bRQj8YkgTI+prnS0HGp6RGn7r8S9Zkf2IJ1XDMGEqF2USbXtodbrYrMO/f4HeqUu4DH7CeT3xzIA
91oG/w+dUwznMeRscl5dePTq1ENEWyIQ8iSV7apXp/2pLflhUw1VZmoGRWYlotqUY/iMW06lV/3R
tw6Zl1P92MKHuGEuklhUTw9sOm0fHK94ALAkPsbOoo1lU7rM7pVAY+Pjoy06iEiBoozdTNULUEN1
Eec7f9uUIuNp7kLOj8SFDitOTPLAwvMmY59UwJqFCcJTflhEqioXKmqqAkPSmFynQwqOnzuM5DYg
EqKwglMgJUuJJmqfC0SOxYrPX5CTnanyogsBTqjUz9w0lxobbVPLlogPQoySZGX+agDPIA//n29E
gcSh85NyjyXr2IBaFGv0HncTiLdjgnzZcx+OTEE/TQv3EDwjxnjwv4veYpzzFM6APajjXhBGrK9Q
QhIfrIayTmZom1kkam1fj2wsPYGLwN0W9I3hY1cnulJl+GUG2DCYITMA2L1IKwkLU1aQlzW7ZO0G
z6LxbjemfJQYS6Kcqrsonk+HhI+9mpWK3jqT/TgGa6CXzjcreFPpXaK268oXj8ri1zDoec+sAKPy
cxKPWlmie+B3PzqcqjLX10wVFCYkjNS+figyon/HV3CoLGD92lyszU5hPCB+Ye50JODyYrUior2K
O1Y3nwNDNWq+ghmX6lcIou5CZhRMFhDkoV0iK78JthIfUsiWxi44ZZi1OS/kXT5S9/w9omwPSv8e
mJczn15jSrn3GWzUctsCmPF6rs+OxErkU9a+O+IurYy1XxwSrpeyAavCunl7IDGlW5jlJev3XFhX
DdAQx3gJNm9N+9hBjS85RzPBGsLINE8mbKJExc9tHnL4b9+lMUPwuD0A/3rIaZ1ays2ea++Gip9R
IDNsTFYa6IdPbBi+21yrFVuBG8pFrcCReUhEYQuN9v4ynBODm2aFkiIiB5uiFBPIEksRSYmAO0JF
2kVBesbgApMA2llNjD769t2FBGTpHBuquRB0A37f7tpS6GerZlIyvi5DYwZIMzOPVCgCKcioGjPh
Yh46FIzP/K6fMs1C5yGjQf6bSyFIGWf7ZBG8A2m8vE20k5kZuhvIwxMF8SsDmLKD3BUEf8tSvSew
McNDikvajAYjZJb4oa8WNpOPNfj+oGoMs8pbA6gVYQaqzavwxwdk4zah/L+BqRakNBWz8S3iC31L
vKM96ojrNpOmpofFLCbBbB+0Yt+SH7ZZfd0j7+KwJeeb+4ieeZffBGBWd8LB5gBHKlRpVTuwbo73
nEcvoMHCXbFwH6qG8Y+QgdrWaMHP+d72UjFIHP4aiUEDOUH+xh+R9i277IGaSU0OkQuvFism4SFj
Io0cvX2r3tYCxbz7RvvMkjsDpRtR6dVqQTI1JufRHEA4zsNaT3I/Age8WV/wOSRaXmjLxs+P2q4m
5IS7uY69ReHcgkCBpj+YrmA2m5JS4tL1TzCt5wuoTAteCeLuzBwt6j0m0OBMuIq/H2vrZXmCLRQA
m8OcgU6dqNjzDI+s5dPE99IMQNHn6y/L6/BmaiehLHWrXZLt4aW7ua7u2IH/zpM1YiANd+sIFIAu
nkIZL5MEbkD0/qLFrkuewl/g5/qSCCRyUiWvrbDve8RjZTYq4SnhMyLvmAkKJmkSXm+b8ILOHnPN
Yq0cd+D56f1mi2uw4n0kD9fIzn2HIV8W+Osgc7gi7PRsdpGi7/7LwYEiaMGMXHumNrHgVKtu34Xw
CW8I10JLy/KgwtDoEk+j6fZ+TZaWxYtkDarVVAh+5vU9owiRn7tQ9NBX9zn6u5XkQlD6SAX6pCbM
u6/9MV2RCWiLExvf1olwtyQ5ovEg6aIcQIIY9qhCdgD+Qnstfshg7JdfYsH+ThVwWOn5YqYqkvvZ
I4Cxprjo46jUBHhXdCUhbp0XhnFmndy59k1jRvMbWd5D13rR3J9uTa9WlYXeyw3QLFryp54T+IWi
i3TeyguXnY7PAXTMAXvNMC9827CEDNiSLmnq6OE2mf0cUtZTFDoU34IrK5j6sY9Vchuu4HHxJ7x+
xQm+g8PDniU2TC2Ls4RLKfsv5pcpUKD5MjdxAyhT6WLf7XJZtOG/U+1AUknkSAZlNQYsL4s00vdx
Ar3nvxEjivaRgeNwL5Qbr6lkJy+8jew5VBEl7o+YBKwbNAH1vh8iY5Tr11hDqzAo76u0XJ/KJSbr
XuZgSVPSqLgMqbn8t/o9Oid5fgYd3LuyMdn+nxHYE/ig7GuucRKln3O+KUGhBZ5DQVKUFLxpzXQt
WBEdYQVZuxxtnCEQr+jDvT87PRLpKBo7O5FAtErWwv3dtSTEG2Haekj4E3nQsmgMJfwqbAds3ken
lEiL5qNBZpZVgqKbgJt9DCD5LEfr8HV6MNIIRr1MrrSEhF4xvg8vFo+4fLczRrY9hB3ZOXbMsOfA
TJgwzFnHYXhUtkgGQ8Idpp331XiD6Y7tgLfaqpmjYJ9ioe2iRdo8Emwsa7lfWbejH5nJElRyLfOb
skbl/WomdCMwWn1jpmJguPUSqj7vq19Kv7cF4/lVOKyM5IZkCfiFz+jdMeb8ElEnYPQAlajVVK+C
kQEdrBbDjB453ObMKXvfvF+s2Z8Zeoo0ZgSvbJZeFw2//KyYqJr2oCe8jpxY7XBtZxyXnrJ9Bl5k
JgimuCotUvElxUzqdnuVS55NIycM/vtvhDfj43Wq96/r4K3tqVDBV6ybYkY/j03a2A5vMhtgy57N
zdE694KFhii0PqpZlfIFhqS+5+hJJY0PD4kbaDEcrw3vUulbny4LkZK9bPLjuB8mrPlJzgKJLKSF
1nGq05U9vVLZVP4aqnxTOHOZJS6/tjwpw2rAW4COO65+r+nYQuR2MzP6UK9KiAhp+ierVpQTwUWk
o8GgA5k1GgOlAm2BvZpdbm9yu5DkMi1hr6eOQfnfsHxK3IabaxJ0Ir4PFiUVxP1BwJ6rH2xWeh0X
nmvVq6ULWc2G4EVovIPkWGx1ngyaMuIDQtkDtu/i8SRdfPBRnTpGCHceAqOQrsbOPptoHM5viBN9
bK0xGUZFIFROTsHTlHpuaJdXP8u+4yhnZGlUnE+fKnGTDG1pFGlfAdSxsTl82lcL/4mRDKaUAf5v
d+GcHo7BdxK2/S4D1hOcs0yfe73hBbek9asY4IvzGYqXcwo7qJrQ/bNtye4BxumV9DWdY7b0R/+J
R72Yx+uTjlDyak8M+2is8BatKuMaUPL/EgelRly+tmKKnCYIWFZm6mLMIULZvoSDWk6Hc3q57RiS
uAt7SJrNc495eNeFJJRDsilzx+tIkCPmww7ed8+duJx8Zu2HYiNsxMwhxMy1duTz5yfwcjIbxUVK
pgXIVljA1Nvr+j2csRT6KMUXc/XonaNlw2l4n/O9BCuV8gN+KpSFl9K/JCPEUqKOeskFCldAQ/Ur
BLLyeEhv0TuRkDgJFvQyXtvRouL7UsaQhbeCkdN2LsSqy69VnP39VFZTRP/5CAY4X7kNUZIkgo7n
tZ3xncxuRTbuh3wOymqmhvHqRvQlZG+BC+XC3OOceB9GCIu22NPXCAeO5Jyz4S+sSFXydz0fQIBg
ELlgd1Iu4ULXBhg884hjues1xnke0ZVBoeROeHZICqP3Pm5qZTw80ZR4r5w5qJWJBVgyn0Bh0cru
9xEjiu40aZpAFIgBLbBH/+sk+yxPbB428eXIliU9ldPp57ma1OlUaugfY2mbmd9kUMBLk5XPnnbh
ctii4WD5oUDPBNv8sdkIebIvHba7I/E1G09A5i1yCAbvUPSyPOdx5KlT4Q+5bipWYahNBhQk435b
Ph7vDfdCtmt51jAUmyWrNP5coyyRAYWBxmHPRZNSFWl4/2OitEAnwnYQHrZIu8KSnrk530chec1p
ZjD0fO/n5MKiQHrQEN64SsUwvDVApL8KjqUAZHzG6qrAO82F9Z8IeWLPeA2S8/o6uNo5hmcdKKY/
BYtXjYRLbeRXnm0jt8dBc4t0wJbjimOmWDC3eh3Ik3x0I075Jr0R5Fnj6sc3Hg9YHAIDPdw7ULll
r3GtHdDfvvXHW2wN4u+AdlNxnbI+5CltVuMZ9oVUAxMY6zh+DCJ/AM5ZrtGKTQNf8WYCSCorberD
4fGjSpDz2HP46TPHMpAiMNYinrBcuRPfpggIuPp3y4sm6nAWqZ2qhV6plMptQeUmuwpPQK5lvtKo
zek1htj+dk9eIwPh3ZSmUB6EG36hiU7uqEwcAeAd7I4cbWQYjQPMFKuR1D9IbDZOnW4ySZiqjOYk
I1rEwPE2pZIJVJb4F/RIgVAnxNC1vkK2yYlFDm3d/20MLT0eizoA7xx/haRRjhSNBKDBRdilMnpV
Xba3k7hrruMSjiTV7i1vVVe3AZM8gWGjxbJjZdYYGcssMmyQZUW0mjPz7B1K4/+lZSFqnUVm5Cww
AP4etAkpWdBqfkhrqyeYp4ADDdW+xJosoi+OSgm+NLGpFnBNO5R/YL6MyhBCDegJQLAp3CxpuW1l
P+KbZnZcVH+Jef6+ZypFeXlGPfkAAJnE0ubDDa48DO4QBp0emBZ8lgutjSE0DJeSWgSh6O8C964t
rAF7/fQaWkrQSPkSIKtq6N07/XnanxHnV1BchvKtcIfwwmUldm90Yx32pxwb3FME2eFsvsLCedjF
bAgyiZX2B0SrfvXT7Qmky60Iw6oo+b7Ng0l06UjK2HNGwEBTKsNIQPRMaxnuRktVRRxNN7WlIpUC
UZqDdvdhd/yRZRfkf9+bgeenGxW8dmMwj0d9DElQ3hPYCnNpg3GmPHPvlOIXF/jYMSViW5SS35tt
P2R9cDokznzjYrtjHVwkdUbQGpWcFkJCDvvRZ5djN8DL0MTUVsCYvRYyju1RGbZHer9fNabHNcAE
yGceElZp1Jxuwoi4z1Go1rJ1gzgYz6Drm/lU1HUiNqcsfloV8fL8ED2XK7Ff+OLM3EbSsr4luOFK
t0mOWFa8mtjmiK8tnsawNQSVnyjphes13/HOAgwnH8wJm1tsWYH/8ZT0x/g1scxJegc9rsJ42LOx
LBLcEgAMOW1y6W8WRBdYpaZ/pkeCPUG1ymv68FsDHmFpoyMz7OtsJ6M0Gjt7SKlXlufhZTR6o0zE
UHfE+zFFm7r5m4wzWK5oEWxoKwOCbbUxlUdxhmbQH4cJyhGbbmb5jGt4uJKOyigZp7NIWKCrqQcg
+4xfNtb0CYHoBmKFFwzZXWEl+VTxnk5ZBNhYxEVqlPUnP7Lg06hgq5WGYSYoTzOd9u2f/2p7ZMyj
f1o23DfevmAgA0ypl09JnisMViH+5AooGITxviWkYX3Pf2s6kORDPE7Zzsd9M3M4/exV/lUS
`pragma protect end_protected
