`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qA4fPvGtmqFTIZarjOkw8L7thMZHBzypIa+NzT94XdVbwgRBmLNOxZxV
bPB3BVHbr81ENtoI38UgGOZCwDb7oinYhwmz8JzL+Rip2eKwijA/UiEMuMu44bvY2NWCxIR6P+zo
1V3S+m9giJHCkl9jaDtL2tf9D5SeSiK6hj+7M06EDLVZwaTyfoFILIvweFWMRxi8WZqv3eWBeNoz
nAwP0sGWcUq535uWk4lnh0FJ0rbI5f3YBoqXxrA3TasxqKcHCM1pacrqC982Kv5vXmmJ9XiBBY79
DHL1JGBuJsODusP5mAh21Am5+1A4gO8LVY8CizggECcFVJZwfJBy8Q3TFvtTwxm3SelHB1jm6ipe
DYYYHiM7jj8rONrteeI66jf2xS8mI9dRD6h7voSAbpwcy/LorUw5G3A3gy2KPzIwEP6MA2hR1rWB
KcgpOirl4Uyj2yNHs8sVKtToa1u0gq9j8uqfT5CmBQblawgMXXN8KMYeBNBmiqIhQ+GWfMj6EFG/
HKIh5TERYHpCab38QUKChLLrZc67xdRFrWyNkhbn/BqoH5O3yl8DjJhAnnIsglOHce8oG//qrxJ6
ofWCsrvSC0R/c0UGvDyf8EVSRZeTMzwkuM1PVDF9PlHauqw/PuvMizbvI/mP3Ib6Xm/VHC1CLDnh
w1Q8dkcU7qCnA1Qqbrz/mRAAeby6HIDYHkqdLoX2iwtoEDiyrOq6bEfJuoRUUoiXYznUj3rJJ0gA
GWog0RBV5s3vqHjNfijePDTnteA8Py49b84GD08PLAuvZ5BI8ohAoT5egUuiOcbXnp5ygBJLv2bD
tR3L597byvmIVCT6B9w7YENND9g/OY+MQXfVZDKpHqEsiUXTEQVWthT4zL5Mc2K6HOtB0SEsTRft
Iwc6BI8ZtQ7L4iPYxft56YDcOR9hBQgqx0KkYDHjYADIgI3FCHJ4v1S/wLlTxjjhJXMA0TyLg+DG
0AHLh8EY7KB6nZIJ4pR25ZbQfvIppL5URRCBabaUGmQyN3JlDWVnZrA1lR+YuE0mo6TnA4fhuN2X
j7pVqk3XzQ/JTZ38H+i+Gfy2Yk+Ndg/tltD7+/L9OjMGOt1g7n94+hp64hv8kNYqGkDqGgUJi9af
RMs1+0fwkOUJX/eT8XPv0V4TY/jhTkHB277XYi1ihKaZC1TlJLXu/jrMiFZA23AcJKQGZ5Glj0OK
VjQfnM+Gv/vwmdoSO0rrbc0wlK8lnYFAyu1VYyTPH5GDqGRTIarQPpocRuGVUn+Pbuv8MB9gUB15
4lPTVomCdQ2xJRATBZL9PuDuyLCt8g7O9Dh1T/1ZT8DhJ6Di/+YrfAX755Uf7p1u5CJ19llfI8vK
0bwhUUZKexCJpCdwW8i5EoCWAR3ypXLKsOJLjSKxFC7oXhBtEjxtXCuLRdXt9vzroi0izBRD6fkZ
9ZxzKGsoZ71PBdAPbsO9Ma+KhJhsKchoDAejsTZTjdBIiSUpopsuZ/+TeQy6gUMTpQQZ1EopEwsa
Ug+CADqUtvh2yZ/ds9b2uDm1/brAaeNgbZ1FenfPaxy0YerBYiRsnymk8UA8KPFAc7jSaLSTYTXa
lbknD7m9yAQFDWss2gOcku3gBnhP8N2pHv84VeKXytLEhilkPlyDHULg1qkOTrud1AV7RjqSVCsO
bzxaS0Vu7bbytqoVWJ9vjPea6Cnf92JUzufHSN3sFxwgLfrdCVXkyTrRfof9W1ZvgZqGuXj1xg1F
z150BpkisrWVLgEZ4OXPQ15I/RavTQceg9HHuLLd56Xrp+7VHLSYQxoZQGBc83M26bOZKIijJNkj
VmJQ5rw36dx5J5u5891fXJbt2XhWxnlACZnJyQGpsGkL/HrKTEleqALcL5CKg5DELjmXPPRVvuc6
ZuRp/5nI3aKDZ4mv9AEph1Omhn+rvrYXixDz+T8McD2hh67kaqp+lCUbm0Cb0hnA12ADr+7u5dl7
sBNyXS2gR+6OcJePPw5w21HMk8AOcobnwqSGqGUUrOiufx/8VtSn1Ibp7jgU5xSHHOoQDLjKlER3
6zkAzm9Q4wizUbwFSnX7FS9f1qOIoyagUHjGejE=
`pragma protect end_protected
