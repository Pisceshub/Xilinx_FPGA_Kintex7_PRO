`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
KknvL6SYSb5dRFuWP4AJqBhO3b64YXO1jXJrKEg0Z3ikGAO3obMtU40YwJiJW7ipQ08/Y8WRYNWh
nV2LdqH0dA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QLUbVPatcj7IWeOM7GaVpOxxKXKrfEAPdOAPmfRnpcapAKHnvWUhcysRYZ/rY/73FKWInR8HJilV
JFgxROZVCNWQ1zJhGgmKt04WHahOu9miHsfm8H7yNJ6k3TsDqjbc8beG5UCVgF6x/gDB8LRb2Vlo
OYeUOl3UjHyll8Sbd9I=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4fDulW+j2qCXqz735RjXksliYlPtal97cQEPC5accAQtxDw7TbdSqrHOiG5KctOIuaRzvRMOO5x
8R7f4K2bkMvIUjiiFP5Xw/fjJySLFuOiZoiNxxNdz5n6QQgBWYDepruKbEU7yj9zlmf0zEFmWZo2
ShS1WpLwP3B9Mcm5hJ+0GZ0wSeVmrvJEKp8kqO3uW6EVpKbiSMmBugVkGUzz9ZrIbzEZlELi+wJ/
HVgQM4hNwGKaRhAKNMJGLkgs6Mi/pI+CqjdrjRYK0X20OxPYi7+y3i6gUy//rkWJVRVSqqxJt07h
XfBm/2egXCeHNQMVyg/cuW80bFPZUcKb/tb28A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eEHF/HRqboErONr15dWGPiKIhHmEp89NzpKM1HVNOPxPMAhm5Q7SHcs30Gyp606YzPvXAWOwIhp6
yShxWJQDMNzjx8XLNdk6Hk4q1OFOlxJvftzg6IwFePhX6CX5M/h6gWDjhSncOnYuNt1s46FrBJGA
DJZ7AbtD39aEQbpRrtRqPKdh74/RGoSXOsksuOHq//+3LZGY5WN1wdVNJTew5IKMLtb98TYlHOO4
w28CobD4NywkdWMYWBeN1weCfLySyzftQavfk/dRUoBAG4mBbSm67pDUnjTuzD/BMIiEezbjKgGt
v5JKng8K28aaFylCDbrjWbQ4f0E0MG89P9bqcQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LBodvKMdQLsL3NITg6iyfn6uEr0nsFsSECbcpJ0VM9GPtNyhu1PCIqop74QUK0jX7gNod2kXTA0j
UPAVU1VbFsW+W9odvoIvVhgiIvptX2ncKxVnQVrYamDTZTPdFxs85ZcmhfukKF1ctZJMx5QHtsT8
/fgDo9EnaiAwUK6EH1vPn8nlJtMakUlaKARMU1hnWHBUkjruM2J062f3fYCx1Fc0yI51VXZXtNw2
A35SpeR68WKPmXnaWtRfYcT55OhdStBuASxbBHMItu7IQi56vUWP8LJm5L8r7e0VPvAGmJGTHM8m
DRb2QSYwaQDB32Ac/WNT/HueDTeVlvRT+cXLnQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RTdH2QVRkLMNeDjWHM39MNQI9JpZeMEnnaFqgJIEgBuj3R1/oXRV+h+0yVRQ+SMug8jz9no0jCSS
W3wRM89ooYAXiOYt8RwiQibqZKat+R7T7m3thhmgMEI8uoi9fGuXrcwO/YAOvNwNOuRc5iytwydq
EbyW4aM2m+CrXKFlD7s=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hNd+z0nXH9GYvgjnhDJoJvhFhK8AT6oUoCmTuJoXrdeSPSICu0d2AmfE/9zKTVob1byyZNQ+dZJb
Ma+7SxXV1+3xFvececBxzrOjVMq4geH8T4yeo12KR/tsEogGtiBVtNuwOoiOTxmMqj4v1JDOa2o8
G9PU/lTBUSoEzibdcIpQyhvP7Mdz6AOWlVWthHuCNvffk52oBkFkYg/wxqRli9uZ+ljnrd6rXIeN
pcjEkI9ALbBEAZnGGMY3do4kdn+d4UrzbiC/0FwIrw+uZYeWK2+A1bCZ3JcBMczd2lYYJYQOACWj
1dr/Sij9Dnl2NTdY6Acp6dQAwn2oASr3Hs8Onw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34816)
`pragma protect data_block
F4D6nIAHG9w7CzDjTOGl41ogLfBDzmuspYZSQk8qjBrLD+fuS/xoVmRkiRkfH8qXh1Nnpil33Knn
UlObw7crj+3qf719zum2Fb4AOKQ9JKcMAFJNKzEIVNEjdvwXnTmBu3rn0djiLJvCAn/zy1iPIEiY
AfPF8PrcM45vyytd65I61LkP96RToAc1Vv7kj6kdklaSjCzuYveZwiJYnUS7l2NnMb70thBaG/8A
5sPC7zQ97HJO4j86NrXEpIq753vfHyEho1eXmloH1z+XBOPiq6HImTmpM8GcLj5XcIj7YL8iqboi
4fyL09nvq///giq3etpvYe7L0pbPFMP7ERKT665SWCCsvT1c1EpzwOEcR0U1p8Xazc93eLDwhU+y
iyyYBxc3NVQw9pGnds7MsR9Fc9u5d8FpnwKpKF7FYbhbzWw/Iywwr7VW0VpUBuwaJuCuOfiOIIpB
97E6yH7DdPtRmeanp9+iLSbbeGQUnpsFhcdPvtEWkIfIiA0oD/etQSH26plAuV4Xs8UdVIm7odwI
d6gD2xmbSsxxvb64zxqXOcrZm32FbLUBvQRV05w7Yqg1TvL1E/6JHFie0taZHpaza6y1cVqzOKEJ
4iR19bamoBK2X6OUsI64FD26dqadyWcxFuJHYKbW4s1WOksOiTfc/Tx3Y+BRUxZuFUmsltuqTypH
/JTXm60VWQJGmVHkbFZawvjMK8A3zO5aySkeK1ZYogAAHtFS599ZgJ/YTjaht0P/BYkq+pt7OLzw
69I3vBHZJJizmjvN9TIh0U2Y0QdSVkYQWakNErpAfPJTzESBE/kFZxZ1/F4IZnQIOwJVO1OnCpU7
FOnDXRk9MygDpjCIyizjHuAICfacMGY0EGrOVaiCqkkeTLuGVu6k2XnQEwnV8OrBT+09dVkCIt+h
oWA93g25nO1naESA6kJrhqEHjvyIdUyFvYqptm/zIPZjFST9G8Bx3ST8wb2VmUKwokCfZ+Jagj2j
dZ54DMjYcb0yHpfpieH/Jm7b1Oc/wN8Gn4gzMM+Y/P0zBhPpVu/Kf7N4t0SbG8TLyzUfHnhopJtG
fDrIK9YR+b3HZ3gknwrdcWWLuEsoG2r4IbkHLvQnXNzySedamwy84iJ5p8nFZfALD67mXGgWRgIZ
gffmTagml1rliSAF+i18xxLfHzqlKeGfPyyC8eptxT21WPmcceCHgOh0vI6gGkjAKJOScVyLTls5
h66dg4UaW4x0e1RVZ4cyUFcfLx64C2yOpJVAHwryyFeiwcSMBetwa94qoj23vB/5//ige3GZIo/Q
r40Ylb82xqeywa04WUZ3qnGa6hFXKn6I1QlKLdHgDMFdpTLZymd//nmM6buvz9iY+0rNQDj7Csjc
nFxV6cERu25lLNf7QT+tvxH673GEhMGITZboUP9OIAdfaF+42rSwvhaeXnzRcmpdjfXseJRfVBLj
79VezdE6HWGKh2uo8hMnmhJFCdsToSTSr1tEUvl9B6PN/AFZR5R6jpf3hvVdB0mZbAPMtrWHYhh3
0yAXfFrvrxGDt257GyLEFkgaf0ZqhEFb0TvsWqqwnU9NpsRNllrV29tvYA4HT75gvoVCx4W186sU
ppniYx6vQGT37SsaqLb6QmbIvlXQcA/x69n/2Mp+88xpa2ZO2rFnsP+S8YalYsW0K2JqOVlKB3Qu
RWIeeYmp+cW/Vk7Rk1tty1FX2n/ZwKigcyqcNP2kh/jVzHE2UkHV9EkU+SGYohjmXGwvGM6UseuO
jTpwlpI2W/FIq+hz4eWlObH1mR2+4gem5jar0GIrFdI+CFDIZAJHsBMFakbmI3Js5UJ8wwOmgKN/
5aPOXARwM26GU5/Dz+YIqSdrt3zdw7K17YRKqkFgEyeFwfqAUYlVv8GDmVztueq/weVUW4ka+vin
K5YJLJufZwSJgSuofd2WK3nJT/9M2tiT+OCufeX4sr8XZK1a+F6OKk4PdXCvP5WKyVeZLUDizq1V
32EI6TdBAS8CF2u2xe38mcBafYwOo2Xi9Gf97B3KRtXyINMzYLwdUv2zpAcxXS90qpM36vmPDDM/
OQOWEkOiDf2El0kAe3TvsPyYO0ScawnrAAJAx+fbJufceO3Q8Vn7ekivdWetRI16zWXlj/nfbO/A
L4To6F0H32fSguuSslxV6Zq7wqzTAYXDoHOEfo0E2DKpPe5q8HRw+/ICpg1a0ehfULxiuX3n20xD
mxH/2cByZoGre5fqFoHVn575hMyhpjJrBFjO++dZCwM8Jk5x+6ir6h29xbdxzRJqdXi3zhFmPUax
VAy069c3FKaqaFz0U5vdefQOFu+lwdEaW0B0uTs10pbRzQKGQ6WVRvcu+BcUAuhJlBvlrsWirGGF
fIBwqg/wfsfYFTkuo1I23zxXOndUuaciZ3wYj2ZtXtrb99b/pnuX86PkhHqt43hzTAnAR9nTxEWR
jF75Pbg1iRyOTVScIqE2YJzssi+2ve08/frCc1+KSAZkaIp6vRAjOQajZ6gjeCHThMsTGV7Ssv9c
/J0nNP01qwpwulTRRq1uwHX60Dj2EWP+ETpuTKRvRzel1x31zo6knday1+hNOw6Tb+ZKNTNJ/8gI
+0qNrCyglVZYCAFLmLSC+R9b7cBja30khkliVxfpzlRRAgZ4cZf5LThdg65RbGSW8FusaoHSvUHw
yEe7vxnBNhVgbLUknZfDotO+U/bKP2ovbeAhXMHycjrstDtwnsZccvYjaSXEZfAo32yclAxKU9XV
tVDdhtnMyw0FNWQbDiS5g18tpbpKh7YkOtYwM2Z7l6YtZWqImb1gq3GjJ8m+DivaJVnYdx45hABY
51hOf5/YCAuifT211Av8RJ8+7WaR4qa14GdVGSlugV9AxyDJFsWrFZHn1Gv7TZ0S7Rn8eULYwWzi
SXLr1dElwlqnbX4dE8t7bF234aKI0NsHpIeQPN6lI10XYHRnz1WoMXL//N57GC/orGyowHaZ6Cbg
FICpgwjtk+qbsuO5Ofy91ohOembjwitTpbzczkMP7M4S+vJapkj9Sd9AWJhPKZyhxVKHnre0vlxd
uDFPhXot9zMcNKqXDjDNg7lrBVMJ1DCe6Pv1XPvmdZ9ibdbX8FVroBNnvuzt2NqX852vOmqgLrVT
wxuJW8t41MlhaYmNyG2XT79zSzuPATsZn4ra3PrVlHNlHMe5rL+woweOPKwLNRq+ILs9xstiVl4T
q7Dp2lQ/dy+Xvraa/K6koQF01OCRSnxnfnuSr8tsAx2GZ6bGBgFBDu5oJ/qW6fF6ObCcx7ubrWqC
y7QxtIrrrQLP1K3qgCOu5jZPGi+fARiG5RPK7BgFwEWmiYDv5y59wb2djPMcGT+q/+EurT2+sANN
h7Ysb8ypU3P9ONlwGZwDuhddCZiFv+474NvjlY8ienVv4yx2D7VpfpvEeY78aXhDCHSBRGb9Exur
V7gLOyQwlHYbKsUU+taDsnE4OekRq69+o9JEPSHXkHfnnWePOJVhPLGpl1VEjUXBce6TBV8iThZz
xrlUc110tELuUkDqrc2zSk+GenG/92qt8xUDTxal2U+DY2ofiCk2UkHP78ni8bACIAEJct07G+1b
g7i73ekEoix474z4/gX0Pj3CknftI+lH0qWKrGV1YontDsXiT1Nb0LG/ex3sVzIaTouxgJdKsofG
QVTY/fwp9L7VUdIu33kbHcMB98pnOyu6iFYLxe6nZr1faUNEzgOom+Am7/LQtQaGQYGG21IYejwD
BJIw77D0s+u5Pf0VX3zDEkrrzNU3q++wG6zNlpPn+KwpwOfOm2Ucv1WUvPWH7nJufecg/92PgRLG
ETmHn7MLEEteD8a9n1sX7W2PulIPTAxjfROVfZPbCdHmOEGp6qUKqtdlA1Wbmy13M2EPQZZ2b5Yq
r1w+SfcXjAGW0nq2QTetv7vUZNcmNCTwOGGQTQ8OKNfktaT37hBr0oSBEhAlRroWP0Zx9Ywx/rsI
UeKmNu+5j1XZS7I/whmThBORhhy+rcqG2Ew3MWZLKW3QYP9lo+2b+cBFKFy/hL3UJ9Lwfk4RUOeF
2JWCCQglSFi+TrDf37SJQz8U5rAPZVrY5SfdyC5fvr32LtNhRRDhdPfsk7glKGovsnYxYik0//tb
6JxEtGOZrOZ6EsS6lvW9bzfh5h8qTpFE44AZrH5H4Z2+T7WVXed+cLbrEew4O0+3ZaJbeU7qg+ZP
pVbbseMeeVbr5j9PyiPv60mmXsQjpIG9NV8JcKIzTV1PeFkLkc26zr/yLkUpVMthjFt0REKxG1Ay
dqsKGytfmx6Xe9rgaUmQ7R/NsND3QjJVWoCWPkMlyl1BfMMA1nKsnA5kdoXyPGPXaDIEac6cHLLU
nRFDh7pIVtFPfZ652YgtBuIoBm2P9G6CKSxJ8uq+L1dszyuVsipCANr2xqsWCGFsPdXGVtDGMYbf
CvY0SZ6KVkuujnol9qP+uIzlYXgeO75yr9mDqATl1HrIVovDd75IXJiJg7viX2+wRGBSvbo6yFI8
oLvS67W6WCs9n2Qk1AacxEE7qMAt7TjedaLmTFCGwcKqead6xYzVDaXedqtuTejZDJc0LIEmKMAj
z/z5RgHEkZpQQWCvL9CTAVw1/iszqBGEV0TjthNhCNYYHrxUzpqi2xtXVau52lxtWkak1v0ShPUM
epa8WM6ar0U4AGeK2g7XYw3tAxFKYok6IGhrka+ipp3x7yTqhUTJrTsRbZ/wvdPaXtmSXzXYpmIz
gtCxU7dR+Q/YcPz/KOYtZDv7Le1HEa9tZJwgEGoOQMfPa+NYS0IZLLIkmmN8UBIj27hazS1DGXvc
wX00eU0R8/GIyYobHfoXB1Zp+pzRMrTYzq6R8MR94DRR2wM5OiXDHkWcZE934nJlTIagy/o10SUL
FmSfAJcudifG70Pv2WQJyf31a2J2pWppRVCg+F4FE8vf8vCPJZwuz8N2wlfmfBYstq+FVSPE5Boy
0p9enVbpYUWGcrL8xc7kYcf9ioQ1FJt+GGxd70bGFZHwoOuee4HKsfQsn+QHo1FojTp2fYQsP/tQ
Ca7//fr/DXxlNfomBxDskth90DaBozr4pvBlxhvIKUFpoGgjHF6D8n5h6RWg3COF9W65iGOGqXVu
1f/ToBVSFh6QYEwtrmw7JVPHVb1/mJOAbMdZRMs1rojwGRBTpymIOzpJU8TIB1UP4llX72oc5VEY
/f2lpCoRoW5zhpIkazfByi8STb9wMO48mILaJElylNmff2miL3TaWCxkobSY6ZweaCICGjJI0Nno
dCVa0EW8+lyM/Tue3kwepWugSp1Lb/wJpOUp9An5JUSx/rSXeqez/kECEvjCKM6JHUZRuFUz7oPD
yEfT6zNi1WZWtZ5SdrnE7UwT6KsxLhVksNn2tBU+iXfusfbMVdwmvMtlqTUw9Se8T0Wzoi75/Ipr
CekiIDWLgoPFn8m8Zh2JpSsO/XRh/y2xuYW6FVqxt4VGdgJ7DZ4TQwL/dYf0SgsZBmBDvAyjKHWh
z+9iNEWY8DBXppssOJCUaPxyoiITJSR11CWgZ+I9aAODwWxZswQ7+yntjTYBQJib+bVS4j6N67HR
MsRWR3zk+CdlNuZJWFg85KGO5nbF9rIZZ8rWb87J/8r/CZMR/8+XTxLQooFtLAoylWczKTVxM/xH
+4LyApdECH87oXymF23ykWw9J1e8mfx4MprZkmzufyCYFrDYzbSng2N2zV5rHX0R0N+1P13BVuAi
iAifw26Odl4A7m1ZMfs8pEOCznrZwHu/FcjXWeR/dBuLy6qbiGX3ZcooN4epTwlSMFIOq8+L0Xhx
mSoWJCKXYweTD4Sf5tiuBmH8agMJlcRNRbdGnLo+HVgxD0ZmMDcYUxnyC2tp0neiIVekmINWqpsg
grc0E7Xcr1/S5Ox7bVyC5k1CjAb5t6/OqVz0T6eZ+xqzLRqWdHE7H4FWtolWbt2TQn3lW22TJMIi
na8Hzvl9Rm8MKYYpamLKdZXMorjGputrD8zbgyG5vGAY0vIIJ24XQhVt7SD+udzS2SegVSyfP5HP
Hv38kiM6YSKGjAJouf+9fITvKFNh1Wsre+ulsHKNHndfOEE8mWL+ZP6SOzj2DlRqVZ21TyPI+s1y
M12GLUXhFf8orNbBiZxJP5AuzfV/wdZP2KOuYm0AqBuitqpLscxc28/T+VatLS8Pb2dWu4NgcSlJ
jBLHKJA502fmVaAiWYkFdYUi7hmPXwxqYyLacSwizXsbnEbecdXIyOVfG84ULglM0pGd+8C/ik07
Nmn3DpQ6bRtBjvIgYPkSZTm0LNXptq6f7XowGVd1aVQJwLTJKZ/t2XPxtFk75N6yYPGx8ZldvE5o
a4qAExHrJWvWm/8YsCcyCeH3MoviBRwd6q/OF5SHNjwGO/VZdyadd30wi9oUEISsnYmdpT+tGzSy
1CRxGisKQl67CXyf25l2BfU5Q3s9Gp07zXzRD0zp2h6g6LN3frZZv26Wq4SPFU5zpKfcJh3YsUJz
tKxgUXIaJ/7pqp9LIBF1Z7uyrETMG9eQuT+8PQASePaxu2sA/jLNTaLu4+/0QqQ71Uzml+8L3L/y
iXqQCTgNV/OdeQmLxsF6Tit1Bt8VWO/v4QQwEga+PPKJC1XPymIgJDarnwiugkSq6HUNemCft4WA
EDl/ejAnuAKuI9YwjMmt7PFAzId6fgTwEflm8D9L/qvF/R7VQOIkaNJogW5j8PiWR0wbWl18gEeG
tSS/OXg+m1NBGTvXt4hf3FZdt4tcg22fRdIZh6/1HIiohEyq1+k8p1RSmnfmC+5Q623nU3iyz4RZ
WWTa1hZyLT7HMTRjiqU6nvUXJS78stPbML8gqF3LTXRZ/j3SuA5Qv/vf3541VD1LgOTrDRetzLVs
Q9W/XvexN6L1+/OF7JcWRjeznO7GrxVB6ZM1L++zROOpttyQi2jtfZfg1aV9vVCLls5QyRxvUWm5
D5QSh1B3aZa78MQy0rtg++4Pc0OTTSxtQNo6PPShF5Ot0ouX3ipflu3A2WnwDNuFth3VriY4VeGQ
uiT7ohLdl9kIiYoA6VSuNqYEmYF94ssB3iwVSpN+9EUI7SiuioePN+icdAj4Vp0eY+LWKUcq7MN8
BC21GpwFWl67192qbHfxskdbebuD9oqVnx+9rgDuXJ6PNLYNyQkNZyGEjlsTrAP3wwPNrTx8kRTU
VdFzAXdQpRgGX4ctNu7A5LqdocGlDvp/87/2MoY3AUZhpcaEeSOHMh1LUKjZOqY8KyWJ43JwN/j+
1jMbe8FbvzIewwIH66vCTxotsC9v10Z/0AFTQQwLIg7FTX8Uy9hpX7PaHE+5gun8icISasw9h9Vu
7Z4Yp3WLs8MJwXqonruFHmSGLR444VJOTSBJXXc2uVSwJfruYcVXqXlxews+JYrqYhngdst9xBsY
SB59eXqX9NiSpSH6R1FV6MyZUWUEMRNm1ogJWaW3k0Gai5F16pl0wNyD57Xrn0oigOFs9tbOafeB
GPIvjVxDSh0xExa/lMC3PoqQIC5amV3b6/8M21qwQh89LsIiGmole9cUkLbAAqGAZFHHsvRK8Lzv
DwnvZjlpX06E0UfuPL0G+nDJ4elrL1EaYuA9bPeFysDFFTAXnFa9o9u58X+4kkmuJL0quFLqkHys
xlPQksy5J5fgeW5WF1JJUdjHo/1kMG7Zc+RXa6Qaqir1xbpHY6RJ0bCxOCj5YpPYE32AJV1xw0gB
gW8X+FZ9m5ON0L+y8Tbc5cgemDU+vBW3edBPxtzdz3y/yU72lAWyecI9NLaqyikbghIyWvIgL6Lp
Lg95ucYYEpa9BLFIGPb8CyHHwbrlLg2hPpZa8X9TE3foVD73XDpkKN8stGJGqTLX4FT275g6DmAB
thWIxqqO/O21fq6lKlMBVWtgoAKAiBl/q87nz2AvjNKdGCC6UWcvFO8kYd96MqwgJYs3OEE2kmOP
QTcXgbiCvEj4T5gJKMDU4qQ93sGEEc/m9ApweScMfuY/Am7Ohss8LiNUkuhNmPW2G10IZC22YHXM
g37g3/JOWj33LMFFMS+/3e5Ztih201Gbhj88Y1uy1fEnSQJJBGMJPSWF1qD7LtTkgsgeVfJCBkmv
evvl1FcU9LiId3SZbtvC7N9fgiYXrtdxjyVMVTmLlrdnKphtGPTRHjd2uUlnafYvLACvhpdTH3ln
kIKXm5B8bCF/KxcQbC4W6BvZUYp7N1GTO3Oo4B/oxPBDvewwB+qgo28XvFopJu+vhc9CrWWwekfx
XNPS73mMiSMV3cOhAIuROuq2KKVAHURlST6SJc8EwYTpV/cJzZHpgxpzEBuhgpONn/kEp92TP8A1
E07UZQZJDvHZ/0j4mLQJmIMX9x0HZztHQ3ikrvrJFbv+45oh5KZLpjf3dRuHAWzB4tvHQ832Z1cB
+d+s/3/nmPdggL5jhmsqCCOjFSKnfsq23RpWgKB4I49LmMA7AOd6bzfJ//L+g4GzFYxbPHpkHjJt
/eCHrEv160EzfQSl/DxaObFGvwHIh0Cf67zyyHOzplz5OYXEr/oMM6O9DDL73FdoY6A46Gqr6y+b
OS7WkVyjFq2rWqvhS5V30IGW3LlQRIg/WsDFTR1Mehm13Vims3xX6wv3+9XQfaW+24ajJILw9ji6
NPbw4fLTi9P/pFQkLx/CDKiPbbGehXYF8tJaXZ7St3EpccI2OTpS2BkkBNXVh9utYwpA6yrtb3db
frO8eG+dzzmuyMVFFM1mj42VaYKMzU/djFP9RbG1hqD6VER1fAsGQ8PncgZH3KcUVcD+WI7g2UBU
1FH9/DK89GNZ8p/KJA6484eTsot8yHelGqF8CqvXwvx/tuUGUrKuG0foN71F8FAHtv+s7wTyo+0s
19ao+S6xAYrDQ8v5w8GQmSEJRCRFLzal67XONoZitl7qPegO+ViyO8Qz64hc2rmzlbe2UA0RqOOO
004NfyY3NVhkSDNBRZ5GmTpEOSbfpXbDu+jFFyYXrR/8e3rnGojUS70TWAccVAfY1SFVUBEXbMcf
JHBMAPjrf20fGCfF+k0QPUhJlyFoYoqkdeKskT3rV6qy9rTaj+l3DMbYAPkR89jZO39GVVViqzRz
HSoGJN70x2V4Zmy6VBNGyPyEvp9oeShr1dPgzjrP5Cg8+xy6b8MdpW+FyIXAV6VUQRFD62c9lOQt
TXfB/qDZtNvhhp6b9mhW3yCflxjlYrR89PFEUHbdsZ9qSw/jwP0YvOfN1lvidGC01G9bVxBr/W2D
lRvfg8YkmapBn4wF9BYu5+V5DJVzBkuQUyOa9liu5OOeZmRAR5U8DGskWX1EBJ/JovqDsG8t5bp4
YmktKVcrRnUrkjsKRwhmzGUlYMppH4ksHwPbtN4JDyWFql/wiy5wHvV0jmZSYRmLDRHUHQcztg9v
Hgjgel9RjPezV0Csh91hTFIf5FRM8oqg7lJBLPvSM7qvhbCMZFBaMbNVxUMCE2mm58t5QL65M0YP
X2/7L1njfLa2DrESbUQx1UXjXcIPsnBCDZ5GwBuho1JU6GPcqo/bqQ9qRt9jr6bDDa4n371senKH
JpYQpnpRKCWj2t1wQ3pnHI6Jxq8qaVHa752ENx6yAZSxWw/b+4ek5H+kWv3Tx3s45C639x3GAIOH
dWCqmBtfPn7xafNSTIiFZ5s9P0RLpGsLQHAr4DJ2te1KrF5Htm84kZbrovs9RF7+B2/EaFJzBCab
5L413zNP35GMyaDldZZQIuK2uYKq+ADiLvdY9y43jPrgQ0PATN3t7w2CoQBhtUeMdlOnX7FLA+m3
qp6Nl2+f553XpgWmjeI0w0pvqgTXjeqLe24C7NunSI24tuzO0RBEU22io9ZxJ3t5k5mOWtcowKen
3xVw6X8VRp8/AlL5xgQAuVAOjUSR+7V9Ni6NHtbrmujn7u8K22mPDl6aeiKpzrrL/nEo/1UGdgKp
tIfdCb9wfmvXs/aSqkmAO2pDwu07hKT0ChPZyXIqX5+51glwkL7WfukaEG2FjtuDNFxQ1bwncyig
e/G4pU9p8/jotfCI+ogs5GAVUUNk7QmU8TpQAYQ+buzqU40alXtYJ9jOGJb5u/QnDpTSBmlUrpyp
TwJOxBO/QbpN+cBwXWWCi/GtfmzIw0En6pfnc4Doe5RlenLtjopCUTmmlAhx+ce7L2QqUXhshm49
/VD4XIFpg3wiGWcN8ckpspVd394MngTkaX6DF6S3x42JWU0qyYqCGwrviEhhZteQff6vE961tvVm
YSrbNHiwI+xrpJUR9HvsaT4T3wQpGEG3s00a0VviJBkzSpWw8OIgknSREHfpWsWZMjzsg1Eg2+kf
nF3+1GeeUoZmR2t/JuRzqnaLR3dehP+V2WWQJqNjXkWmGumPBPr4IeAYedPH/Viip2Gc1RyOHEgi
cotiprT58YpAgriznl16bAsx8A+jLSkyl2itY0VNeGTV7Z3kkP3l9VaC3YKwjbaFf8BMD5LwdT9a
vdTW44MIFP4RFImhSHgGyW/wfa/9rqAlqkFSQbqYTV2KgztEaaoh/qTCKE8Y/fWerezcoAfaR+fw
LUIpt3UNf1vDCGrGcaPelcftxxiBpMcvI468w5bg8Bvp7tZAHOR/qs24ca6fuNBFkkHuciy/fxYt
9+sy/GoQwU3XRDKFyuowwEK4+xjcj8C7KEPLwDJIoVO+FbKG3N4wgahh0Xm+j21jTKPV9n8s80jC
JpKz6S/YiRpntaFaanbQhTO63Dg7/4MoXYiNZIOPLWp4tDVva36A0Yaqh6veJnKxu1qyW7XLdtly
/4VA+W0C0qW0KP6MRc6YJRRU1wZOW9XnwytRy5hmLuX5I7bMuxaeGzsSiDUuk0fsG8mhEEjs4pcu
tGjPjr5m0F+hxEVJGpkLQT5qI7JPOWkVa7x7hsMiNq70gpnirmxOdsLtXEsu4g0hVaK5vdacMQy0
QVhQY8W0bpqpTaZ16SjkVto7oAP2sIRt0HwtAU44vEaJM4MZZGky1IosMCTBmq/7Q6u7yuwI1Ros
t5QbHZ2uKm54UigA2m36o/xKcZfB5fuzXeCKxPymkIw+DE5GfVMrxuCBBjmmA2HHhIyQPI1fqJ6t
oSQzfJSnVWUQuhNN1zyfWCGv/Dgs+o9vypIRBH2QCHeVntH4iVIbBjq+ymAHxOHSJraRtZnWIbtm
t2eRWUrxBC9tyuOrXkqtSIuHOxPwi0h+4F3OpQ8oMuNbSkm3g3R8tG/9eP0WZCTklUi6W0lDubov
4Onpf+tZQUvwj52EhA7MG9nDFNywFZ/bB0tCOmiJTxCZlo1gYVKpIpbRFuxr+o8N27UZ5HzfD4lJ
0w+YzWeqWxbJ1kmCokndyhhwfnshcu3SUSp91XGFDUdpEzy0T7mRfZD3W99dirRBow0X0E5MQdAe
scJemX1YBEAhZeV9waKgiPjQ26KBOA7ZERJDAiqctk8RRtvxz2cFO0tsWVTL/PqEMCg3drgvTJ60
qr2iID4rhETtsvXve158JUWtpX3Lb3VNMwLhc1pKWayCXke0FytWFWIZGC0qoY80kWGxE024IKML
Y0pVN9tcW6uofSe14vri0nz0Ogtqsvi2lhRWQLNDzgAoXgNB+cB8M0RA4VwCM/V+fhwZOmFdosLR
4HTgeiVMij6/HG2IqYa0Scz0S+rNJ8ioQpGg/7nZ6/27vt/Bvnbpe0sLphtRrZq7/eUqdpRz82ya
pUt1YbLwi5OkN9jpjT9uAiDl9T9atVd7BzODv74eyKYQe686DHYQ4WFTMElPKDY6MLgxceS9IHcS
CtI5PeP47iVXY2HCOgJtVkVvIy+JRjtMlLcXHR7DByPMyZ1HDJqM0v8h8/syGTQYZYfVRKzrY1Yt
7JscAJ9eQ/29LX/wQ6lgO/EbODxsQpisOdNhelCOoCyDz5OFwOK+OJue2wvNtp2405uIn3wNU+Yb
144tFgKGDbUZKdisVze5Jm9teBEqHxk6VtlFa/9tz9mMwLgomvo8hlMhWs0GZgLcodgKqhBJSpm2
5PS9FqWI/yOE+/smn8MdLEGACYdBa6ZmfI94/jBo2FoXXaR9qqJFTMsL0gvZHXKT9z/CmA020LtP
UvxR/lpw97WkQRKI6GA1CHstelorAwUzOVWq/TNGfyel8kTBuAskktncODqS6YkNC7vNM0+jpQ8y
0fOmULQY92LdUQtfzEWi+YM5PN1sSB7wuRfQ23ZlZiOE5h3PXa2UawtyxSPeHCn77/SrY2Wq1GRj
EYktkPQQtcTY9tmmBPLCrGbuilBrr5CjZHzGz7+BesOEkzYK/xkt0FcIARzzV2L9199ax2IXLlOs
lN7QCTzgmCrRmJdUiiRG9ORrJbiYBP+QWIAmWulI3Q1tGz8m3IA8rF3DjGyM+6x2mJIz6Int019G
KZJ7o7dXysStVVNGc67qi/rGIFwIhr32DuXDmbFMmciBPOsYIrr8bh8fVdQh9PRha8Y1L/aFjS61
55rawxWYEDIGi5lBX8aOGVIAf0AmK0Q1BXMWmrNqCvmdo3Cv/sxqFjXPuf7Tq2XrWFF8PNgir2Oy
4uYLBvj2NqH6vqCnMJX5+ejJ3urnapnFTROzM5XzhKNvghYHiHGeM45dnWuKF7x6ErJp6HOQLZkg
5vSAKaNtyAiE6sFngcE81pg7kEw9rB7DJIwHr8OHxN73iGY5wi74MijoUcZN9Wj0cRbGT/xR3uLN
a7IdKp8Ny87bYup8N6X0lhL7Y8oUA+UZYb9oibUiRrDZFKoPYf2BbnxuyilzhmrCvw3swfe6Q5Pw
s65wZY103mnLZBBFqQ6JoaSvdWfZbt/eux1epa2sIb84+Tv+nvchJw6UwIug/fdr6Ze1WXoQpJhN
nwAWZRuK2t3TiJuJTw615qnW2DQe2/84VhDMBcx/Vp60fcYngX+AvKUyXXCrJ8+uKDkb4iNJQfUQ
7Uz0O2U/Z7C+ykJ4prb+N1WhaPwERbdYUM5Rmfim+EHnm3xR+B4z1p1Q8iTsQySF/kmvFtLdd46t
m339g3zqkM7dVepwx2Dwaah1vemOiE2uZqs3GOO5xUWFlij8hn0u9AMBAS/iQl5p2NjhCXOXs+Qr
c5C07cSqt6wtZ65tqPN2SAusF5bTZVAOnzE8bkD21c3y/i06p4DBpIchjci/Xw/UynuykxIijFwo
pl8OsXge+UbJjIlM+PE5gG1C2ZrkXGCvMsuMJWu/stJ+i0l32N7DlGM+IqM0M+n/yyGWLYbJwncK
/ivrtRu/N0M0BO3aoaqGbnNe4+uVoWl6gkHoEOLWLDjbMYvTC6WphE0HoWUscnT36CC5ODwGOsj6
8MFg6Qb6aNf/tweT5wTUmE3VCgIIB9Lfscb6qaflyJ0ryBITtH8Cb9SNbOHnzoaPyEbFvOI2X481
gvX6d4EfY/oWkUMcZPQcA8SUO8oRBAxvi1OIXudd4fuKQpRdWmTCESRqxm2uksysMBorsDWG+J7x
f/BbGrzgtv1a0fSU0Vp/mWjPm4qOKzoC7qWrxW1C2Gag9xTthbZlqhN9D8WogyqsbLNlEIDwYsEv
qGZjxk2a/oCZpFx9qdHDryDsBntX21CDgo0pXA7CaJwQ5ekoivzAGnVzaJGvnIw/SSJUHBk5Zl0e
sjIareY6qozEB1fqknxSyX3My9EpCXa/28iiFD+/Y6NhH5DxLU4VAKgpvd+RQ29CWZRJjS3as8a0
RZKTrjx3U5AXXgsfJvuALJm5Oq8rnLyzecta7jDI06mqvS3k7rB7a54oHmitDcpAs5BaUQIcAddy
/qVPQR+hgU6h9ZmFAtKZSyAu6ThXtJRYkNt5d3hZmsjGmeA94L8nuWnjQbTQlTEw+NEUPkp9vsvP
raSAWdYZHW9OmRZCSBl+YTcYhAKv99EUhPejXPEZ6N0gwG4UwOICi2l4wkJ6uqzsXXFHn/IZziY1
OwmK7zkZTOzv9O9dWdlpKNgKraep4g/zVFkI2GpYPASJjqfF95Yvcqh+O60qHY5eV567QgzlHc5h
QOmjB9zSwVI8Niuq8hO/6aIwQodEvC2q1sXB3mgTmAjkk9aQt4XGKLPExiToUasbixf0ZQ7pN/q6
9J4eMyBsRm+g11UBDilmfPe2PpvXNiJ64DFpwKl/shtuHpDhuB1iqqGPCEKfCLlFGbc2TW9G/nMv
WQEq7+8qLhzg+5fsqQla6gbz5lu+bkAyUbBZ9Q8Fsd6NPU+IaWNcaSvWn9BqGBA1K3JX5+371TW/
iFq2e3mI0trS47yloD6e3n+04L5TlGI+gUeozmL39V5ZlfCumYRbiPmcleBAjwhgc4r2fl8mXoai
rcr+Td0g6en1z4NvMoG+Rb3pqslZAg0oV2IWbQhIR74iot7ftCG7ig0GKNsMbvugtxe2f5ELeyPn
l11OtlT+Nk0v6t2OeYWYZVZP73gnF0/sJpZVPjXSLibAMOxVuAWLZh/KS6v5e+quEesyPZ33SeCe
yX4gdD3roY17kGe4+a0zF3atz5aXGI0jIQfK1KzzI2N3s2ne8r7tkA4khj7pKbqfTYtoPGPRELWa
aof9cxIBh3M8R7kPug13wpiO8uWJcNFvdjV42q3z9kvrfL4QfmhcT6Lp8Ox2NOoil6tykrw6zjxX
OmF8wkGReSmUS/ZVyMmcsmfwMQBamXp9Tn2N4NS/vfb3Y9uIxqc/VdC9Pmv0P0tu8+0fl8/eO7nl
SJSeg76FRZdZPfCO1PQOKTd18TL3cXk92U71kKa85Ydfs8ufmAVOQ+fGFF3Tf/13yyjCau2hr0oQ
sNwZhpC24Ce9PhBK5uoCQxdVgGncTtYz2GytOUq4THNJdYZi4rcG/LTGQhzp25S4g0S1l8N/Is+3
j0S7kGS7gaaeze3RkE2drTb5cn1qSPYuDFelX7v3bbERLiUx3uaVCXgqm3Ws56XvbTuTBptJDNwm
IkKHtMr7/RJJv7qM7tHu7twSnDTbYu9Jj7Qg4TPL997iuFXjQpxUHHnOukmj2UDuHnA2ZjAqR5Ur
5Qwmh9Dt9AYdDHsZ6vQPd/mG0IiN33qQ+DOG2Urtguul/uvlCETrIVhV23ZEDl89VQiVLKcA0s4E
RhO7hN0j3oSX3iqYOA+fwFeNS/aRa0cNuG5db6wKKcRtQOWsoK2MC+y88Xg7PF/GseZ0KgsxNJvG
wsl9E4tSks3KRI1nIp0TpRdnfgKcfdUPp31CNjgJ6quj3pAA3eQcs6O+vlCmlsT+nAhPDKOgJKYt
dvQBWlleiPQbVethgzrIsomK03okxzSRaE98iLiOiPWgWWuULOCLRL+kjJFI/xgCOjj8otWhaBiU
k7PUBwlGZeWCdufkFjfe+t9W9pQmQxH8dagaRFyZ9C64ISeY/oakOVdgkTgWEaZlwC5QYEubnjCC
huBH9n+57WS3ZiWlzCwFTVW/noSYlYqVbtFD4WA2qqqRofdEerAlSb5gQEF60eEo4UC2DLSs8dnS
ne4tq0dKOOGuIMmmQB3+2USJd7ZrF+FVE2TOYaACbRXw1PuEMZf/YV10U6aH2ubXQW8CsDzyfisu
g3hV936up2U1SDgNank1JqUi2v/LRDvyW3KbbfK5RXsjou8qQNuN8j8RzXdpD+l43DxIMt53cswW
CtI/GYk5PfhxIowtO8EMskv7D9sIO4sNqaBsIWgJdEqv2sEMM7sWEHNFKkfs8nLOE3OjzjDVYnIL
7jAzc7LjxPMMCmt7CmtT6pgjA43RcTxLo+ZEgRbAJ2yrETXhHP4HKQTiFTECle7C3EBFhh0OCgfX
pAx4zAx2+jydyN+u48ePKulZGs5phl3BIv0zz9m7EZiytVALr3vcytBykv3wjm818jyF879DjgUS
BtT1e4wHRyq6I1MSWafIZ0afBUuS/tRooXXuAcwT9Zb8dYDCc1m/q69yF4zsjDW8PT++uS0AkFXq
fgTrY7lo0eycoGd6iQ46jOyqsA6Gbii/YFm+E9jLpBi0EGMa2+PYWSatlOFO3FYexd91OKowJIjU
xuKDjcGqRHgb8Yxfzt8sNirUVulbhMZc2FHyS7Ea+Evvb8kBrMrAVkBRtgXKYX1Bdqj+w67qOxE0
cPJfbY40QsDOcsy/kbJPWnku43Eu6tIaCmaJm4SeZ1R4e2t9Rng2GoaJic4BokI8Z5ZZQuypY01k
lyquX+IESoQpM8vaBLwOFIZZw9OKFhPA6uX8ni6aKnq60VOcuXrmy3FGYuMm1v1IA8Onwc8g2DhV
XMRvp9V5FeqaudfhJPu/NuEHowNwxySbMpW0+0HG75CWAtf66QLscsF5Q+cRr5I3c7/Op5+YuIfX
8W/Wtf9iAsV6u7FYeczZ1tkCfWtd1IB29ny58D84HNbe0ZhPvUzEfK4aZpbQmHEBYQrwRXFiUHY3
U0S0i42obXme0ZajJEGpQwCzk4PYc1OEzfRiLjRWhJwe0Mw2QoZE3wkVmJdN0lf1/XX4DYdTkMry
UDh28a7knTrfBQOmKe0ZWu2WTzF4PrkDhWrYD4JvAKWdbYzpjFfQ0k6x7AZt19Yxla07YH0e3umq
pAE4ccBtn3C5IIKes7m9RCbB5NSZkMN2qxo1cQ8Fsiz5s+GVdv81u50TNCwvi9tjjRE7emRkT+yJ
MKeLPl0O1yEaqI0WJ7BlEquEsL0g9pxKi/wQeCKNDK0K0wQTh/oABr2ZDG3nK+k0Kc6KWaqxDYjV
NQ6SJi0uNPFTmlV5jUfF6gaI6jejrt0/l5F8r6Mw4ryVwIPpzDGrc0RKp0hP7Qg85rl6t20Lpf8q
HaiN8HSwQNjE10LHqWh0geecb4IaMjrBNyfMfA4UnqcxJvuAJRchrBCjeT6TU99u7r1tVCDVg2DU
Jwi+SkqH1Arx3jNUgVsAeDOvBdP9Ebyi3a1Kld4zQUY+If0OzhyCrTZSBX2FVEkfsfJaHZg9rKaU
u2kwJMa8ZYBw3EDEN+2QUxWG9QHVbi+2y4XK3+ucnpxTNyDsfxHH9dZLhseYIcYX0inZhhXAoebh
ahnLh/ct16WU+0SCKT4uuOBgDEIfdsrYW/OaeWCgwWeTeSNvMIxwIAlEogdD7kUrdc8YWletpTKw
/d2Y+wOt607s7bqI4/YepKO3opyTpiLR60Pk0x5DZlqU8Xl/5xbRWXpU+IOC10Y8hlI18w9Vklf4
ILWzWkDS96NeH9eSjG+nSODLDuAHJoLg0ujQskwbSjvnE/KuOy1dQZVEal0nMBI4pIWdn25DXQ8a
jPQ+N6neWZRwn7F+JGXCJWc5zV+ixZn8XYSntxQvjwBdWepI+Qmpwvd0uTfMwIyr10ovVyH3tguv
y8i8C0PwgVakM5KR4PDHekGzUF4letl7Vvydn0IJ8yn4xQtqM22gndhMhBipwyC7ZMP6cBeyqaQ9
4m+iYBaqiE/6oUirdwTvPOTLVXTkx9Tlr6pN4+qYn0qGAumJEtaGpnwZphj/dstCqpx+hdFwq9VN
IxAPgFPKKBWJ2bjizufLwufH6mTR7uN0ffIiM+F8X1/zHP1Kv3MGTKwsh0SGzPy0jVky4Q1H+8Jt
nXUdO4pxXZOJVHRcRel1ACxM0JZdnOHZe7SkCIvkDKpRQZPK551FZDHSKpvaZWpR/mlq0rNpghzf
G3X/1UY7Qsw31ElavaN3Tf83Jb1HmxfC5CPNOsRLVq9bha2LUADltNfRiAeta0LXRdNX8e6UNYOr
QAa8vJdWGQjvuCW62/D7vsVOp4esOcEVZ+gjQ2ACeGrsx9MA8bp/738YGBpiMyPVWaKrO3X51tEd
6TnDJGSy0RDqEStmi6ohWGz+VIt+Zw05aKNdqiYVT4gm2WMKB76uOkFZNMwqw5vwfpuN0ftDJGpA
1YLcTsd0u8wCLZ4xNQpK+JbX16RFioEeopbqEk4y3Q05pbBPiKHKX9XxaFUjHAub+ucwDPRWA3Ax
FR8jSNWzPAL5iOpIzP2FOvtETTjXARVVz2y44SIDEtOiwBlcnTTGH6Qxu7RXmOnQ74aC2finkAOk
i0aOyuanU1w8jRRGgRQ692V2L4Bf3WAedIIaZibrsIMnXGn42eJmfjXevwnCwvhAMe8QfZV1Dmai
5W3wV/m2NNUjN6MfGqkrvQE1Ez4fOh1s9DMUWRKSp8negEwCGHqbMJ83/pFRPALwoWTnzmGOsXQT
MlDGtBTJVd8l4UCQYVPgxii40CP6cqX/yBVTVVvugigualq2ZROUw8VZkGfbu4b/G2wowr0GegcP
mW0rvKxxcw3eRK2gkBeMYHs292kbXhGnk4Vr1uXSR02Cbqa/ANOulmsHhGiS/QvT+YpT6nkddypx
QwqUxCwyYU70ZXpXVFkIRrHgJF6bMs86u1h/Rw6NZCRGFZ9yXyRpyKRrwZqMmx9AN0TKbvRiUnV+
SVndMXvMavg+i0rlkXYdJ/DBMaKG6eo3Ep5UwMz/QR2m9Q0PbRNnMrs0W0uQrmDI3F29RR3ycPBF
OoJZTyMZzxoiPxWhYYJnYRh+zeIulBphqXIjt18ayBrA+aW3wb9JEZeYPk6tw43BQQ8te5VTWc9C
nEl/8SVM6fHf5qI34TEfsF38Zs9qwvAwnPC9zFS8Bn91XR0VAcyGtVsNYC4TYns6gjdwLDaFBeds
5x6tcIzy3T82RoEmCYbBHCoO6uWdKUE2oSONMXw9TjTGOXHHphUxuoj41Fd8NUGE916J4h8FP0AB
PiGdX71uHF898StAxx1c+7beQtSjVOk8IkW5kM5BpXlkzPajSjEq5Haspb9MT4wmpaGXfnYZqcy3
cqFZ39AQEhEY996fOfzlg7FgG7Tbaa8QFjO41pEF1re0qtiCfy1BlJ82x0S1+6JOUy2ghWED/ril
8rrX2nR4iV3fSTTRHE5THPouru2Wt9JZ9BEcVxDHgL4Uweq8fHW1uEp2BgwVra94KyAMwtoYBBOE
/hb/4kPPvQ/0akG1JqG1uPmt8N+CPB5JfqMfxNnNde0UzJ9LAEN7EwgUKMbRNFoMWiP0ob8rMHOd
OVZv/bZMYER8BPn/SBioxW0DECW8P6EtPx2QQix9oAlxe/uKqgN2lPB8mW7r6Vr5sjEUwdtAWK2t
g8HIWzn+QXBLRIIyFSLRwPfvi0Q3yXeRtvBvy6js1a/XGkDEXQTLLiIpwb3+KhlMiwXeu64B77QW
qHk1rIPpRcVnH80a3TTgt81WIlq+sqxYXtlKoMWNXx66QtxM/DkhzXzvusvMPC/CJCWEl9jKx+my
1bYdJFdS2hBryuK3UMC6n0ZjlIgi5z2GMs4i8MJOVCtlMMlVqhOLtxAuZdrBQgzlYDyA8CLBUP5H
icKuB2E9hWAD2UnjYdMWfNAiaXM4wFtZpX4lnQZqNFRl14GkEqw7PZ8CloAL8yQVyuzCV9vey8d2
auri+kmk02Gn5ohORFR4yiKu8VtA3leeDlszHcnARIic5zjdo00Z5ucQQY3t/Ek6aruoyn1EVeHZ
PDUtEfnCv21pkf67s6nxmenHD8W5OGfCk3VHE3RmuXtlYicm5w8t/o3snifaI16VaWvFVKu/gMLe
iQgTQsEaNcam/83FnxO04meYAhU1mQejVHCfPC+oGN2xzI4ZfdPH4YrEl9FdEmhoWKirujCnflD1
p54gCPrA26XVkzs81LPpHhx9Wlzune6biDwhW8qOOc5C4aixlA6ngv0d1HOGjP7v/Bkg34j/t2wF
A2o7c90eqab6LPPcTVEsCdgz29Qawp5+PHa5rMTTUuk2+TTRc0yivY0LKAsShjr4kaoO9K9NGb+D
B/ce6HkR1ZcYehrunkjPt15OZiXtKpQvXCHNlhsngJuOyywJfXwda+OVqzuC/aJVr4vHJaoFkQ0R
NnE6o0LfIDAdr1hv1pJZ3xi5EHcnASfxRGQcZkH8BO8W7d/lnOVc6UCfsmxcUut3R6F/ru/JI1Qi
UMnKuhkMj4o3XqTNtY9Pk5WUhbHii80kFdWodWpX73YGCEzPG8JbzDbp3+l2t0iGdtVWZVYfSzUM
RA4AAJ+kKCEIqVVt+WqxurfqfNqH1Cozno/YrKVoSHVoS06xDuubdKv5iBWR60WtzxjtQVAF200V
XhdG+pphN7EhV7PynWFJ2VetbMC1ZdJQte/OaDYhIzbPmY7lvu4y9/yLciFBTAIQhqnv0fQW/m09
ZQ1tbiRM7kMaV2O6LEkSz0Zv5PnlDrOaVsNU765jaHwtm2CpuVd7PraIy44XJtd02ywV1PcjtkCm
x2FOUw29ZgrwG1Wutd0/WUVN751ncrV6E0VmzFR41+7UIL0w9APeDrKayHcW81vFF1S7ekVkUoGz
3UhfFgNzYs9B9Qwx2YeNpmsjdDhpQHEeKz79Xxa34yl0JrLkHumDUmvMK/1IbcaCrRoMu00nQhkb
HiyWVeToPfZD2iJ8Jj7g6hekUr2nvHvdLKqIKMRee9gduUzaX8lV3StuFDM3Z8fGQQjA+aPY+Kc+
VhttUI9VOb8E9JP0CBswTwBQaJpUWLSFVjMjajZ0/BKrU71OgbCzSV+Hgp58rjE3Vv6hw9HLOnXF
aedNpdUQ6bqbOtEynfIhiwtWd6EOWpw88NOwJM3qXTDAWPHiwz1J3GK+AxcJ0gcLwYJeA9A8QsK0
wD260N4c6Kg/FwSMF0l10fuRAKj5nIjkzbHfuT2JyFrYJfPT0ibzp6egc/zg5nFJUNDTFIbPhkhu
qVXUFBy8WpmIdtcoCymIlDIpvDQ3YQt8ErUUq6pl0AVfkyPNQ1ed32xEXFYChcZ9+++hvKvSVJlX
fBXz2epYRiX6/NaCAyf74I22Qu38pXw/iSGnXVM0aP6JetYv257Gsb1nVx+ROtMUFEbSGhToLFrh
XrOtnEZVd8/Ht9Ys4OZ8MiMjHEAmx+0rt3iDxd8bpzn1gbmisMZGZ25wxTdRIiphppLX/Nwv9j61
8TqnsX46e3JBq9Y3437kIGcYk7sIbsPdi+XqqKeYc2O/OuqZTtTPZFjPHXR5mbFJGSE+kbYNS+Pz
DTPu8yu9bqLCeuXNQYxfJ/8jXx5JUQtWa68LbKqFj8b6TP4J0BY0L4z+IeDOIjpv1mKw1qewtWqb
/+aWhGqL6EuOlqinum5VjiSKCWbREsp6U1aAVZk60L/0AZn6Di8vzGmOkaWb+N0A5VNipdhlFj63
8NhS6Vu5HcyJQXGzv3l1JeQ0jdcFnKxicxMAqbEFJPpr3Mb50BEHOacNePlpOrnR+xu4+rszF4xN
8T7CoTgaBImYP2j32vQ/IxUYWym8mgmAZMh95ZLiM7DuUogZcUoR16JFdbIjy4wkgfi8UhqHOQN2
mttpK3/Re8FyqkoxVNrTwH6ItJ+RO+8jE0NO9lUIL5MIM+kEhjDQGUL3qSTgAdTgSnrYRHbvdvYG
I9Im+1CeCdtdZozi66Upadctjne9y/MgWuifRNDYgdVeWvz5L9k9wGLgu0bVVwMP+8NVnKAjn1zO
mhaxCVamywzcmD1aXKikf6/vkx8PO860UcLD3ozeB/zq5ye76AuYsF5uHFXkBlmFTdsGA/LWRD4H
VC1RSLnuuS7+PePRdKt2ew2qeHbfvPWaxD4t1l6GXtzd1UYKyJEAOWcaL9jxSlp9XRhNKidIzD3/
YG1C6IERQyjoFjh2AyTrtDhmEYSibj5dwIXvZZnghEM7tuDjMQR9Ge6/7LP4r65KTGPnHNvIFIzZ
YtOE7bRw3h0bU2uVS6hqQq2NlhUy9N7KyEFfET4qw0lh5H9Myg/lmK+3XFKX6zwWbfCrtEt7aTdo
/c80PGRS+A+EXJXktYZNrOhddz5p2e20r0n8GHMOKigF0im47YyB3LnT5IRC8bn0S0kbNqJl2dpf
81FDWkQ9tj4aUSqu5tDEfNFGDCt++bIDhviPHm5+JYQfb4ZSZ8Zi2Mz7Ys6nGhC2erv3YTylUf8E
b/subTL18KDNGKpTqrhyz4PL3H4GoR3G8aaJ1Aq0MpxH6hz5gNctziYQEMIjYR7Re54tKCNrO9TC
mRK3Q5bGrC0e0sxsrtHa5ELFqjBvVaQzyMsbaWdCSHgVQfkKgUhpadFEs2GNoEG2QH0bflqrcGvG
rmRBwLSjFQlJN5l27w9n25wz+YbZ0epiT85hyN2Dye2hQaaPe9lCNVP0E47b9pd/w8Tm6mwpDNaY
TEro8uMJ6poaeZhJw9OGSdJHnC1s4NK0hFkDh742gPkeihsjxYaadmK195c/P7Z91lHBYXxGUlrW
A/cC3tzWfz5rcDSExZPfR5kpwGmYJGp9TwU71Zlt+ymXi8rWYlcASBlBIFMyiFedUI1aMOI5tvMR
5O/9xN2F+itLic1BppeYzqDGBa0gXkkZF5aWdFZwebh1N7ziJS24JIYSzFWtTRtE934IHb7O0yKc
/vx7ttiYNadFlPspGzf08ryXO4iCfirYstNbu/x5T1YJy7SqUXnyMsibVPScWBcxhlHTIGbrT0Z2
0AshentKmxi9+IhhUNTui6Zw1JSQLkg/pJbcKVyHrsK7DUfjpbX48SYFOYNCwFJp2GimBxGCBbOW
brNbwLh4+tAOd0u00j5ANnq9iPBttSOIurk02a41vlESuyyVsk5k2wwQL9QXQgLrhCEbgRAsSR/R
W/97nxPba20dl4fz6fNXuN7xLOtGqR8R9ZnUGKHsB1KmovqMBrwdHCf/aT0Y2dqvXHcXO1H6En1S
N78ql73EI0Jn8eSVumpY38LQIFhLL4Esj6cIXy7dZdj6DR2eDjYElCgXbL4nsQ1w2TxICZniS+fS
Ysdj37tbJ8TEx7ZVCcdoN/3cEf9cbp5wZDIkG4sq0yIrRVekDYA67+29QgqRHDgMS6cRJOOKrB1J
i98VXHe+HX/jLzy7G/6B27UcoLZ+CyUDYaekjSkFxan14s4nWVmOTXHMbBYs0cDYh37z5ECQ8WBB
Q5bchcGEFYpLSRzYus4ip54VBKitIg71AES0//qA32VWfkkmGYHaqRNqvNYAUgE6Fjf2ZzXSsMhr
JlDwvhg+G0WmCf7FMbzE8jdDT+Tw1iNMsjBPHaTl5F9KkwYoPkLj+pdh/7xEz/C1pBQ+3eCFbgd2
aTJYd7k+v48NCse4evinbxAylN0udkxZTCbB99kO67ah4SqgtsplKZ3VX3lPHZ4Mk8tOtcXKGqAg
iUpPXs3LkJKz0tc9AIJ3AW2pqoyQOE20yecHtXmVNwhG1yGN5fkMy4zsL0HrzTctD+tQ6VnaMuJe
YaphAK1I7YZvUEJCa0mHyqqh/n7M2tKYUI5teT3it5Tv6EGnTmVAMLC6NY156Epcns/T5z/ph+oR
ZfjPX3zAMapCqundNS2RoO4bbIsl/d4/umJUearyMZt7cZUjP9DICqw4TxI+38bgF9XDepkGwFIO
QbsRTrVIJ3TKlkw3PB1kRWNu/qk+t/bcmlpIcwIm6+URKC/zauWf+Gu+pKbqrF8SM1EQBhEY2ZuI
QwEYFsxq6pV2rkvQaNUT3nXpfsbqOKsJcLQ5FGTog12Y2egH3dM43p6e3R8ISgv790Yc3NJOjFEF
7Lk9sqvUUexa1S1sWbJUKwLolJEUdlFpfp9OSLmVoLUx5AyU9OViBkMiL2khr1QnVr3qP0tcjXV4
IA/jObjBvffSJhbivlpCC49Fw3UKLJzpLORgrGfe2nfH8IvTcUDGyY96P4VeAD0oXoEg4onpen5U
orcBcO1rdGObtsgP9g+hOZ+v2TDXrwYF7WqqiILrT6VCdImOSTAbHyNNKwYQ8duGGC0Xw1JegO/G
n1m1htRZuU91MqbmyCOw23cfWX+Vf1oX4hyw2ruOSn0Voi4RFs4ako2bga/NuQTktGfLFukCL5Be
KQbL/DX5zyUX1JYNb7XSI8Q5PBK0MPHokD2mF67YC18IGEaPLe5SLlk/eJm9rNwTVW7EdnR2EoeU
cQ0qwqdvEhMsxoF5qWxsqfkW7NclgB4qrkoG3P5bLHVW4d+6PZHAthI8NMod1Vn+M7nhdZxULjyW
2kYuW02XGA4Hm3zmYN+kOodp77HyA6NJtRb3bvirE55u8fKcNbnWLNUiQdjOSwfyxKCBjRyGVR6L
1KjQEX+oap4YP+wenIJS7Zm7uW5KSSQWKjVfAEca7jYPNTRqzt9KwYDd8le8I3kkC8LBPG84f/Xc
m7v3PuvQJNh96t8ZZ+iCoiPDdrD+3C8ShljfVfdQ3dGoj1y7EmzzWqf7TYWchX1qdF21sNWHtDda
qdgr4L3W1FrMCW87LaYQeL3C6tk8Yff0fIcavdZwCpDyYqpYPXo0kjedgGURfBZ/rMAjUy0CchyE
ie5tvQ4OPNtNhUQFlrtVjGFkkRxvgRvNbH7MctwBt/KgY2KnMHrsnyzwSAmaczj6pKxuTYBQ9ccS
FmE+AhwwH165xOGBcrdjaWXAPp68sxwiHKJc4MIdOOfuYeTsYAFQuVWkcilwlBmf3SD9zpZlO1dF
VWfvfFfJ4HN7W0nQLFr1Yjzl4+9A2tHWdXUrTfhcqA8NRYd9gATGufnuRrv28NksdwKClqCSX2zk
uZvgmlLRVDs1XT1oKZV1PLCfj9huNKUuOV7/Q6ITyyeTe2/tZJH/Ty2O9+QX038XlZSkRMZe+mN2
JhwCvays/5nQfJLHKXxFDu3I+V5L+zCXxptwP8Z5xDjDjF8upEufpCb4Fe1cCyAOUgN3i9pIjCFu
MZhFK8OUFJHGIt0IJ7BVak8ISOzA5a8I64fRvXUcCUsET7lYsmxrdloCWgLdwMaXAJxqmQoJCj+X
RMOfFuQ4cEtzrEjTHgq2tTml0fyfduX57I5LAtCfuobpVmc59NEJ9sF2fFLFjrce+hdmgqO1nRJa
SwHETBu2jSmI0ztyZKvNJVPlUmclpAdoojXFNarvozUTg00T2kiX0jaFExg7gYBNChsohgHpo0kz
q0GP0q8y545yUXDuDX/43AZfy+WTIjpLRrqXvgZmgc8kybZfC9Ry2HqX9AqXnMy8Jxsg0Av+fZlq
4UB5GfkWb3Lk13N71Sbx41XRJTFmd3tSHyDsmJwSaf1p6Y2mHfHsCQmQ/Cbz8cdwznN2L9Ms6UhW
WiHoSZhGYL3X0tN4452JmVIQrA7jeBc8IcNwPBNX4d58FTHhYn5J1pCGenny2Y43vRi312Ny2B9R
ogbniZGybtCfaXTATIZxbPdsH/9mvkswwtzYMpv1vf4zy5TAvITCk0oUJjuWAIFGrM9Au0nmRIIE
JeGRZHEwMtCoqYRoJq0Da2eDjsN9C5lfEgUk38f43lNUddHeGoUhIkXl33nbxacE424wAvLV0dxl
evU/atbFkSOywF6jqb69p6zg2CVK6TjKIXHapDDgzabESzMvEPWtORTw0WRIASc9shbfah97k8Cr
RTdn6dZA4Qkuh9Lrauc2DClDIIx0zdGkPm6m9SAGVLehu+WKKxHLkopIAnNDx+yGqKAB84r5pnJK
s6FbLOH/hYU219Mx5gIpA+4vA3Mkz7ZEp0RHACdtMfHulEXVFXaW86V+mlNeeo6UEK9aqYsS/YjC
J/D9c1zrXv5ulWm6DCX/0wMaOR71I4BIb55tuH3rKrmJQecMNNB6uRBoB2t6xXsQj7a4sb0+EkOs
VDk1oaDHmRYFihukQlP712CZ51f0mAzU5cwIdjKNiamPGYpYqzIXCmnAhHjO9RqgDkHdJKW1k0nl
/WEkne++CTAa2MR+GQs59YX6FXnDfcwtEmevCR0y8fkxmWXqaKSy8X/wQiTH2QwZwf4FFia3wukv
g6Qn4iKkNl3GjXy0i52kFNcjHm6QgiwJbNkeIiTYjNhf4GLfFACbH+x9bpFacg9MppYWhKHEHBYQ
D+Rx+i6LnXMEfH96KGwBuOwqQquRxxawWsOx0nkyU46OFJc14GRbaAJyC0TPHanYvAdZ5+VmD73K
LZMrYwsX103aik3cqNoLd0mF6pInKskqlkQVKoZH/S5J81Ji2lYASSgECu+hSs5A8Djg5QBo1Sg9
/HVJYwabUcpS/fRSZeFnsmop/n1KKa9Sm4AbqyjUlf3GyaxMZCFOD4yoNm4YD+pHoFPOzuXYhrin
weZzbnsTrxUCn9r/PTLaC2QX1FvprY1MWlNpuK84dA9rG826o6+C2Pg61k5f4VXMqPcAcr4G5lho
i8lZc5n61874DPF6eVkzn7BSMfhniPh6WqrPUd4HYMbnX6XHnu8QO5gjdfy/QPfArluxVbVXe8lu
p0GFCpBRMkK6vp7MRwZVy46uzF5F3mzYOBZ4w5xfN1Z6E5HZn4Qzt+QAZQ8tVvwLSWGcBl53XMUF
E9EHPH5HTQt8PjLl3JwBm6slc7zHqm8zYJTAPKPR8qPM+lEniYM2UQ2yoyIEbanR+3h9prOAO3vs
WLMgFCVUcUjyPifnC0ssSSuPDtUBtcPnAvo17x2olbvphHkGpn4nu3aWPKNNoChuFIXC13UO5UBz
/74tBWyLFIQhlNmCKl12PQak1NpuslJywQ8JoZkeCPVzhmfIHkv/mb7SciYCKb4cz1atIhyNQ2l7
+1Djrby9Y57wDlX7ZWDqXdv84CZO+Aw3NgK6HEli0o+ptb+z6ungqte8kxUZjkEyGAXMhDhQN9w6
o0uNfUd24PubFxSPkUuWuMvUjxDVejbP9udp5Am/sMtuTTAYjqlObU9zI+BrtNwkfX+8ClOYAQek
I6zQ5RDdr2cDF9BmAYTrugYVDCt6F+8+yXbB9LPWNR7xjeBq3XXh0FLTqyPFvfsvjr7Anba1A9PD
ZigtBpxVRE0czcF35z+QhjJT+zpIl0q2mwwTdQQH4BIztYUIDNvRiGGFCFX+Z5fWwp9o4RVE8Gqk
b+hHFx9kB5RMFhkx0yQ7ZCA2m3iyd0KY4Bq1Lf1ml5rWb1TQhN5aTA007otVx6qGa119Z48HQgjN
yowDcCDe15FL+ahcXhF0TSml8Db3CLdDWXXvzCXaiZj5QRfgJVf89CHmYcap9VPV1Y3qPM4zNwW1
bRv2lmllBXdjTVYYVwgCvwFzLBMRAnLzbxDOsUU8I7/8e91yEJydhrya195Uu5tVEXbGMLv9AqVj
K2046eGoB91LT5gMPsam7Wl/y4u59Z8psQhE16LFSfVZMeeaOJaYn6iJt/dKuAS1qtrC+6fAkJbe
iSUnpu5tAkQ3Sz5vPVWhaGXXTC0D6t8vmgVZZ8Dpzch/anre4IvrN5WpNT5ZwLHsEbedZJ0shIe7
P7rnZPUonuIY86g8rSvQi1L9nJEmuzrEy4foe3zJi+kvF7oJetVutps/Xk3pCFejv5dBWl19zYm4
vapgLb0+0dENDtn3T33qZC12WIBtT8MgXGP352yABZ2SNWSOjl1lJVw8jTt11XgkS2EzfGZ6XHy1
1zlwdyY1OF01jyD/s6VJ9pi/zNiI7PwuxAgGijOpNn2ZlP8hfD6hgytNceXOycBRylhluJ4bdrN/
B9BruZmB/bGtvrJRsI/uKyMel5Zi33keUNfMhRsEUNLnflYMUH2xymuT9V0wbxQCOf/B72PHfSzq
CrP1gXa8fxhxhe9K8f1T+v0O1kx4refkEWnf9qvXqucZ769f6feM4AZkdeGVQXmN7dHRIJQM0aOn
8n3I3pzVkv6KNG4fSb/N05UD6hWIKBDJPF9gswy7EX9C/1jpJNbT8xGwxL+fHev7u9QCi0QzBGOC
KbKcLpsJ7/UQ9casWeFTCJId3e6jEAh96vYpW0EWPE0oO1SzGnReXKG1w1HLnxQRIs/XLPX4Okm2
lQW20GzpW9WwHE9dQe7YpZUfj1uodQYkQnbHJo7d2MIRphP8x/MpsOBHe8qp5esx3pifFM4LVXbI
Dxq/NADd9qSbStFBgD8W+0g/6y8rhHrTIpVXcVhOQgPxbL95BvnvlVgt/HonZmYefFcWbAfFkHWr
OPHDvdpiUJRROhLyWZdjL2Q0XYbhykYuX8lLLg+pwqToQGrQbGIXj+lCxMz3PsODdO0xUCx9gVok
WC6LDrhWkfXspVxTuFTjjIocZE5MMx2glWXY6jRC4CBE2FPP4RW8JJiByoR17QQR/1Z3QvqgXf91
h3VFtCilXTKUrX1HjMdXKAbeiA0qlbmJPqYIzpkAWE789AuNZCqebQRxY8gqB7OHgOgXLxixNko9
02hgOr9ugHPi+EiSQ887ovmw/wvW/XHng/Ynm9S1VfoQugcMJpvP2s+/1/rAJAvxUFDERbDneN0n
CubWzkrmqxsjX93JQbDO+MNGeAk3bFRG5Lr+pbp4d+YDAee4EGoQvNOUhFjN4m4xAWsr2JQjJQoM
JSzAGaIyKTFN4ZkkpiRwtnswM3hd46yylXgYurA8zrZUKOgydIP43WwNUlhRN4o2HcFozo2UiX/Z
4kmlUSq6MSR5uwcOonfK9a3CTnPv+JEVvYf7iUhEluiPvMHq5L4UCNkKMkBAF2Knz5m0zv+Nt4mZ
u+Fept7ITzLKevvTOcoRrBW+fLsGNkjEL7xbLibEWEfnTlylqcEVcMhOtzOFoHk0Hui2qAhH3D4P
JYU9B6cOAjRORoJasc2N12jJeQXlUA02zl/hG9zE+YkPcUwzGX/n5nmLM3Nm4mSje+gNEo2jJgRu
D5oFrqOF9tFzqL/PNUd+ugE44/Dg5I+k5aEy9oLAUIu1Mq2vINCktKbp3qDj05nHbxpuXJbg0rqd
jQ16zZUOYdkm3mcvZINy5gAGFJlcYKOtVTP8qjHGAy8Bj3V9aq5bMdEpjMsu3kqm6SSi72tkeYrW
b/Y2HXWNs1hZvVubh4cuyz1ysdd2wAZJezNwQhmSMH5h7IMRmdpfjkzWGK3RO9Pa+PygFuCCvnBW
AFpO1GmVVKhwB3xgfxeQpz/dc+Xh9sT2l3k83hYPWGKDh/bwtb9FgVKRVMTqamx1yg12F6JOsgTg
dv17uNUvwS0/7keqYZzBBKU0yM2keN8J4QEO1kN+Nn1l6uH3PxpIWOz0S4nxbXlboJImBK3XJLl9
eaB/5HxfGMxe2R3ExjuQjKZTbjA8XUzjzvh7cWvlGU18hiVyYDFRAiCHvvXRaeBx8Jd7spvmamuF
UI4OWBAOF5rGsJD1hivHLTEtQQT5cGuq5NEkU81cHgxfDg29NCwTJbVlZACQFl2lqEXrFCWfv7B3
T7xahXmu62aobDvFV/y6T43fi4WjusjseFFMrNs8YqZCW2nc2zg4Z+upLPVB438umWB4yZJXiIsD
G+joAPb38M47AhN+6NHxd+S+GpvJzFj2sAJ85KiQglPz3380WWpSu1rwnllPgB6Wicv4WRTa3mxU
fCeHrckZo5Na969a9M6qqxpjHYpmemOiUtWIsmutneen9nnyJIYW4q2FnPKINa97AzZcmsqRrDgg
zdCr2UgunXIORMK1BpmKfVUp98GdoFJmw0IGq3eNYkMUCtZR/rpsurF/8Bec2aLP3D+k9stszArm
QwIuwUdAmeDbYlt1pfK6FRdjRM19E8N9GpRafNULom+gsktIgE8ecuinV0XykjRlCyb9qKOjqR8Z
qOhMKhZKfetjdsMn7aYNkkru0E3IDtx8Yy9n5swGWrkFL5WNxWSCiZrRL7f2gkq6TNot/1gcUnPE
RuGQiUUNRkJGVe3ZQyA8jbXC3LmdYVSmJ8iQxVINwpN5HkuxplBu09v4rmBT1fy0sJpGoojEtZyS
1MJ8EVKxamQTLmJXirFdjRDw49o/0AKKMfuPzzdbEqcLIM9OQF2PuHpwnVcXjgZR7hiZhu5YmEqt
8l5jG5AQKTLeJ1BaYrnDDCOr8xVZXLTxNhvlSuQk8LWNM+NmmK4+kd3Xpi25F3Ewy+TVfjPxWSWA
JM5BpKh+XaIXmocHfkOYgVRW6baLThtOpCQlwz9A+Yge+hjvxhlB/VfsHbCFnRrRt9jJStkTEWiP
iSqLUFdrtI5A4rPCt8bPiu6s6+QT7Z4J3/US5L4e9CoAWwoGgVwY6abhCoQnx+N9B5VmvBGS/Qoc
pw0C8RTtL5FEQNf70Xodm5qnx5lFJzbUcPUnHnYhYfJjHnT2Oy+gCtnTQg6vsnhGfHQtTT60mKUm
prtGxL8c8yHWOLMSXZeD8Vs6cqEgZ54nZyShgxb4j+OjUcjuHLseyYE4rcHbpdh30YeWOabiZB0K
9B7A/qTLZzg4M6HfGl5cPXQYJiVZF2VQ8EPUbeCS3yWUCD7Z9mJxXI3wXNn+wGb08B80LkqKSFQv
zcLlMRj5bYA+oRYRSCoydR1L6imT91wSJsVxIboMPIphpT2eaVpqAz/INLl+uAxyplHGZfiROn4L
f83fW3uOzjat8sX2d4KS69g7gymMcJmRYed/zi03BLSuKQVtcX4Kg6H6HV0IIXQNrT9D9UhvTbMI
ilzFDpKJEUqZlJa7NReFNV0mcruWJVl36uWEGc5ItG/fBWwGzBRrc8Y36axoZREwCl4DQ1Q9csr1
XvmD4W6zC/+Ow6SbdoYHDZcYoNaqS3gL9DTQ3aS7+TOkeWgmj8uzhLrhiNj20ehfqgGApljdiMJP
HyjQTbwMBwktsnvL4k/CiG5Qo9FaKUe1fqYh98Qe7LskObjkJ2p88H/eFwXgozYOfwFnxb222nip
JeuChuHRFwaTCLE8SJKOQb7NqkKPsWj7gsr7bmyTNeftBU+801wpHTi0NCJLp5YcY5FahyXws/rD
pQf9L/WFR2dOaWj1qEeYo1zAUG/li7oapu4+ZuQq0ZmAjxdNJpc0vyUUwecS3TxfaqjXU3dNry5W
jK//wAiwG+3IubuTccBWZb9X8Lv3Aiwvtb/XBxKijz9GmkIUy4VMWwH6zmc8DRlk82S1Hy/i++ZH
DWCNHupZiYI5HnqVv9hUj5VhaifmaY9aQJIqDCFWGsg2YpWI/6+2v9NztFuHMkWw2JM0Bm5NZ/dM
+6c5OgKDgJ2YFfvYJarOGFFZ3j26+dpVZqoRuxbhGz1Oe3kUHXMGffsIEbJmarcHKiDDg/s3ff5w
2Edpkm7Cj0TH0r+opP0nPoP9O8viXgUsIkaEfSfD2/3zL6vp4AeZhZ5A00HUFRpgYMlTSYIqPEig
GJaCLOBqJ9rVQG9eq0V2uRWa+IurEvQMe5t+Zdop0rIiLGZBmbpEjJZJtJHMhELOVC6AkOCNfLpI
+ZbIoouCtB69spOhM2RzesODXhjZdCRkt4SUPpQj9+3gJzWeHQyIkoPyCQRDh0bNKLealstmOPYE
BXXPww8DWRx4W6x0c+LtvfUpUD8xjTAoPecrn60t7kmKrELfnWyck+7Ynccu7F8tw1Sm1lLfI25s
Ftr/MS8ls0plGLQNn4MqWlS2S6guA5lQdR2qJvKRjtv7p1JUMA8VTgMdZw0x5W9rAseefb9FEUCX
IPsSLgGLUR0j/O5wegmEiwzh3aG8JEfPa08TLV3//1APnr2roYq9rmd7F1wz+oXNWMAyNqihB9Sk
g8N8Cf7hrp4clP1KF/Mq1DUh+iaBEY9bJvrV0GvjKK/j/TbaskOPZZb936+xJXdO+9RTxjV7vdEq
e8VLnbUwmGzqrj7KuF0b55gtyyWcTuMsDyoDKwLzASyxQF35UxVg2rev+tMNzViD/0AmgaMmtiD7
goAqVdGSO/ae+7eqYbvphv6qFHcQ9gjClFhvzXyCpJ1g3inMfBx7IPb6Oi6D5OaZXnHh5XwKv+CU
PWFbpR7pAek71eYN5YC8TvuASWktQq4BKq6+96lCsPyPYIsgjXL01XILJ7fWnvh3Q108tppxC9X5
WRXsrzdkGz9EUUO8B/2zQBVowNls4CYsZcigQmTxZxe82KbryXlor8EVCEuHBnoU38anhwznUM3C
zObmZr+I1sXYQHBAQoA1rJ98kKwlhwZBHhdA7lFm7XdT/amBef7O75pt7t8m/PAA8ihJ2zFOOrM+
CEJB/okHzIMjie0RKuEaTPyxeuy/c16oE46lGpIB2tZMvZKPkXJH9OF/dA+cnVfp5pxsNAk25Zrp
bNXFjlETY/MWoMg/zzNlhy2aMVYZPm7IK4B8BJgiG3clqUXfI/zUuDK4k2WqToTALyHoMbasvIbP
FErHW4fqeAUuWQ2iklrihfUgnDYlsxjcn6seFxV+/B6ciESih47wEqGhcpMVIVcYEKW7tJ8X/y8y
HUm3Rlm5ewcs0AhA4nXseVG++t0u9Z0fwOpnYBT/rrK6fU0RsbbOiIcH0dELdqCa/5divM5UlICZ
ptsz6hehWVuPn9VCx2ctH1EMY8Q82UrW/Irn8GaFZBvjHopdxUuLcKJA4DB4uzFSh7RjjqlV5+/7
ZPhQKI03PRFw7AD5vp2cg7YXV8ObhTYYL1y+Nu0wXKQsTfOgkH+qYzMzQpEfmjPjAhhK4BXCei4d
cm4+yuJjhw1BTpFfVRsbJOsA5wmzI9i6MkPmqAsgz58xUEIZ/6vWq1Cn3K2zWsBPQbIvduplKKM5
L3VsFN+yTDYYLCphK5hCyzVNNmY6manp/eoU4QVuYsDbx1J7rOVE/OgGpwBgqvUJda5H+XkG1mQH
1QC1w6lcgmlVUPvnLRC2XUTeAk9/zn3s5c48rA85PIvJgZ82IuzNRM6RusWv7PEXc8eEG/mQrw4x
Xj5rEWLZbdmsUir07Ava7nCdTI0q/p6hKtEjqsZFw3RC20oI2LwMKPijUvZEydcPbqKMAIoTMR89
sqXatntkjuqdXjR6JBoHCyZ3ckRpz80dVWy6tL7I/hpJ5g5K/Y4zfSUMmqb4YtmHbXkvMf17Xt91
2JTClpgiAHj2SoiquG+oDl+wBQjHeH9/yIFScm1nWUiYTYhQMfxW/PxDGzfkR3qXIikb5ax8+joy
P30oFfFlTQWMqXNek+ilyhdhaFeRCODR7Vmjkk3zQQ6N4Mq0SbBZDW0fT2lIVKFpUqMvEcT/ExB+
mbEhGunnNPmg9e3/56dwBo8v1DNa5fTR3Bs0eGQM8eYtrEs994nrtrlmxswEKev5NrHt3+3IWNp1
G29BAC2rm3+fkLKv8FKTR7acoG2oL4Oqy6wE7SFWNnEpP8eQ0jl7TE8zRgsEBARKL1JJ/t/XrcOD
Ms3pdtmiTUk4uwN8VdiLpjs/+axVydPy/Io09S13kkZHaewsQ6LYYn75HJam7Q6M9VyFNdT1Pn8h
jh+Spfl06ULagaqMirBh/gVG6BE5kJF31nEEJLzMM4w1ypOAXeleK2TsVEi2Q1vN8mJbbDk4CQJk
88y1LMIiWru6RBhTxK2VB9UQMoMCubS+ixliI5b/lQj8WZPo1ursiLzQ6CTHg1qHhCx6A1Unz91h
pTq3RduEb2Vk6VAd6IG1k3njTIzJQqGsPAktzFJxSzWYJ62xDQNMQnoK8p9s9GHIgXPzL72lfj58
HOqzMWSwI5WKqwrmZfDYNt/b6BfcChHfOjsv8CuAuAq2iAcig18lZ8KJj2hirRPfyUmDpYNvQSwk
omzTEm7zns7hSHaChRrPllbpY96mNdh6C1z0uW741JAQXcdglEpDjDbjweGaplcyL9dDwK9JgfVt
J6G3XJKBWxXOsYr4DGYCCXb12mL9RkJFF8JrqsK6rPgBChKCrb4BpfDKfBmFaIkiQJmF6EOR51kr
Wxew7dff7yi77VZv4MWtQ8oNZ3zDtE7z0hhWu/KgK/mYRsnsAHqz370U8kK2LO5xanSTd4CHyt2A
3z+u61em+h6PKndm/KJekKurvJKsorVO3uAMlKhnM/NPV3d2pguytoK5q9OAuOpKjXYVgsqXl0pI
iOlDjlnJf/5889n1Nxi+mAZdKUAb5UZ8ojBYkBlDM8pQtG9OeJumX7uqTKcA+xm8sCi/xJLaDUDW
vREMjUjEFpcTxgpiq9/6aZNPo+xg9fqKbLpXFXRnB6ihvewRLZXX+JvBb+dyMc7Xu8kL52uJHOSg
0ATKRDcx5Rc8FnzlehU6wz/sMh7TyPz8ldXPXAYIpxyTdm85Q+7ycRhXHWQFs6qv38CMGswO8ZZe
B93kVXjlhRzvluuSlGG9ZU4Xri+FeAq5LN7p3YNJYwMcSr4cFoFyZLSJN59dqV/I48jh2E9xZ1Dh
ZDiaQCbs9ka9357Jgoub2i2JWXj3onkWr1flwoGvb3yeP5PWipu8LP7hdVU/ku5whDTFuQnk+ddB
0OnbByDAjM6L3EeSOG5AC0xjfiUkzzNrUWSGst1DUU8SqylfDR34weOFV0xKaiGBCJhB2WeMFlr9
F51zFN8B6Rqx5483NgxT7x4kvZmL3AuXHfnRdlpHEEOM748IAlEv3Ugietav+0eU3QByfujEVYV4
aaupm8WQ+9ToB34gXceh3bks1RXAHwpPSDglweawgVaqfryN8LfDojpqKM4WXAALJnk+WxuEZCBH
7H9JZo1eyl5EYDFjwziINzDXtiNl3rTEKGYmUXLneEslAcQLhR7oD2MW0zxclINZOaYNDVWkSBiS
3V/Q+txoSx05ayyC3bAxB7VbDE7WQ5sWQGFOH7ogpcS+hWIWFj9M8Iis8fNfxxT8OFotw9iAvt5P
QkmVRu3dnE5y8ier+RJaK/yFIsxraWYt3ILJ7N7W65ZZjl3B4XBX9BeODBhsweJIlHxDgb5CwV9c
jHNgJVURhAwnyBzIbBsPv/JhwE+x6ei0iCf0P6CpFmnXhCeby7GIrZi/ArfLwJ1XoUwIUfxZPcfj
sVwuajjQkV9vnCqkmHMtb3vKCUf3MPhhJHF0Cb3KNKx3/Sbf791KgwvSssQjHDNyy+n+ecENT0+y
1RTuFxd4wgU/FuviOt19RUd4LJ4yUFFaPX8XIsG89nWo0DJ+bkWtWF16w9MtJDbfbuo7Cpzwz2bG
7JosskZO3LF2tlqQnS9smt/m9r9cM4rsHYmvEAUwkBAZ4PQkJyupbmtj6ErdQSkDM8jtxSLsNqyE
icowZ9UtLnp7pozvG5oopYHZMeIICn/Zv50OzVbZM4AFZ7usx7GxY0nbsaQqsBwlXRaHY3e5E3/W
T+uBHIClOmSpAc/nGZNLlwCb4bo2c8AWmXXnkXQcKshQqRZ7xaO1BEXOW6tPbXq5mbBTyc6fojBI
6GQCsGaOivKJ+aCx9cRcp9h+bN0YMDrVcFuYUmWFsobqGsvqC3NGgGmjOcwyOAmyntPRMPuUs1fR
DyGofiW2MN5QpM+Skhvbt5GsiWHuPwovomVz4UDGGvIyB/OKUu8R/4CNGDuDq1x/ogIkEuMpZ5gB
+TF9eQ/izKtg/rTyvPLTE+YW68FIreIbi/EIFqx6efEIVQCepEbTP+A4cA6LDFru4erlPrUUpz6C
1dlFiAKldfXl7rD7zr6ZWWxUs716KbtVTfB1RoBV/f9IJ1WYHrqS8uc+DdVHrsf/DfQ2hQvbcs/P
tsql/EaoxBY0JkiEU/BCtz6AnAtTOe1Ogq5oxEiOKuZQlnyboaNmLGJhnqJYIUvIi0lNAVlASHhP
ETR2hf8Fh6TXhnDVB0r41JjERIB3gfMUxspG8nkKaWA7TenS1SG1VWUmJ2pCIM8BXo+J3qYu5JlA
jGKhwfzGt5bBwaxwySfKFrgcCK5oU/OK1xczzuB31xJh3OCN1hW5Hm1KGltwy4/M7k4CYfxMTBRO
MHEnDcy1rdF1m9ZMgMETMyL1NHUVntMS5jOLNiegPKrN8gIHhhCrGfWBOtnnFy4xef2PCtaBN12q
oG4JZnHgFzUcp2gySejheTP7Bn+5GnRvHor6YrdrOaVEb1psaphzRkkOvSniSqii5AJAbsEgnLif
oHqw2mXv+0mZbrzm60ZOJMBQpVmWy7SRU91P4ayWlqUn9YxDT2nrxgJ32L3qPIe32806aa8NC6N4
dXHzTd8Y19kTBKe2zEgxLQID13aKSvwmhcgIzE5Zj4hTBDJ9mQh+BMlmm0mgC4GCUYJB03LgS9yB
1wUt4Zpn4L0K7+7+nEvuDHLv6oKqi9RFX9F+qr4Qd8rdY0W+SlrD962c0qPdGpwFUPR1bo1YnB/+
PEdxl1YOl/MLx40wQZEC8EXWTfeggaakQNrv83Mo1Uivx5C/AH9K3IE0iA6vGEa4gkOPytBdtSXQ
rO4x9oWVzL2NAr3a9cKd6ljUE3+EnYg8GGqeNOliYlgyvYh8/GCaZvukIGSBOiQ79DOZiGBw//7t
bznykzUZx5WAzSz27qCAjMoyZaffpSoxQBVL0+H0PuUm5cDG0Gjvtb6EHR8MSrM3+GbIgSR9Ltwx
eGxLn4etUno7zCaq5s+twsl7aQ8UaaEY0OG/SW9Jr7/n525rNO+BjowZOE12um3rVrs91tt7F1T2
4fOUIXSxsRR08rDh/gD9xv1SqMxePyhIX56rJ5HS77pXifvHy2wJz6D3MqSv7MzLx/jG11kFFNG3
9QGoAOTC5nHj/8d5FAJhNIomDcjMFCpoIZw7Myx4t/28ti9j94WmPDopsJixzjNIB9LMIzi3a8Hz
G9cNLQhoMV3T62GaqMTNr6PsdbTwMUEsElZhOMwLdEkWT5oyyhbWI4BcwEXieABtFNyRuk6OvlwQ
Ylz8Or+LMp31+zjYWbyRDzt8CQsG/lQFLCat3iPL+94Vk33++E5PAy32PHdSyw5ce7u+0zee3H9F
k9s1dDfkHCuVoYkJXiMtr+L7A6FO//ub2aSIlEVFtGIhUknVgnse8y/ick/NAtsNfZfqLpBTQh5/
4kRjEW+yiF41gwQhsS9SVTaMYQlLllWwFMdHME8FUMHFdHMPqLz1LR11Cw5wANRkUm3r24dsg0Sp
xlYa+m/tbdfAkbXq9qvGnT3g/ZZHZixLO5qAiyfRrM2+Ggjzf7MxVaQBtuPmBU5WIDeWaSoHKRW3
0AnK1dehb1m+b+P77fdL5xh7Z4Pp6KJp3CFNPVWKnh1+b0iHpvx+Ph8TNUuUS7lZW52QAIUpDX2M
mD8kRl4ofmILteymSefgTHfInV98NF9T/5iivqS/RNqpKW9AZkosh3UOGbE5V+kTlY8FDAxloz5U
F/aqtL66poRAAICyKhTaY2CfvPw9+eb9ESxaTSFCjvveIOK3Ua41QZA0kcoJw/E6CdUqpxpQx2qH
VE+3dBts2Xq+tooUkDEbzHHY2weTpOx/wrucdNRfckAnXpv+M4WbVsx6EUHfE5hPo/Y5F75ucYSd
RaLXbq34JGMzD6LRmX4fq5yr1g68X5dV774VWVvcOIuwK8pLEBiAJ3RMXgseNDX3kSoKHZ82qi/p
fq0XyJmHV4IKRPXeG3NKYSdgSc0MTfhLEypcis82Q5XDubSnmRRXHTJZ1x1mEMKZm3wMx9FoGR9y
9GvmcuDN0yR2g/LjJ34VlsGkvDVwgOYau5N9zQ113qqDfeLbQHSjh5HRSv3uWztfqMec26jmg7Pg
22nYGDD4VjGl97EJdzs/zB3YnzH3OL73R7GE1FQkl6MjGGsYezr90e2MAFuknewBC7IPYblDvSAt
nKtlxDCZFc3Q4sdl7RkpEDdR4C0UihfIK5iBHlFVJcLQD0ukU/FTb9UQ9YPtFJDvT6F9BGxo+yKt
eEfinxgDZFqI0gxKYPHCI/bMd0ICeEXY2Ov5mZ3mMEzCtq7VixM94DLLPTA3WRffgy8fs3plcKTy
qWFGK5KJ6HmTtcXP/xqjk0ptnWQyfzV1hvTa+tAclvn/hck+gzg+FjZZd7qtzMYGf1V+g/Axn8/J
ACFPvrMetky8cnTP+H3XraSwzskyOte/Vho7m0E2EsgziRO7ChibnszotYYmUpiccc+6sNjtKrnd
EhRXC1CVTa7deE3blTinbQRnu1nTth7yDBD7uDW9/lv/P72rPOLc4vsN63hSN97s8clwCOYfZJoP
T6ewMhdET0Z570yuTEyfzknrhVczpM8auXoiW/w7MZizshM1/3GC6IjrRlvAeorv4i2gYDllavuo
0OKRZter1ANYtq+USi+IUg3nA4amwQOEBhvoc4Rmzf3qAZNTlLDHconi5Mus9xPgb91kPS9dlRod
zSr5DhBU+ilPMOwKzXpgGlAQGsyKLQ7xb7sRPva1wGiJG/ye8A9wJHIFJAHtY+f4bjo1Z6nX4dC3
d/BN9SIdmQC5+OI9xQrbHXFTJIpztYUo6+0k1IDwigrdoghdXNzhse/Ntx8sdF3nQpUvcuBVFLvT
dGGrBJo0roFp9T3S33Ea4vnbSvbgrBSEMdnZDZn+tJ09woMGaraNTXscgZulgpVvjW2bFP71gvJO
jNl9izDnX44gS0zyYa4xUj6Vb3gw2apm5NhOQyAN9PQ6h8qvsUp022vhusC0FqRKJc6WhuZJYQDt
b5nEFxoSh06rqEutY4db4sf/UYEkz8D11zvVG7pDZbZmj7dBgTrJ5y08rOsHxnS7U4q/NEWo0/Ad
Z+1M4LO9lw5Oj5VJvb6mduukDjaB/+m/E9ANMBfksl00TrTouOd7CzE/9mPcm9NlstT1wEZM+uLe
i1PqSacFi/J9JgzsOtZLHCKREzTTApU8QGNkB7M2n5FDh/CoJrG1RvxlAy1xkL4H1Rk7zaFsKSwU
2WdSPXiyyLvOrS2lQlAbr3+ZbrraIjk+nd6e5GxAka6xX9oUbz/50k6IUcHrt1jY8XFGqjiXadFr
mXExl8xWzMpAGEOcK4AM+Y0WJSdP6l/How0u87n1K14T4sK28ATOqjMJX/P1TTFc+l3bpoMKglBX
8fZOZhGs/VAStQ+3eBCFI2kOuzwx+jsdC9yHmV4fnGBvueuUsiN9S9eJMxIabn7UceebFTTU+sa5
m3kVRM1mfbI71+2l+obor5SK2ZFroKjZfLdmrm7tgb7rCbM4XA66S3C/CWru0aS6/579OrsbdDcV
3C8c7a0UbDIY8u426B/zqknoNC1RtEcDGgbYy8uvXDAqe1r8XNIeZhfwO6b0PM8Jp7MfdLR7o1A8
yF5s4WNAH/HhQL0NjkQMWRISrsjq2mWbfmxzI6p9LAizpG5ww8B2vJ21smo5d5MgLKdWSjwgbMs5
jDI/66a77dO1Um97auVcSdireGxmrHXr0fvXvcPIpZ3ttFTcdkjW+UBDQb8RYgv6YEXsC2v5TAsZ
CpMw+BvlXGZvLxSYnJe/2nrrSsJH8FAUxd/I739rPDZdxLd19jffeKCCKNuMIRFgxUkhyeMPu5IL
roop2WuHzGed5yRpOftepdGynfI3apXCoZDs2gl8S9+zdKnU0E5J3hS9sOywIswoLEMBkdiXBt4D
PzTnoR0iSDl8/khnbLMT85WkAmspNyVYA63PdDgW2/gYs0vK+sAgJOso35GQDWu1xXYke0bgCi9v
9H7poIkC88z1juQONuVcVha4NS8gbYA/JTuWl22rZ6VQDfEK8v4vbnyuWYs9DMyPLgyflKnxELmy
CZcbiiwPGiUnxwbSrVZuPumDPwoqH17eu2YtjfRK/OYpaWsF7eqwJ9smiLhTGmMuEhz7CJfY99x+
cZE9teQdIUCuElY/FaDfkafW5fB4OaSz2A+yiA4x4qtxuBytW7MVxs0F63x3O7xKMVO5v4TWWxH8
0TzoiyXb4kUrKWksztAVghttHOFi/gViIFg4uPKmc13euFvbpd0WLDioOLr8gPSTzLumTUU9bAqU
t6iU7/C1a8s5yG4M2VKh3ew8Q45Pvt8RKndZvyN2U9dF4vsg1Vwm3GHuYk8vRfUFgsUoBO0Lh1SN
OMQnDLO9+RI2hPZflt24tbMvUB0MvZUpMB3/JlASNUkpMgrwZ2ZFFMbhdVwDjXppOdvOE7Penr6I
y80VFucEsy7L+3IbqhDXlnfFfjk5pifk2zBK0TytBUV/fYXS5d3JLONRA/qJuVa0C9FcCa/BZW3m
nnJQ5jPFrK1+Grx/whOY/HIor+VgsmuQq6Cx66j92EN9UVcqGSCUXDEGaIzHJGXnbY2CKzyAC2ZO
DBzHK9d6r4YHsm4tXHdI+xwG12voLmxf//Muc4lUuQYDJD2Z+RL+SW00Xxh+U8kIzqfxI8L+HBa8
f78MHe4/d99XNbCq7XoWwyX5UygdLUkevcmNQQef0J43iRpee50FcABcqv5+iQPPZ8v7c1Jb0rHT
IpWhkOrsf4GPFDvY7Xl87fv1g3+p7Y6UaLGlbDW8J/Ld3EkyX8ZOPhqQ4Pm+KF33UqUq55bve+DE
ndFPT06OXXZd2q8mx0RsoCo6CIeTs5hBu6SZioq9Carm8yD75tRIen+bealKOce9a8i4BeRAid+k
mA+IeVGSJAZyvH+rMJ3yuIEwBWy5IMxQUqmvg62o5AIpcLslzhcSx4Du8NZgA2Qh+7X9QTP6bm2+
CR8PlV2sJRPA0xR1h/d7m/3ba5bwOx1OToBRMRa7HZJoc/gO99Jz/RK7kIITxSbHS7HuUoahTcxs
icIoaeITBA79vKJxo2kEo/U4MKiboyr/fg+78SbQlkK7h/sJBOtupU76NtI62Sb2vlWyk7OmOYR+
oepSczQuLLxv6zuRrwGN/QAd99UTa/4OOMkyfwexb0OgJf0dhSDzGmXigIpUs4wppSbNGy/2new7
LBMw4p08vBNcqWwQRWkmyzDIrvsJh/YLDvPjXrTTNVXb31qc2MQV/9/sp79Z7avCWck2axas7uMP
OctCoTVIqy3KZqK5YUtjPXI9ePamw3UnkJRhSyz3KMtUIzrUBpJsuOTJ5jtLYxUTfAEAAzj64rON
+ESqeoXgu0qxxT+YwRRPFv0wq3mVWs0EVaOLnf/SXzWzFPVLhzSnha/IYEQwrKQWq7H+A6Ev8KaC
k7yiIrdd4ZVTQj2H6jU1cwca74DvubW/dkAw9cILoAk0zFRJccOml7vrUNLhTYUn6KwEh5Hh26WL
X6GwsjdYdbNo2NmBx/dMhWHnG1bsxtT2L79s4tM0HoXjvl56B0Our+1J5BbQ8nZhAFaAqxBf7gTN
djP5xZvvQopzUsdPleQJ/EBXXg/aWClRkbT3R+mlATuJhaTRFLhEOrilzpgRXuPVnYsUcKYzVbDd
81HFufOze/NjPVzpi0zcJksWwTG1dxk2RyYenpVRdCjgPKyB7MOWqiH4LLnuIGMWnbFLKwQh3Ijx
img/KTmE7NJu0+Sh+wNy79/HkMeiAFkrflRulIakFMIssxGr4qU1/88TC7GCkzQJ2B99aPdvUhHO
DTvZk7jMXojgSdclpBNLGa4wJdShi6ZoegEybpUnFnLi1bAARPz94V57eAoHB3QQzkaTzC02iSye
v8BDjgM7ssO/EtlNYywUAbjz5Dvy2V6j74V2bLXg9gjK6SPnTBYoFkD3UFYyZ3Ra6LvTq5fWip+q
mM1ppdPlfFCmRVsKSWWiOWCdUKco2KgLenA1WaKFgIDq4gxMczTqcIwus+X/BRNgAOpjGFMp05kJ
wrNxXGaxqp4MVbkgmxXdHZumO36GUUAxGMXq37hqEynMy8ZVnT7Zy5hxFaUSI02vycBLtxySWsB+
vXfthFHHDSTmCUgg+Wvs4BB85VM6i+ANcofAU+9c1+UfUD2w/R5k1A4TRw5wyRbZzbkK+zlJnRe2
qc5Qq1rvsmHs2U5wc65fxt5DEN4LueFILpkVECw2yMpcJKhWNLxPZtrYeUz4TLm69auUYNiPz/RT
kivGGocqANa/pUyNlSmJd6OREJupAtkHIXc8F2IDQWDkc4s+IClEdeUMZlOAYa97mJ8nALqYNn+R
T9gO80shNWaFTinIXoivUOeGVdnUqyFTLFhkf3smUkPzYp2sKpYEIBDpb3BcLyajbhBoMw3auMSV
T9mz1tYk8mAwhf4LZvnI6kNwggHBKX2oXb3WUTQw9K1pztaKUQknUfYZpWb2rcZ2VEZaGCo5JFY5
fgGPk859aEaM1O+MKeKh+/zttqUyAjYKYDo2xMSqnbjmlAsWcDT5Rjj4bIq1r592PTePG70khTby
ycj4Ph6L21GWBKTUEr9LLhsd/zgDdHyE0EIIV+6B5kcOLiRxYbDDU7EHxF2dP4VRkjq0IMW9GnUm
fPGBCtWpa0lVkw0H/7AN3eVsHssv8vpx3eHSD7odx2M5nAiVhkY4lR9y1ylXHHwLs2G109+hnOJ5
PeUFxJI4TfN9m1bU1ilPUZ+xDD1qYuN5sYkOYyl6xHUXGTXzFfq3qezZC652Dae9LCSXC/uLPVk0
QNt/A79J03bp26h2Mv/vOaH2pfvD4B90nNzneI9TawcwSPxp9y8TxRqx4lkrTPOLC3alQna4hQ2J
UT4vW5TCbTu/e66Q2bI0sILGhNMaXE58dcK9kreN7cIuGbj61d8n71qbsdk1q/pJI8cwYGtzVNpK
MEJl1/nG2DiGO0Af1Kmk+6dVKrN0zYiHAzX7DWv6oRlCqdTHcnHGiCXuWOiOOPdoLdjLYeScuk2q
M1DOpuDDtu0Avb0tFrVbclj7E6ZlZ5gORVOAXoQ3+KrBD1SN8ewWzCxiJApV8GxNkHHB4NyK80SU
ckie8CPNafJGfUohp8T3596P2mF/aO8vkfa1cjmAUgUx2SezddW6g+ZW3wBR/XWfm0W3pR1HTcTO
ybUVfMvRsfMvNqP2fGgr+0N0P1bGlbsz2NVHlPMWJd+xUNx01nmkTqUJaNv2LwuuqVjjDYwcTJom
2j4LVg7oZOxA+O4CdstOz2zGq4WCWCbBLUJCtiUExQlosEsRFCJvznSoq0AsRyTbsPttdg81/3Dd
IzQxf/NnE9cYWe7UK7qYJlpd5iyx3hpH0+iNAP006TXR+lkVCS5xSSFpTxYiUSLL068H7j+Hdhz6
a7sLZJvXz6azjIkIKOvq7z+nZsosSo2v3FoZnrSN8FSdKiugSqjljgsnRRosyJeffvSUdwcO9+t/
Yb1HmdJjyQHf2X4WDXJkRrQcMC+jfsFN6iag86fTVGW9toQABimd9RiV2edjnuXVBYs7Icwhya6o
Kdu6AjN9euC/BNcOzPdmHxN6hBnZyJwJRXqZA8g6DXa0z2KfXRZN870EopMd4xA20+eYa9tHXYHA
EYKxOnqL+IZ8bL6xpmg8k655NQEbIIaKWEaX98KhhszwFuu92lerjElfEZGLcTl1zE8Slkb+V0kF
MCaXDXDCYQMACADjsvObRcsKtk1yQRvuxO14BqgsXUJjrtfuNR+D6Bs0mZUKVKDtXFwTcIbNsFHI
ZMKMhZtEc9yV9Uj5TRkjhorgEqDhD4As8/lEDiP4ntvmtQ+4SPMuZXvAb0D8vHc5KpDtCquFmow3
O8MbzP2Q+pjoyOt+RX28+jabNNGY/rklABM+hTVzN6eejbGwCqqGLeRnn6yYxoKXAXmjE+Rximo6
+bkN5Wf28uuER8xslDFYseOwEY6Q0Qf35gnpJvbB9kA9KeozruafkfXjuOcu3+6NQlXcOOjVtKn8
4fPQ7GqA5kO+5PD8QMVqswdBT+/vTPlgW5ENJXb1YS+SmIqAoBL6qiSqtK3YaCPPWHx3YWdJyJOZ
i+cajvWTSlgAlWVMee9tc1PgddNGOVLri7WlBb2nNwnRtgGiDP5YF/leD4T+VkJZ9QleyYHqJDZr
nLhO+KZoOmqe3V+xslzGBOrCKp/0TSRrLGMiMlIkQfVyOFCDZMxQF3IViTRk7oEoZts8de4p/xXR
NWuHMghTSgRyBxC0WK0K9MgC2zVowwIl5pYtjLH6ws0DSgJlvEhPGbCQwUoLJe0WFflv9/fcVBxu
WSX0s15XXoYmXTpSPpzEQ+zIKXoJ9wtJdu9V+BwPW9LmyvY2OcMQ4DaQzUXUuVz83Ak9Yx5CFrvB
i44O5BlVYWa/peyn6++7Ca/NmxL/s6xm63wsAOa5wspGdrS69/HLoRB/HZg+EOmT/hW3G5MoMWKx
16C6q2Wa2tWo98PydJc5MuQjvJ4yOPODj+Qt/9mufhy+EFyXDmcPG/lvoMXgakLP7W3iQoCpShX3
VT5SPrOLjiBL1+v7sCaRIrXRN8/7eg8YkBn+/NvIWSV60C6BAbue+VpNwzUNjlvn42iUz6kypL4L
8W+H/yv9QIz0lweV0lWgIWn+Iujq0Qe+waBVRSAA2I39s+/F5FUxdIVwAjqEDu23ALq9OH8g8f1d
fKE0tgbu9BbhFK5QzT9FWzt9/VtVIi2py19IekrCAp6zQAto8Sa+rnlesjaifq1b/RoSKKmThksx
xEZdbW6rMGGHZOs/+AQX5BFPDO22RWCXfeXteEea5iWAoLGJ4ef2YIImDNHBm0gm4XVwppnDfbb1
kaD+N3QUHgaaxt/V1OJzvV3fnAbIcKFKIz3L6hX5NkLRs97bIXQiVxj9M8V8XtHiaEs5GS6sW3me
nbJU+nd7JBwWWkDViXHSo4mhAivcOyUvOiyd0SD5a0ZyByE1j2wcivV7JOkD7Fr7b+ADSURZOCoo
UqepQdHhEHt4Ke7MeRJeUYP5EWl6wjAcsvh0nSO4rLb/DVb2mvhBn7W6QapAijp5+/w9CUXu9pTf
3iJeT6qXLd3LilbwTshSzZhIQ1/53cAbVOwhjie6q4SzU9SX0UUY1mLVXpS6Jds8yXZLCW4asAyH
AxtsyRU4Gpmq3q7KSu97RCR+ill7IeTjWKJfclqOtXtqHias/vDG5AFe/APvC6sV6QzDNlm6pgJ3
AtuYPwSZPm2Lr4LwoHdkWNljFyAJDU+ZN97r5guoONEIEuUoSTHzjO32JdNzmGgb6DIQMc+tevk/
9e2hcARHrJc4jOl/6lQv2hrr2gSVWPkRPRGfUB0V51ymvSW1HD0WHZxVQas8SE5JFVS8Gv6o4rt2
IRrivqJIT2v51eD4SXHFbaepf65v+YOatnM8CcMLQ7rnDwHjLaqDSKRqSYVC/kvffIfUxbPi31wO
JBmpbg71u1XuIV4i+hnvT3fVnNxdcW3Ccj6KgFjeEGBgkosZnA3vdSVipOcIV4DjpoldymMMfAMI
gfIYC2YcsXYUKB/H2AtAdZxLo00MVyBe9eg8PAdf1KwAQy8Ra+XwDw7Lfuyw643/A94s8kfI179r
Mv+WLvpw+I05U4HGgZ0No7VDH7nYv/F0vRhpYkkOnvsZ3KR0w6XLLaLuY6VfZHwBXftWQw4g36rc
6LOvcv4jEgcAQGV1cfKFwMiTX0pSaNWAGXhGpG4a4pAy3qooIac2evItogwq4ZcleigF6g2Sk4to
UMai1fFBLq66KLcfvN8C9Znp4qc6F/zE3iOeRUcC954A5Jj419rokrR03oMSWe34FjBRxHaYM/nY
OKXBnQN26BJEqmZBimjN+gedEUkgL3z6TH2PmOB+BEjEyWAg42sb5T0wFYaBxlf1qfZrfCviFEd3
z55ifyJ82OBOPuQyRv+pyzWRpsZbUnAKD/TmzsF8hR1bjfYCRDqy9JOE5anwMT3Gt13f/vve2d9h
k0Dp/k3Jp0xcqgRX+XlCUjBLRpyYjt/LlEcpSH2AZTKdStJpHYRHpW9upLsrZADuFpC8SIY2tdGh
bwaK9I0BT5FSWjlqMcTgjD3dHqEBUWMLvQQchSotgKZCGxwdv+VSRZcukXyxHYPQ8Lb+xsuI9MVD
FU8st2jvK5ok/gEVQDxi52bx5GcaDnHmTp8n4krwR5Hv3sxT17co4IxAu9JXaHMWnNuwxzYbNaU4
DOOpn3EDzRwL4PDAKINe0JTOvH4cWppFgYu55pw5NJwFMnQd2SoEP5vEOwIaRtQSTSIsXTjD68no
hprFaNyZmw6HHD+d7aTkZkpt2XEHTUANZXAENa/32G+2buMzsMDVu5owtxIxaUasQ94Bfob5EScI
XiiZS7fWoDfsZgo72RvAXE33UHEM7fOFVsPThpQckKau13Y2CcTkIcqGXppNoDscMBatLGYr0UJE
SwLciM0hLvhRHwtqKkTHbB13UzxzD1Tqq1EYfIas5iqiYIUbd2u7QPil41waaSrpMOY2nMS8kbhU
nzafuP4EHmedkQdWYUIrIuV4a+onHFKuAZqoG2uqOasnsgQ1r499P96L2sWk5gzxzo9sWclcWzqJ
BOfXg+doRPetq8dhjm6g08UOBMwNo8cql7phr2htEEfBAIOc9vDQPxdiICWB7fAlB2EzeYsSmtFh
oHt3M9HwYggt5fqB/2a/2qWmY+9d8vDEMjKyVBXdNoTmyqRVY2dD6n8UW7CPJh5ekmF4GLI6DBKd
9F2jkR0DCX742N/R/L2dohPb0DfR22y+L1amPRsYTXGTC+QILJ8iaWtWGEkOXQ4pUCU/vf9vhJe/
SgCGm7DBqX08dON7p1TG6z/vg1JP4kUujuoSh6fAzNaa/iiF6dBBQUPwFPmaWI52Zdy2ZrVDsVr/
8tQarryW8hS+keojlBGLCc0WyPjZRbDmBtXnB7HX6DkG8STXdsD4gD3ED3tnZvoPAQpNYzlcYXuC
L3ojW9dW7smJvZuGVeNIFOEQ6cEhnbKjP8Rxpr5/UzNqQ1PCVWoMD4tc/xEG4OQG1bP7/xzDtTMn
Wz8qlhDrC90L6asmdVRqdWs8T3FWtQWdq0BjlSnPWWQA7Z7fwXwcrnEFP7gJ0qzaEdK6njxYN3Bh
cs2RFJx77qG5Wj10+sGawflbFxeU0hIGDkQI5dlWuui0fiz2NeXzSeJ4qEtZpwZxhyYWjLpIuh11
1ifb0plmncNvgGXiZxI2nBf6YdvGvOQFtHBQ6QicxgxAHnUOVTBV1QIhD1wjqPjqdopCgPSt6dlY
9mXs5nlQ+ffq9rsyxgY4+OVZ2lerJtnwO5m9kbdniAqtPhrr2QBiIfntmriPAuzQaaUPYz75qAB4
WZUPfuuUQrqi9r2PzzqoC9YcfJkMNa+LnCd5PYLAT7fVGYnVGFk6D+3My8RX0aklbLBAaxt64kwJ
Sv9OXfvNjWCXxtrVFRXCmw0OmF52pM/q9kmRvt58RWGXol4IIreq8BlSmlo+CQ==
`pragma protect end_protected
