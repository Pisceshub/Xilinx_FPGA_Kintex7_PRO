`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
BCC9rc/UvLO+60OKG37h+5K6XVw9+xBlmGSPNNtCyHiGBNAs7uE+P7kAaWn27GhAeEpR/kFMWCax
az/GVqBT8w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KqqDQUWeBjbeC5Do4n6RoTO+nx+zDp05oc3Bq7j9aHdTCyJc3x0fyRiN85/GGjrUv39QuhEX8Yfc
PQieFCLLhIDiLcaO3g03QeMtoC4gucQf/+wx8FMN+etUNIAKvGSpHcDF3sE+QU2wR0z9UkcquWwd
T7s+2xbq6nw9IgjIn20=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ArQFRYMFjfIqnM01+3BErkf89TR7vHqh8+aVuOpf4ehtdLgHJ/5eVLEiyKB8J8p19WP3coK1LCXX
zKhiKuxxeGtbGwfm+yWYlBx9ENRZgRCMJMCvUsDVN2so7XdAPwkjqSnh0W76/Lhaf+d+pvRWlgkW
9DQk2DdXzM4eoYWj8692SXfxs2GVr/LFsjE70VNgWii3g4b6hbt8arRzcBGb7WdSP01/Vrfupwes
wvc5UsRUnFw41z3BPXfnJG4S7TLMUaKkpXt4XkwlgjRwtf/TFvPay2nUHGQKbMhpn3k11OWjCVq/
je5H9c1eGYvQsLZXkrE0A7BXPj2zxOkaxG0eew==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D+ZRBE6u1yF80QejORI2YlK5RectTc5Hc3ZGgcNzOnHuwsKdRLXxgO2EwzuQORFrUAcI2O1GShfJ
cDaxaqcC2RUD7RA3O2LsbI/gqaNLWKfE2cPM5kyY4LL3UpWPM0Uo5ak/GypCYQ+UOf0Kv83mOrCw
gTGIytvAqr7oSLY9s9w5ayy04DJKSe0dAiinfq3BJ0yg/LnSWrLQBOBrA4Wdb3lM1weRawy6ucLs
RISAq5pL8KX5nYwI6yisEb3R/a68Gt9JyNzCGetfTfKa/ZmZFgr4Mj4aSY4hNGRM3OGia7fX8MI2
J9WLaNV+MP1mjqAewxP7QuQOtPQpJ7jXaieBRg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ntat/Y12i+xTz2OshnCjcnc8y9zrqQygo70X+7SJQZtc4rY0Zflni9gN8Z4mJ875xuUjX+lsIH9Q
3xBNfK+u4PKka3FGIKhp3P9okYAJ4aQHDoQHPys7ay3p9o+QjpDu+LoKsYOvKcQvSTT5h4JB/ADm
8cRL+CJAT0lnMoC1oD+FzJaGD6rbUe/m+ozDAZO3EXBxQhmIERbrgUps+YqPcCfIPBOirPKyo36x
gPacfOHCAyEnDGqsYlZ8/OKD+fUUWGYGW1h+tcsLksdUksFOzpwjaG/aylVqeGnpGGdju9YCZsxR
FTDPxHHSYbWz1IdEVen5mJ4AEFHyNM1FWcDu+w==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iooVi2sFmNJOwue8KHSUPRW3tf4tB3uu74gs8Z6LDvu2knYgcu9jq++JPYpGEqao7R4n5XlVPf2c
k4alUHvp6Q50up5xf2+TM6YAlKOh56q9Kx06TJnkavZHpzcVUxjTO8lhG7ZWXd4Gx6jTrcXay9Lh
hZnVvqIrYIf7F2M9BVU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TKJ0HbePLQGnDE6xQ2nS66ju3E7NpHUMIS0eN5TmIrTiavo1ur6LEw91l2unykROGHhJ6ADO8P3+
+vp5WK18tY3bqWh/q6bhiVRnEA2oMtztFhG2JpSy3iPMMzKWi7QDcZAMQdJjnf/G2+bGK0FCj+pn
IcyQWYXOLQCp2MP5UnYVxp/1/Rseo1YZ2mplACxSxS0C9v44JZ0uWfMD6EGmpBALrJusrcpykUXD
E/ZZoTwRUL3BWG4AsvhqsJUYITtSPAjRUg6DenJjWOgD37PK6P1nngWyf9Jjbs53XYO39akVpu/l
Uewa4cLxL6R5/kYVDFXX0OuYcl7BxOYxaBLIeQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`pragma protect data_block
eAOL/opCDzBH1z0QvPCIvO3t5YHaZnTDBeHrraC4no+qmTO+C2wkd+zvRhR4lO0xnYZvFdljfnl8
bc9dnZZx8LsI0m+KPrTnHbt8g7ipH5w+hK/P6DerYD9tsxaoruWijvVZqr/2gQxTIz3r0IoT7FbJ
qN3kDD7ueUqCi7Zphz5ablbkuUciBmG5Cf7FtDUsyquGpA3F9T5Bflr4kTPPA0oFoe9An8u0EQ8C
o/U2w6DzEXH12qOOwQJ2BSacgbimgXbdJUGelhAYvhl11iHvrdTDgAUPO7l4/ZX8Z3AetCREaGIi
Zk53hRXOK8Yo/Qtn52/7Rk85XmDYU7EkxL3zFgUTwxixMjMAFJPYEYV89ML87OZa2KVlxSrEz/lf
q9ik1Er2Zoi+YX+vQzHKICPY1DxzFuR3ubkesJeMVT9nm0MEHxhlGXbQD2PmgvOOZUoCzKzVLsII
55KMKomno5VuQk1kMAVJgTR1QYb4i+ZlPnUPR4xfdnfYOte/+YOXY6EkVwcPC6e4tdV0BHdChDUF
cooZX7bd1eI/wP2QuMF8ycBVAtzxOYGGWttRaxUyWL4Kbv6GWqBeu06AC2f4pzSiduzYDG0Fg9Cw
VcKtHfh5208XnBwpbhnW68vdmnNUR/lE2KjTtAlNs5VmMFlgyzTBnEMOKzSatmsmKW6d4DNEzEEu
HKZWDsrlBGucFpCvjVhDyPIIZy/O2eY7c6SPUWtvKHXUVjz9LrO8R2ap5EohTk0ry/TFnU9uQ7wL
TJJNU4ZR8lGsNqizNrxndwX0AUcC1yVfO/Y3nkJr/MiG33k+skXO0G6bhMjIEK8SVTF08fn4xJ3R
M5AvyA7u/TuJFOd3gTxCj0PoYj88bplOTbpMvTu6VrfTlGuJAd85Vy3ubKndKfPULNdTlF+S5TaP
drq6B+YKKglEzTcu7Tm+M4J3ZZiBU9yRZ9+tgOOCH8iYoh4g2voC3Ic0WkcuUe8f+2A/iaVClHca
39A2r2QjbgLupMlvCA/OTEAk3y8HB4DJu7dPlJ6zvbnuC9bQYXwxPcWzmSBW6O7ba++FcK7UzhP6
MZz3HCN4McYS+7qK0Ljvo5yNohRJrgj9qXhd0vOUt3gTAGeqX/WhIVUQjGTHoqgSU5U2sqK8sr0Z
8BYIvCod/nryHO0W65u+2plq3Gqwl15a9TdyoFK4i0zsrATWdZ51T/CtE/S0WmGneUPa/IywTlDq
+jI/VoasKXcJ3gP1AhNaSETwltiZqapyuD849blBDgtkBpweyr+KLNAzppm1BAObLUWFAteW6uBi
X2ANOjlua/SWW0vK7k13nYQ9Vso2VX5h2RoDw5SGgQompCrC+VanI2BCWAQZRfkuatGOt2kIoHj2
SV8E2FCR0w+tZnnjo06xiumTV+YYGt0u1XoWoAdKJqusMiJrddO45wh3MN/k3l24lf/mqSb81VlD
N0OEkr8El7o4fiGwZC0+lHJO4XD6BzQi1uzTNm5K1h6sYaaUj9D1zPtNZLVDvyVbUXWVq/vEMRZG
w11dAOIwl1BtD4MuEobZHlP55hmR68cLTYtFH3JnPOkodaNp8BsN8bmBaUde4xd4yJhYbb8cjNWt
SeOT8yLU/VqTHTMlT0vJKh22RjQKydR8qLMtCwPFb/d3jCMqkQAKXLGAt+YxIj/Lguyukez+sWmE
1o/mnNu/2M8EjKiXg+8WealItDWdw4lTwkmgWaMU4gSkMMmtjdk4BSXRlDA8Mhi0qnyFOK/7nL16
HCYkLhzBAsqRrCDS3E4P0l5RNNsl5F52G9yts2qA7jZuX/EEecCX/u7pP1jtR/Oj5KVIMpQTuEIX
mVHfR2Hd+hruEZiVg3vbqcRo2F7ARauouzYTyoa0Lo3g+0cz/QS7B3FQHrx4SZDjunNayWb/K9/p
g1Hh/s5+fGBoMQ0r8GXZdRKtykzCYYCNFtTb0R0zOai4IwC0OiKvriLX2O6FFssoVa3n1KupCKHY
900k79UVulQNI709n23K/ZDFtuJD6T+QkMScHTbKSS6+sHwGuXO9rYReUgDx8qDDS8YHeJxeYaMu
J56bWW3y6B2edzLVwlEGq91qTE18Z7eLaFPszAxLPEUXMDAFU+ED5c4fNOh3qw9RDiPGgQszawBN
8BimPhWpRs/BP/qGKaQ0mlWZI+mJcflStVkUzzGpV9CM0hyVgEzi/XY6o52OboJ6kT5CVcq7DLiz
3ABZ5m9eH3QFMcYkHxyzu1tvpSSBmlpGwFcUlBDPFfcs3fAYtj9oYRvnSs4/9HPjO+i5yld3X8uY
aPn6iA/iXsv9hyqQrgbckGhwKouU3EcmrjEJnXg38zLm75fza2GHhfDGqDmRzeT17xePY1GJ7iC3
qMDJUU8dncaa/6p0MVwY/jUd+7rJ+yLIe1oa+2Qkv+vtK00Qg9fLuvoNaVhB1TT4hHiNFmluQZOr
/ncJtmeMgZCnN5fe4GbKzLFylVXtvDNXNFmkLGpCFdh5oA8UVnmKVfZ2RILH87QPc21QVV6i89dX
ETVD2sMg5ruL/d2EeCGVqGFTh1ZzJcOROz3nQwqvR2sf+PIiI+6UTMcsMDTjtwQS1/9MrD8o6ZAl
FInwGsnlZeBAZkvM4liK0VAWvolbzLdlgrwiQIer+PbdrYr9YkZnQDvtI3wPq7x88lxYsT2z0YUi
7SAScYLIls/5fK0DbWNTsbDrL8zIZgP+1+i69Tod2ncv+S1lh9TVZS8qe3CVw1J0gu9qmgXfWyEK
ZVCF3xpJz6nYi28LLdl7EVyodswiX5rmsXRfPEHk/9tcBzMG70ExMreipVZPENFe1PTB6aGi9yfH
FEbN9qPyB56JC7O7qj2B9aSqLrpDgZ54UCO0QIK3KuRkpdJZyCkwZRseNxS6iDUYsBKW7/KUANc7
faChFpuVkQZdGpQrp/uEaphKHiETsq1lkS54mQCrh13GxFiRh5HoKtKDAYIz0k5/w+d8hzpXGR0L
WBwBeAZkFGiuCxV8yrEUbHMiHZfMsJ0cYNjyQVT75OFLbQHWtrcVVotHjmC1FfaZKY1V0PDhYDuz
L7p/6GTeS7fa7DedyZoEs8N8Mmqdnfa5i/41JX4Nbi97+maB8mEyzqEpOesD9VFQmmUngQRuu1aE
G1+qHMyG9AUDUk5DA1GEP1L4EDj3pWChu4z/iJ61q5AyAFG2XQ82sPlm4fmh/u3QmFX5+RjUkUJs
J8pL4HTl2ARGb9AOiTnqET2LWp1PYwZ0R4mx7wtl4cx98K3PtI7o6Sq11j5r1Ji2aB4yMskieJTE
45WhCAbLn6xWIGiZRix2X4pMQeyBf05PypPeiUMvrEtyV+orNB7L8k+LIBTIA4fJj2ArnnVhY+So
FEEjIBLu8DrtAr5g/lVeJj9lLTsyN2zKbvkZMU8hX+IiFl09OL+rDYB8ZZbZsRRHSpTFeOEODKu9
CrII1fpwRpM95H15kkdQmsV1igII5fQiosdZ4cUW+Xqa+HwanMcjhunMXjRH3nLY04dg9XJblTBD
yCCzHCsvgds/R9xtveB4A62r7490vN6/BvtcSDalCwHoYdEvsFXZIRV7/ng9PxH4lfXNL5J4gZ6o
hd3TKS10kshHdVNUozdgHD9L9/2xqLl5d9ONLD7ae8avHRGiat/hS78xuebUxP/GES1GZsiJ0hVQ
t9g7ggSmjqT58Tk7rW9bb5C9nyK7qFske2YDaCzyySjKN/sRDEjT3Fdl3N/kA/0zjVvQI7lBOjq9
sdOdz03Etcc1eX23aEo9oH4m0zhEIdWFJgvNXIrX3jKbPxbNAkj25Vdv2zoePqXfi7R57OBZbUQq
bI8uOjPYC/3VBRN5TF3PluZ3z3wcauOy00BkiCM0OCWtHkgo+ddvsezSP/ugzaJ5Hmiyo/FgTexl
XzT0B2ufw89C4c2RFDd2kHA22TC8aK2I+C6hlUvCslvynNC/BZr2nLYaoILsQ/Io6Apx0dPy7tnR
UX271DnaAWyww4eZFxSvMtZ4ah5nyTMCT08wir/7dKNxBumJCPAx/JPdcWVZyGx6RkFn4oUXnL+U
1gGbIOuat8NNLLux+vnJg57Vm0fhlW4Wq+6uBvvFvSCyrYV4//KAwvHO2QTUSgNfoMa2Vh58e3k0
huUaYRiebEHAoBrRW2ToLOy6MBxxeRzfALkNyPZ9yitF2kckdnaRaZM2zeTnz14QwpAScCFV5CM6
U8bLXSLRY5Abnp6KINToM2yL4Gtcks2kdhba/z/7n3uEx0iyVKbwbdOKweSKpQPD+VQOjEK5sVsT
JfpXSmqai7gsZ32lcvg/kBLKd6jhyW67/7CrUfxsakhm7i3zP+NbliUGuo+tCKtwqCq1Htcepktl
NU+tz3cRPPDVzK2Il4kQYYR1SdA8LHB7AA0TbdEbUVPGRDngqsZE/f+5VCHHSN5OzFbCHW2ne/nB
CX7z6GDsSOtFLw+kPm6hu0RjJ3AgyLkstUVaWXz8wt5u8wRA/TBDoXekjlSfwViv5X9baHk9f8oe
bmMLEkY9AffBYIU8UKbiWxHREBhfnIwZrn7f9+qz/ic65JhzCxabXFzJMnC0j2WPwKtKKOgpDMh0
j8qThrWrIFr/ed7r5Bc4vDGdeJtCyZM6nCTYol4BwF3bza7e+U6WLF9L0f0sA++ukQVTwbXTycRg
Dcs/ooCKQ59+KzVvOS9efER8ChGqYWFW+F8H2izaS9AFGoTHpVa2AyDt83W3BtfH9Uenj2Cv1aaD
u5Xu6ozPJC/OvB9+foyA18UvYEVSy/fX03RoEjnNp174/L8AYc04PDWcC/c64Zha0UAsJ/Iaak0L
8l6seNDJMwcXa2EdutZbFI4c+umXADZFV5QuJSPny2Tl3af9ZzdpEAxcw4gk887lzxTWhMkppqPU
Dn+9iUNq/Cu/EQDr8LXNivPo/xhe8ASpET7Hkk/oYek2I0GGSivIYF2t749QgVmyHEO5fVHnDzRN
AnMulKiaeGMvfrOCWj250soGu2WvuLakHL9MrsrBnNWrv8MN0BWxu/ivOTo6pfx66bZui/MFCG0m
i8mR98XxMfOXzYjBMX+GAIeg7BlGx6IYRW05KyKPYZ55mXYce6UXSiQ5AiVOpFylarL5nrLLGUJs
SNfbGT6lPlA8f1wyKq97vMGigqVydCelq+ifsk5ngnMBCzCXnVf3+GX17k01R7+j0en5X3XzM50r
lne1pTrt50af3dXDAYKQPC4giLaBjTEj6mMMtkz/gg9adhHHwW05GGDmFcxUW3TuJwpiTLH4K/xc
3n6wFTkTzE8aZ7tpc7B4zgh8YYKQJwupIclllx93qOh2kCYbEWat8ivTdWFd77D0EoIHJ7FkN3bQ
T5duDrdYxRViCapS3XwQi6gZimzGkMOy2UYPgjg5Q+zVT7ey14P8GoRmLyL8DM8/pebvS5Rxg5sy
fWoq1P6Z/oVp7YO8LB9prJGSyvmy9bK1/HktQ4ksvma7W/Xq225CICvxW59uY/VQKPnKlCvk8lGY
M7PF+n//j511flnzNuwuzn2G2IQvDQx85pEg0oDwKiW3kYGUFYWjVvx3uX23AIArfGkuRdMMSt/F
QaVwKIdzBmYjv9Ht2H6pLwxHfxV+d2507xZ2LK4vkRNa42MNsffweL02xMtDpx/z9K47csumzAhT
ryyLOW7+Vi53VZWw0flzMhWhcBL45iGrBxFOkNCKh94/1oi6rE+RhklLahDi3GUfr3I8lKuz1Gd7
vi5ViVBqpGY3gn3nX4kxgGo1M5rcEF4hZ6VRks6UNFTrNMScDNjxz5ubP1p8u073Xj7Kn3SgHaVo
HnvO/NDSMTrjhwqSlEE2Be01fkFtZ7e0bU7umbCgmppR63KGJxXm5yhKlAQUZztXnNRcbmK0nYc3
8UH9f3fW9nyhxXDfyr6dQt8c+jnC59WXs7YTDLNzqHFJO8eg9DP+CqXt/t5aopDw0yuObcWQybMW
CBcPcDfP4+CDmLJIznqzkhEQa4T5U9eQjXfXYoe7ex4RbsRVBNn1+A6fP4xgmZf2/Lo/I1xLnbFA
qnIk21EQH4iBYwK1EA80omdgRAocCKi1p4siDxfQuRcwuxvuy3Tg1w3o998Kx1jPMZwSNKj5ewPX
UGXsYBgQdDFQyc2pqCYTgShqq6O0P3DtCHzVjDl+UIh4Ky7xG9o4gsay+yCwQLxfQ/S+TtaW9awg
niCspR72JoMUWqxtcwASYgcRR+rHjXOu3SrC0bX/N1MwUYFsYpA5kj/DXKKnKMd0azF0DyPmF/Bv
B6cIMiSBtcdSA15NRzgVLV3qRcC+/DHmaGgNVhoqGYP6EHO9go+dtEL6TURTVxV4kIW6T0Yc8hxD
mvsTV4M0znYrtZpMQTiD8OnOuQwdm18cX89lXGlVsLMQxNyPuhJHUEIC6bREYZdFoCPYfATvxws1
BCebvVPZYP6k8rYyK/s8j01HuSFEByeWQhNkI8hBm9XzMj1Dxgyw9t6+e8J/TXWkGkXV84oQb4lV
XruXsMvXXq5EAXfwKkiQ6dckm6aFdTxdfZ4z94Si6q8zZ5h5CbE3cjuBKdvpLi/bqOtYpr4/Rhfb
NSH/QLvL/15ifIu0imoCsUh7qo2qxaUFoDdKyx7uR2rFt/oP37jg8EDAh8zZoYu10chm+++RqfPO
x1c2ss/YH+9lAsfffqqQUstTfyib8/UrORsGrSxyGfhIafvtfw4i77i05Ylew5Az8gJeomeFMF7y
g94fMs6ozIQRwUu4ClrTPz26fL4xWH26hylyINp1nsl+YSytDYxaxZf7siVY0vcKNVuHSAid4Brd
7Zb+/n4dPdbJoFI8wUx17Z7eAz76NFNFArSmp4oF4/kJEEk3tx0JcBNf/ef3xlQLZTzYPkyoIkhT
+WsDg5nFmolzGtIppZR2WFcFOw/xCV4cdWrn7F/b/gS1S52LX87td8TcbxWA6OyUAFYDltyZte4V
tucTVSvUNTZq2KkDnXs4e5ofdco+h+pYjGqAEq8yZg73vl88S41pYmPlIm1f7PY21MUMezbbB+Mr
WpP4gfFathll2gqkcdwbgsoNVXGnaXTGpof2wdUo7TEPyJ88Hwzl4HacaWT3PcTxbOXsuujznwak
LfFTExRSJ1iFnHvwZ/rjsJc485KnPh7d5qFr9z54rmacPw99ysK8F10XJKt4U4Mw+PgkGzupFGya
kyu+0IctdO/oACi67SPq61MzCKX9YnKDzFWl2wemd/EL0TuUhfvA6cwr9vQtartKzMxCJOo+3zX/
IUzEtbK+VC0h0MTBrGdn+rE5XwvZhSOgmsIVXjcCOhUrwDsMc3+6VLrtgU7bsdwcbWm6jPUjMt8S
HLj3+Fwqk40adgmYuiU6GUslNAKqAyJ9oLkqFO8EeN4wobMPi84rgzF/QOfOJsouon/BGDxtNBPq
dql8j8mqQoc1UoinYQq4fEs5Az/NX7sc1FcCNAMG/VPJ2hfKE6QzJ+wnH9Zmo111xxUH8vUiFZD0
6lMAvPNE+s8eBl30kehj01LbT5uwROJp0rTSewcP7uyOUPsi7eho2gBT5k3KkRcOFC9qgszwyxFj
O82fVmEltHTXCppEy84JQR4sYggJt7BBUmaX+mxNCt9miAM+uozvnT0Rs1eRxAzJCC7K8Levmj3o
FaeuzJCyUDTMZgT2o9V5+tZjtgjBj4v64un+eC8lUyCaQKzYST43N6M4ox5wqbS67fFayAw7/8hI
4Gvg8bTMfWSBXvypxrTjm2flExKXgtKmRTwI/IjqFj0kq30VmCVEfJHg2NBtUT08grOjtB+4f3sB
kGfyi9HZst+6SEpQ2XwCJ6/sgKuMNV8lJU5Luc9tMqsI5BWVpM8T5EzScc2z+2JmGFEPINaT5KCi
F0qDXrPJgJ5qy36qdcC6ATVg+2OcciFmvqQ+HbdmuIWEDrBG4x84h3pN3igGEuNUo3ko/d5zWOo8
ZrzOANu3BMIiwL4Khfd8yVRluftD49m7rrSTJymI4PAd/dSGkvWXcYqhidi4s9WEKlZw6i1pk9Sd
ZA0ewe4Lq5n2OeVHmzmFmyFvpjYiP3AVXjWjasf0V2LDbnpzW+T67zfQ243j4XFKbRseoHSSejj6
Mx1Thae2xwiM3PWTNXjLz4BBoejmCG/eJmW9yGKsZIYqJYin5DDroCUxZ1r6Kc58yVRLaIjlBLKb
ynzo0sQ3yDXMFM/Rmyn1mtyLfJccuPOgGDjuBlTNAI0fn0dL/c4cgJD9A31kRwbWcp6iFDIC9iWF
2ayDe4uyHgZUK9RnajbY+V/OjLPQzGezwekPIyrSlJRXBQlvGn63cVKVOQdP0BIneTpEz3bBPGNE
DilRAsldAeJIsbhRtD+4vK6+k4YZpWLedP/BPVcQqlNWcMWrPDR8un+6q0Hs+aIFknLkieGYrNLZ
5wZZf7Rq9azew2iwU30Y1iNSOawZPMGh90nlWRvWNuIWFLqFFHfhqPlzFfi3Vyh39wFb4LZFIcmW
JlL45yNlLnwdql6BA+i79PYeNnSy9YrexjaYtYD+IjiSwcYA9XHHeNyCYxAI0hb4wNeH/ZCrUINQ
BE2M3a6Sq0UNo8joIZJru/vJHZFhaNVNrAji9b13WvPX0zZoA5zcVkwstYJjZiTIY+GWc9ZOwX+f
7YudoYHyCDDRDLozIw0xEwwq4DZfTsGOAf5NENcceqcFv6w6NaHT0ifNrJpr9uqge060/Z+NChzZ
YPjGLQJSY2IuVCS5s4m4UdP+W+ZLTcvBZOwFR5UoCoub9F+Zbmnfop+okQwrLQOHq7Gg/2yUIuPK
aocSqq72awtvrKvpxzgsL86wvhuoDC2yBZn64zJi1YrCOaHLdrxqoI5Im3/vLcWY193ZYgbng975
LWm3EKaakMvEC5HIWjjtF68UyaGXQ3DHFhrMQlP827Y0E5sBfYz0PamjIxVm4VLt6aCHGU0b39qu
71+A/tcl6Fzh/E5e3iwSnx9FfTsV50mFdLwWz96Hh6hDouzbZNyHc5H1YYu6JN2b9AfKP+nd6AHj
fqZqqPE0foWUtocoXL964ibdYSjkIahB+IBJeiEPJgHzfcqoeGfE99SJoficduzySxNOm+y7rWkB
i1jOiVnemZFt1ELKjcNaiRI+587FS0/c/4lrOHKYQCLzLfQp6wt+7OhOBT3IbUBN2bX09Rfhg7E6
IAHyChaghqnsuf3gD7dOcjvsEfRH9lMyIyAAcMiAOZhQN4x3u6yr7d5YqNRojkLVY8wqUpgYhxTD
TlNUKEOooLNAK47GqN6pt+X+TIurtpzxPLW+bgY97+ppAaw7geNsg2bNDTGfjZRctg0yb23y6XOz
JtcXvqxqnh2AVmZ4+k3mU/BHwRns2Vl+ht1TH0MeS5GATMa+0/v5vNO259h8H3vhdENkNUi4x3WY
ELlE4TL/mPnyG11kff9bANngw+8hRJwuyyY7gf/D3scYhzBqAMdXuqfmVhu6UxLOxvAxUaJo3uAK
CrOXCvAqgsJKC/OkLnaNRHLA0+kckXmXMp3ZPiKMvtAn+st6q86fQbT5QcW77Y2unb7iui008Kno
jp4joQYptESPQxP8xv8Jgxb2rwLCtDwR5+qkvM6Gw7yzUhjbpcFzEwA4wWMaCC5/P6vQ25e738Cl
rptZzYMJ2f09EQtwc71nK7zUKxeoqQZL+f0r9GjQyLl7OMYiuUJZsaE3mvomEXbYivuxjAzijR74
RC5ANMc+hS9BmPMm+zzHLt7Btb7ET4I7FfXNWCWm0qyHHJjsQpQhkZu1nkmUBGxI6ZI+NitvplWF
sbTyabVkruERE7roFK1/xxheycTzooUjp84GeUfMOUONB1D181adPrLN55XOf0DLzTxyFY3Idu9r
zMeJzg77r2K+2bf9Wv0o2YhjUdD4Qvw2oEnxfxLjgc1SOX9fgJD4Yt2fiG02R6uY4POHS6yZYu6d
TTmRAEGeYMMFIEgGmHoghs663PNn25uHPpvngZUQCoViHGRt0UFnG/9ZDL1Yqtp02OR2/HGY1hWg
4xy33ecIQq6xjFXPk6Iidmfveq7q4KNky8uiWQ+57IxEI+w1DGp9gYDQfgTEXJ7cLRyedYZY6eOW
ZKZLAb+/pSoVXrPD8ewauBB+pptXHnRZPIwgW9mzpFVidbFBf35h0aBYJcpaSxWJcVjhTqLso1Vs
pjSoHLSYyXAaft/2VfIe8ADHj6PfgDe/TFox/FR/4SXycGG8PKHHNAooeazKy4myMk75s4Prvyxe
3laJrFjNghtYdLpufK71oVv4U5SggoQLubuxU93sREJTESYyZ8x4RmQXuaO43+sm4Ay6VFAiMWIJ
fTnNKewrHcCwkwg4EgDHUtb3odfpA5pZDuWbyh+u/+bkmNzsVM907oATziVQROw7Olg6/5o9lUOh
Uz98iwfhlr9GBH/GreZSKEHcbQkEltp4GFRQu+xyZbBWtJbm9q6K36t6+Gr+2Y9URtfMKuNI1zR9
LnSnObSLkroIPKPfqqePI322FoJkvdtpv+9dqUIgP13OJ0WWGM16GCsSCPzYSfgxsctwn7Tzyrjt
CQ+kGXFvVjkeu5mbc0p+5dvq1X4Mlmlh8o+28L/DXS6kQCmafQ9t7oNZIt+BYp4SVdHv3VtoNZGu
GcdLpvM5o0YAUmmwL8pCtJbfivSfkHMrXa3qgqxZNFHzTKC4J7fP8YhEA65/g9BTaxxy7TN4FSAI
dISaW6Wj/IdHjKC1k0nVvGCxWxQDdvwlO+sY4oLaGTXduwZn1GrGln1CIRDvXP6HeQi8jU0KB6oc
uebZrnKVqn/YKjCdpSVGPiyRt1XpjYCBUfSJf8rlzwo3kc3FzpZgiAUBTlUSKy4SK+fshzpfyJhS
iI8sGhoKkf3BHKaHuD0eyMjIEX/eSiSF7Pg7oDe2Wa+R5+MkjIfRAFXFW/cr6P4DykZ4o92rWv6i
rt1d6w68R+WnTzBhFmeYOunwdjxT+1PJQreEJMWrlkcnT5ZVmxBOGzl2uonPkqq6uOOOuUYyD+G1
owM58k3KygXxVIlF0Ea75vaLzG1Ey93qtn2LBsjPMwTT/PwwGQozbYdr69xtA88gSSbjMLG89r55
nRJC1gmBtd83DehhXVPaaAaIjE9uzMgSJqAr5y5IU4MCui8q0kHzZ6aq7H8ROsXZmACD0Xz8v3jc
Q+tGAG50pN96u9b0TS+U94nP9cHovDz7YTY8VnMwgqA2K59USy+If9m8UbU2WnRHtqfiHehAiklg
sriDZ/gD5wlvMgeVlWzGce6cz6J9I+/CCFgySw2ttezeGkm1pRRcKjhkWLQIiC4BDPRXxnqINNF2
hOz03bIkyipAtQ4Fm310MVLeg0k/Ewr0jvmLB02FFstemKAxRLDOVxfzkQ2Z3hqozMAqA0t/6OFX
+62KSDcxZOtQ57IGDk/Vxzb8tvP5RIo5Y5nJ1J1oGy7Bo7mdi9wafAuayq5iuvQ5GPx7oUR2ak5K
ZRa5lTyL1l3z3ZxaomCPe2N+ydQxJUEIBgnPR4sml6z1KJeBIO7i55LuyDncM0+9k4qonDqbHx31
uP7MwGjZE6rF4Y6r2LyK29Bi8ClXxpQppT5wD1+YW6MaVqikbt7X7lZaS8z2qE+8MD4OlEiZlXHl
ajrsgKFqNscx8pxR6BYBV2GzWblZldb1qJJq6XIENYshScHGlfoClWtNOLPW13BeGK5cWlVIk2uP
v9BUtG8+R3ooKKdNNvm4kf0kEqWxSzX/PB074TFYNqujxq2MuctdI4nFzOFdPhKb28ZS/ewxuwM8
bUY+sKPYguJhDTSBz62yCNSloPmtaoWHKFI1n5mkTocUdBnEpmRB9CkCS9Neh/s1uS4TpTlsOpbv
VdI+zbzskeGYVGDEHY0SP2YPaqSSWYVpL+Ivf/0bV4MBDaZQX568COxgUWA6cp6UY4lZENMaRCDA
d7TEQfFVWiAKL8J4kGjk6rMqQqWvILU7HRU/gEwureIEUqjAXqevYG+EXa7JkK8aVRTOrPIbfgjj
L7PclVP+YvVB9VB/wepE5IQM5zo8DmW7jSeQoQ0940xsNhULtffrfzxik2PTRUJE0VRunWGCpaWn
MGlhFrecVcgrZ9CQyE9rb8B/wkXP6ReUxagMuAztFqOVbmAZL95ed/+F/kxZzUqf0EeXUlqfSZnT
H/FpsQ8dryJGuuHfKC/RsSzxGTZbpo7qsSKxYe/rl6t0cEHabz1uEgf0+p0y7vrNMbD3/B7iXHUo
1uAF3FqIaYgu1/9QB3tCR7kHcb78CJSa1TE53K3QUJGEjymDCL3yE9S0avSUTH2//+Eva3k+GoBl
18mTU1lWT+x1dU5kFT423gZWqnfqNv2Smkb9j+hS1Bs63c8dAYq1Jun+YASfQ1JJaZdRuWwKzPo/
PxORSjGk+fn9eeJhYVowhTJvUTj2ZsqqwNzM1sI5IOHBHww4ZoGYA8dg2e/3e6D6Jq4mKEmeGd1j
PcCM7p/NqsOapbIgxPBxQ3WZtIOHkb3HlEiiFZab/Ka/w8iof6E8E1jLjc1xGmIVef3YiUAPIEaJ
+pYIXk70QgixHMYbZjY5oxPzZKQHDcWhIoUfKJzSPl8YlWxYoSFkaNP6n78XXbTK5M9wCHuqPeV6
/QQgZLhLzqpysZZM+7WUayDgODgP9Kuitkk5SVbE3A1R4QOobVEySxeGAndRLN73wrUHoATcUrjN
HB46fbctN8JTH22F23K++pItCa1qF4qoepALzv+kEbm5fkz0z38/194mzmOhBoxIcxZlN9gE5Mey
xYWw4F52FzyDwmWLiidRRFyU8t24jG3qS2gu/rKfHg8sCpwqGAlsxuSV9u0a60dgqNq2ZxOaoKmf
/Kn0JCwvKNgCd3mR/1n1Lmd++ZnQVMdNXV9r1Ax2eV2lLP8O3vjSPrLOJRD4+sbUVyxy25mpWdsB
ukNEa4auJ4wgnn9ed+VSXM4s4LGfW9eGH5KV9YyXkuF3qvifMEQljWhBjNGfEH9lyLMy98VOnvyM
T1Vjp3tnY4y+hf1DJbmhHzHE6kuQaUCsPLlWzhFnCjCE/4Q1yVl6k7LmKF24p8kDFyvQoJukHUdU
Sq7QxFhp2Bz53KQY3aihE95kmuOKPTJ8lV42K9clKVk3WK0dq2Tm2MvBVrTCXx47dH0TkHlshNjS
7uxlcpupBfgs+x8YijFNrIh6XHK3KhXtSqOuLgxF2T73/ADlMv/ypZdUyECp79ehEGfenF9Bx1OL
PHMyWrGPYwrtkkZ+xwRpBIxtE96aq8StBXQjekGLe7oRao2wjeXOpwi8lLKHY0fvNYGzULHh6h+u
WxE790ioo4GU6bS83zzsrR0LmUcAkVSrYBdu8TaI5wfwvL3BJNke5cS3eroQrWSQP8Q4GEm9LByy
mFtr35w5f0K8wkv6fw20QWVPod7+y2DX3P/nY1axjijNsNC3WsjC+Opqzkp95KBygYE7oEeeFmG2
sCYuRQVhGH0so0jDncbTMxIagp6Rmlo8ZnLJBXGrikpr1tct9X5gI/4HAU4d3k+BuEzyE1WKAsrI
bwJhBCJp1s7POBAHeyia5XXq5XbzXOHqsaf8iNsa1fOkpA28SAEN1MM+qLIGKAnrCCzBnC8vN7ZI
joCPd+Y6MR8hdmIbY1KnsEgcN3a74dcBozpOqd1oYsud9HpnwCkNkGu19a+yJV/Z8tLPOIQW58mq
TnOKZGHtQoze9r6uEwvVY+s4LGsTV8BzdhrTfkQr1DBrKlEBFGO64yGqXUY/vTCIDeRVcIfxdJcv
hybYMxMaFS879PjKz/GcfIRQwIr9BUV1ko3iprk9HVYjTMV50nixEpFqSSWapm+4hcv5Xv2LspHB
y3Xlu6EWwWrOJICRqlb4s68SSgUfCeru7AnqoGboMHnktioZYHs8Po0QaBF7uVuN1P7jhcHVHjuv
I358hXvHsXM3EUZu2gu4qFIV5ej5kYdjVz+t47SjVutymS+GPc+uqjbAodt5vxyrujJ4xtOE4uQX
MH3NLwdISKPSflNzl7c2zjwW20MJuDlZdlgI027Laj6Ln7ecYtYykFmiXBcU5nAO/Hkt1EtTG+eA
5WlFc4cw0Lh0EgOI1r4C0clPyjeIP2zoSrU+51NZ2bfnn82dFS7hxcWkUKwD4vw4n+OWbK/pz8d8
r26i08a7LPXBhgftm+mihuN3XImWX2NC7w27Yih071rHpqHkOXAaBEbSwewoBPhMRtWH84OyBEFk
dqUCOIVBiCw7NOP5/Iv4RyQnqCgwLN7CWqizemc+Hbaq8226UoDeR+vli8ex91I3ICsBR9w/vSW1
aBAURGouYMiaw7QyhHK1VjgZxUx511DVeXuL7Oa4jSmVXwV3jAUKvDzhTVp+OlPhE2sSHs1LM/Ef
yfuhhjoExK0XVAuUtFfwnAuSj+EBClpEweByP+Nt0tOs1+PXxH63tSJNAHRt3ICLsOdjjaQR8X0a
xVml2/CZ9UULc6GtKjHHNlE4yhR8x+7MY7VF/zOlK04IQIsB7S/8kGGln1HZE70B4R8Krk3apyZ2
oQEshOMLV2nIgBRo0ohCKmhO+Ah2VcGOFjyqfjipOrhM/NJQt3iZizE1zc+IGIZQxN6ETovb83Hl
PgeKQdWTQ1ws1hwOb/shYEwp17x6JA31qYgYQsHEOYFsyl/i9XgD0yI8yKfyZyUw4c56THLIJnHc
VpPs2fs1tSa0M4QzLtPSuSFdHYVWasHBeVxzQVUMLLqJggXiKa9RjgOavlQMVwfFcHTEPvmKXCQP
FaPXIm6+3sDDWPE07vynmYtW/YeYnSzju+OhCE0vqipo9Kq4eYcxNe60WfoxqdzlyH/Dj0CzR62U
Zk7whDvLtEBj1ntB/0UANl4l8WpBvKvmFcZic2kFzqdr19PP5czVjvgCfVfiZl+rq0kv6W/n3h3q
JihLZf1nCA3O6lwG/ynBTWt9fBjUH1/0n6upTSuL3gibgmmrm89AvF1DmvafwsOLQBDhcI09L98f
Cv/M2K3ko4kAtwSN0u5MDL62wN+l1oaJJ4MDXjncuZsXMY6SKt+bqdgtsgYgabLTj8cwfH/8k/Ne
52NJCDTAi00kmkFNoIq3/KH/XQ0gxaouOYdPwqZUTFGX4XrRYgaMRW2nVx+MsJ85g2vIHU5uBnWD
7jV2KhQQtc75bncogrOIqIs63+2iUizl7bfEzVCW7aARpMRd1iJnBC3JW+uXYluTio/duqMWgDlj
de6CP9o9GqlZPeCVZEKap2fS+RhcDXhXt8jYGmGhp5XkKKzWyNQwSM/ZswKeYH7INXJA2iHFAe8n
t6iH3EVIOrfboQrRLWZ9QWVkMZGuCxKZm6BpGRKXd5T5qr9QmO4xr4/Ywd/dKK1oHxXqU6oAbU4T
7LfV1kRH0H04EnjDC+cIxgZi1QS8hJln32YUbmTWhX/KxrA55CeQEI/+GDEMhI4kszrpDllanizP
FUgI5KcAoyT+MmsSvtsKG4nQcqYb/FGgHVSQ9ymmJvv7Va59wkv7VUo1tsHrZzMjTeKs1sbCKLC0
QREoA0gfpkQqN5BEKxv2z7Kb3xbGT3pfXnOJkCToTwvVN6IPi/sVEcJ2qYvw9g3zcIM+D4mc4qiA
/0cM9xVJanFjKeYCUJIs0YZinGinVwa2fy8FB+8jm/9yxV/ucgeKBuVQovUSXE6uaO9f5hMcGKFj
ZjyBcFpuZRp6X2P5xby41cpdR2rkHY4eX9W3dh5IF427lh/9tHJsTVLrweHdL22i2bFDeVefOqfS
p2sOGV5NNqfB6FHIDS7SCIjWCCv7y+UBIkLqe9IGXZnv2AAxo16x6K43fTk3/OiLpCekEK4rjHue
CrSOzAiFhwiTw8UQoaC1EdqeBEZEKIo1nVh9eH4Wx2vD5KLG8mZw6y1VFRTklcFxReyUeDGrmINk
j2BJDAAfZxLVU5ABknNqvLBysqEne3jhyI1zV8Qag0nggznDsLjAokXXwM7rwLJN21PROAGndnSu
pCHNdBwZKLbQxTX6uciCTY9/fihW5auOUgoZ0LRxfneVqI43Yy6et0DP0Q7WNGBglSdAlTr6D8Vt
JL0s7jypPcaG7zYjtV8=
`pragma protect end_protected
