`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
KknvL6SYSb5dRFuWP4AJqBhO3b64YXO1jXJrKEg0Z3ikGAO3obMtU40YwJiJW7ipQ08/Y8WRYNWh
nV2LdqH0dA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QLUbVPatcj7IWeOM7GaVpOxxKXKrfEAPdOAPmfRnpcapAKHnvWUhcysRYZ/rY/73FKWInR8HJilV
JFgxROZVCNWQ1zJhGgmKt04WHahOu9miHsfm8H7yNJ6k3TsDqjbc8beG5UCVgF6x/gDB8LRb2Vlo
OYeUOl3UjHyll8Sbd9I=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
N4fDulW+j2qCXqz735RjXksliYlPtal97cQEPC5accAQtxDw7TbdSqrHOiG5KctOIuaRzvRMOO5x
8R7f4K2bkMvIUjiiFP5Xw/fjJySLFuOiZoiNxxNdz5n6QQgBWYDepruKbEU7yj9zlmf0zEFmWZo2
ShS1WpLwP3B9Mcm5hJ+0GZ0wSeVmrvJEKp8kqO3uW6EVpKbiSMmBugVkGUzz9ZrIbzEZlELi+wJ/
HVgQM4hNwGKaRhAKNMJGLkgs6Mi/pI+CqjdrjRYK0X20OxPYi7+y3i6gUy//rkWJVRVSqqxJt07h
XfBm/2egXCeHNQMVyg/cuW80bFPZUcKb/tb28A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eEHF/HRqboErONr15dWGPiKIhHmEp89NzpKM1HVNOPxPMAhm5Q7SHcs30Gyp606YzPvXAWOwIhp6
yShxWJQDMNzjx8XLNdk6Hk4q1OFOlxJvftzg6IwFePhX6CX5M/h6gWDjhSncOnYuNt1s46FrBJGA
DJZ7AbtD39aEQbpRrtRqPKdh74/RGoSXOsksuOHq//+3LZGY5WN1wdVNJTew5IKMLtb98TYlHOO4
w28CobD4NywkdWMYWBeN1weCfLySyzftQavfk/dRUoBAG4mBbSm67pDUnjTuzD/BMIiEezbjKgGt
v5JKng8K28aaFylCDbrjWbQ4f0E0MG89P9bqcQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LBodvKMdQLsL3NITg6iyfn6uEr0nsFsSECbcpJ0VM9GPtNyhu1PCIqop74QUK0jX7gNod2kXTA0j
UPAVU1VbFsW+W9odvoIvVhgiIvptX2ncKxVnQVrYamDTZTPdFxs85ZcmhfukKF1ctZJMx5QHtsT8
/fgDo9EnaiAwUK6EH1vPn8nlJtMakUlaKARMU1hnWHBUkjruM2J062f3fYCx1Fc0yI51VXZXtNw2
A35SpeR68WKPmXnaWtRfYcT55OhdStBuASxbBHMItu7IQi56vUWP8LJm5L8r7e0VPvAGmJGTHM8m
DRb2QSYwaQDB32Ac/WNT/HueDTeVlvRT+cXLnQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RTdH2QVRkLMNeDjWHM39MNQI9JpZeMEnnaFqgJIEgBuj3R1/oXRV+h+0yVRQ+SMug8jz9no0jCSS
W3wRM89ooYAXiOYt8RwiQibqZKat+R7T7m3thhmgMEI8uoi9fGuXrcwO/YAOvNwNOuRc5iytwydq
EbyW4aM2m+CrXKFlD7s=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hNd+z0nXH9GYvgjnhDJoJvhFhK8AT6oUoCmTuJoXrdeSPSICu0d2AmfE/9zKTVob1byyZNQ+dZJb
Ma+7SxXV1+3xFvececBxzrOjVMq4geH8T4yeo12KR/tsEogGtiBVtNuwOoiOTxmMqj4v1JDOa2o8
G9PU/lTBUSoEzibdcIpQyhvP7Mdz6AOWlVWthHuCNvffk52oBkFkYg/wxqRli9uZ+ljnrd6rXIeN
pcjEkI9ALbBEAZnGGMY3do4kdn+d4UrzbiC/0FwIrw+uZYeWK2+A1bCZ3JcBMczd2lYYJYQOACWj
1dr/Sij9Dnl2NTdY6Acp6dQAwn2oASr3Hs8Onw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3200)
`pragma protect data_block
F4D6nIAHG9w7CzDjTOGl41ogLfBDzmuspYZSQk8qjBrOpuucVYT+diiwlidT+yzFw31JrhrxUWc0
At8+IxdcQqoDHB7xEf6RivHeVwIR4tPA9dOMVXaVcf8VTTav6EVETUT9Z1TR2imO6pt7Ojhgs3LH
tY0OG0Q0VHTZ27ctPEOylwm4+mLbBNHDz8DGOnFeNrrsxPOCn6Pq2JDQEpXG3QxY/XP/dHPj3NZe
kcDtohDhwDI2u+3/htKlPt5EHWMmYuxTrsTf2jzlDbEe4UZsBJjbg3Et07/bw2/DuEVOBDo7CyBC
/whd+auwEri1QHgDslwWSYMgs8E3xt+5YV58xdsyVgPEu3L6FQvGcSgdCizIyi1MQFgRy+x0og4T
++DcEsPChq76SnSHIIv0R5km6ibsZ22U1qKU8V2l8cuwZPTme2WdB8UgGocRHQjuxBhLJ8Nsn4+U
TzfQPrEoMswwtZyrNb0HRqJi9agCdXfGS9PLSNobt6OT8VAEs7pfftaGj3Kl5B7k4B/5/gTSQD2i
cPWQ836VFUAx6yLdB59CUzNphyWcRsqHjBbNpX85UfXsEpbBCz0l33LJj30jNSg7V95quAz2tzSQ
jpBUa+IvToqwY7dPNIIgE/7WOP0BKEGk3gF5xtMbV22y+WJ6GgXMF/itWUxumox6zH+0hZ6avXDv
XJt6SBM2o9su68pFirPbTpKwbEWr4YAM7NpF/5Q29RyWUnaSrRq2Og/DKB4AJqOdUrWVZkmocfRg
UMiDREDmgx+sOcytLmGJ9BJz4iOtIzJ5dCYX+v+AMPLnhHwIACZaXj+Qi4liZSVWAoo0Rln+hGBy
AU19tM7fWUco3NzR+doljj18XeqZ+9NEmH9NflJ15kwxGeYlGjQr8UmMdmpDCR4WG07BS5QWv2fi
4hcjd9sGRsaRIvlh39QgUZhuzS1gzjv9ZuYijTbw/OtZiBgfcCgT5OFoFWw08jHXH5xneOu6p6Xt
c6KLC/VWnQ1TLQDM3dOptuDAITbwKIPh9ZfSWwvvyw0yUKIXLAeCPH0tf8chXacRL0zHRE4U8VQl
VelF7tRSp0LacZuJC4n6zlnBXdtUDCCjOMqG++93IKCRCROke2UPK06+UXFUAIn1CPUpgiVbXJ4z
iwZa0sGck4o1SmM8usNE5lXVK5O1kHLn6DMvWFIUTA5S4pcFGPL2ux+4MEFDUZWspa6CbXuwEhnX
1V6tuqx2Vm7FLyJrlTpMOsD3DXuSW6XOHym7+lu5rZH+CEt/x4uF7IA2tm960vTkaovQGtmlJx0D
HgQtAXXu1D4zL7vU3V8C+zGAOPEb+7f/al9QiaFW7mBMrLKNhE1n7mz5djXWnIh1ZDgruqBFa879
aZlJ/chnELzK7i9NnhsOuL1liaZ4QbZHC13Syp6J/fYeBiZmWmmeyLCpKzNnWeZIUqfgQZf0SH/w
/B0HtpfksSRbj+82qZJOQKQbcdPkqs4jAcbwpnRVDGbSnJUIJyHHpjbJegtWfpVwRcFNv+vspXo2
PZPDjloQSdpBK3hCmW/U2R7kTLZDzcZOH8xC+fDa9awLWzTdK/wJqBPpn8M1txhOlGaUA2up/68W
SieirEDrd8xNPuLY0qLBMo8+/EEaKAEkB+NsfOeeD56yF3iavizoM0E6JI9yhYhf3RXuF+gKyR81
RA00DPQklqcNi98spWiEeUBvHHikKFYK88o/s9YYhIms7oGi3QXeFz1tsPTSqum6Tt1jX/YoiyUM
y9d8rCrzzSuuHKZlCkNO5KWJ1gtOyJf6tWfaVkOFi+X2R3k4mWLuq2/gKlIRWgGVMjfKFKbq0fTn
aD4K52C8mIXExOxdNBkKU4/eUggPWOyuvZ4UcRPsIGIBTaLTkFPeMBcTPwVxBvUebF8c1WVbYhFu
VcVz5d+9m8DAUTRZ2ajUAVo9zcoq4FCDpggWdT35MCR+8y7Lm1M0MOFoSme/NBFCQQxAcfF1ww7G
mmO4eeqqC80lCsp3cL+vgU2g+OtrXgj8u/RqACj/fEmFZjyybi7uKt97fi16MLhLzd9GxeKz3jJc
DV8uKTvhOgmNneLC+9G7AkDtMXOgjmdgnF41AbPKuDhFXEVTlenTYh5/Zn5MaC1m8G4OAXspX2UE
4RzyPHrTa2EP7SFKGam5y+2CqJexMgxzS+sIsv/7mHzWDWmc5jP2hWVvEnwAfvj4FPvy76e4De6x
4M+UPW4kLZGQj1nAwgD/R6Q4ZnoWj+VumiMdLecZG2vtrcTQx9CakiJLFHsW5JS+RdTKWyth1v0L
SDrWNVW8qLJ3k+NjApyTBK0qWyQPi86MEYybm5D1okOtQN2qgj09kvuECadimYvOrua8MvZVWraN
2Of66653HIZnnGv8utCf4g2EZa1lDK//x9diW6f/6/ZoVg9sAFz3c5DNDpAqNcFiAdnYkrliEXdX
NbAjO5DbkMtdndN4ye+cbvADrepExScvc5trPgfbpxt5TJtrhd8Lu/+kNRknbIFfzwzdNM79Inbq
TPAxSlKf2Zk5AnGEIeZAZpYqzcB44YAWdH6M34/oHuUKRlEW3xCYFPIDz4EodBjf1A08J/blWAiM
9PpEvlwnAfYlJhBQt+5k71DpfXdMJLwGYbwpefiKVurovRojR8FGwESYXpUIb82sZQwzcQ+2fNl6
E9aFXnWInbgWu0pgt6JBYoy2Et/rkYM6Yx6MHwfdpYw+ZKwV/Wumu7xdUO7txvXw1EsTilFiwS/N
hS9f+BH7X6RyZYky/7qx9QAPVVTKXE/WsyXPr0sSVBtFpR+1Oh/TZG0PvybE65jlurwbnZcI7lw6
xQJiiDvVR1DeEyGpBfHdZC9s+1p0gyUZ9YAsJXLf49NwrWcswOFJsOFXGrVwHeG11G2yc8UtLI8Z
EvzHM7wCODtugyQ0rUcT9N1kq4TmsoVUHFUONweJXCGl/EpOk5vJJf7Jna4qJCWiT9ja0dH5irju
cQhvatfcL/JoVeRw2/2GPPqnyWb7ZxGlmDhv5cjIMRuyjXWMEz/LKSLrWGzI3aIvcXA+wu8bqDob
sfdc0I3Mf0Yqe7YzkWnlDgHXG2nVOhM+SXs8Smcnelmo8DaGPM/W4CJwGFWnDzmuEfdV5yhBGKLA
cQlN4zZy7SP1zbeS79M0cK9Ld0uGXpQZOMci0RFw2QvgolrUhhtRRYDmGHrBgIllDLwkNyGfukaN
PFds66EG9R8yqGkhpqcunCduju8e/fkt2vnVyL2fGDcoOOBWaN26g1eVNtkHiEbRGjTF3fiYRI9U
M5SgteumaUSuUIYOjhjD7ESXFobvN8r5tYLuCaWK+1FC5Erts5IsOs1VdnBReSHXFnBrvb1D8luC
Ch5qVYZkHjH0r7nrV8XedlTHHDCiJ/QFeLZkoGVa1HX/LTl+bwIwQzDcssUCdJqyHtcp6XsJgJWP
/2H8bwJW7nlrn07rsIs8N4S7dGl8hDv59aa6emFMNqbQ7Lvgwq+CHw8QW/Dle+6LHMI7ZpKo8J6K
BXsmKISS+PA/eWWdBscmX0XMPXva6LOvnARZkulxjHjhSq8NyRXB8SHuRJLLBtvd/MeXCP/qeXy5
kIoFT/JGJWrHMRdsFzH1II+SX89UUnSKjoS1QB+J8efNyutPg9G5yLooxwEIn3Dmt4vy49O4ugMH
C5I6/wyG/yPVpWFW0/mJ4i4S0+hZ0SCwrkPmow1bpgwNh4GAVcs9uHFLGVCgPgLhCYAVmB4hXIht
0D/zLJceqGbw003QmTbUNOMfiRDGK2lOfyC7y0/VgnzT3MZAlECxFwWwWDSs9dKXpGyp9wJN1SxH
jpj/173CO0Po1qaprh5RM9KgJAsK/tuFZJvxOfbPWkRowZvg3zhSvv0f53yKmvJX3o4GntcoNSZL
nd2kSUTEhbCkOsqWt00B5SHx+bG3c100hMcZteLuyWgmO6fNuRtb+0m4v9enseWKaCy33u/mAgi0
4P3auHKPtZWfIxHUI6u1q094qusm1Pnb3YyM6lIQ2i8iDUfnexz/3XLeKxQQffXowYpoPwAs0GwK
moV5RJ23gDtnvYghzxOE5czWz7BVndiYL29/uAdils9ufsSijHCUetmgMheFnDKWcjbsaQxhMrye
u5CisU2YkIzfLA6lrOQKVcndSSfzjEA7KFvpkHcoDpcmI/tsxria478dIs6fIDSDfeYNoptjSfEA
K5sM6A+Nwtlgm0DO/NVMcBl8V8ro/xoKIjJoUSM3OLUg/kiTOZZZKcR6PSzdtyhptaGytBihH/Fn
rde+DA74UZ8=
`pragma protect end_protected
