`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10144)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qFsoQXy3Rb46uY3SWSugoMr5v4BWbdiGa6dprhYdL6h0bJnvwuazDT1y
S+A3OMqef1TgZUTM+A4Gflp9vNdnIuRWMNlRwEEaIseHBq/RHMEaWty6dSBD3jkQ78ycwVdbPd5+
UAmZnRta5uodDdw9UOrGSigE5Xs2oezK3gd6oj1C4tfCndYONzUajoRMrXealp5iqfc7RmEPnmHJ
Ikqf6z4c/VLWVO1c52tysEfjnH6SRaP+PIbAVbtGauEGGrmEvU3iGf7KmUJm774rHEeLUJiaWIGo
f011jVZzS4S1/YTXcK4NpVmntxfLFRmK2vYJRhyymnysL47ysjeJVsJGmwa9ljYKk/yqr/uDuyP5
CKmi/8tdcYqm+p4vbg0r6VPWrWMk7gdybHWB1oM4skI1snwq2VgGyroEXBYFuov7kiRXScCmX45J
DpvWR9gXhvoTqtBka7mwV6G+lgvDEmCji6vHrr6dt4kw70hQpyASPIx9gCx+6bYqUMxDJ4abm4yq
WTkTfgQY70ia3SM5x6coUnKS+IF6DityOSkIwsgcUOJrWxJRWwrQwMw+K3GnZWeqasBqd7nhwN/s
GhRT4G/o+VwBtha0d3Ec2nI7LJKp7nhdy0DsbQGRh22o0EoS4kr8379KOA8Au+yqrsQr0G75ttw+
9U8dIG3rim+dDBfLQHkwIFxd3ecBzV7LSfkhaYDKebx6EYsdOUaTF1GhnqhDKDRvWPM89eFdwpEx
anFVIYCW1qte+e2/PUMisXm2X70vStsaLZ1pBVolHUJUEx5QpwNcBTeov332975vMF/oG+RBqpHQ
sqrRgauHfAmwlx5AzJRV0BpritMTZN5WFl9BRGnl0msR4vJ+TQimh6xCN4YRHL354a99BLxcSyIY
ZODUp2Azsg+2Rnwzj8KQ3n9cgPd3VZzog2O66dtLm/WTiQTS8VlSanbGLT523FLS98u9Sh3zDZVN
EHVPI0zT6Hqh2FuDDe42oe1V6qoIL8Jrcyjxxux69kOSjytWahD+0hLeZSDdGIenwWGrgTjWn4K2
qQdlvuZNvkny2eDAsiM6D2ZBKMb19RzQrhkhewKAnIiJ/AUxhkgdYWdryW35SpcxD08ce+kr1GOc
qY21hB8rWlNsd5sib8pqQ1BBf5rbfwEs9moboz1rqOgNOu+SyotrEog8XSvKG33PUkNf499PaTXR
q098RQitbIgbHY5nN+wfy10Bv/vKdtGSpQxig1edHnWrBhnsBUlVW7jomkAHlqjIFKvZm6Lt/IvA
QVGXxU8XZdlnC4Ll5IxIn8gnH0PO97sz/EGYOEWdKXscHNNaar73v6/tuu+2xG2tXTNO2Y0WHayh
4vxIK8FCnsZl8PgpmsbbaQ50sZrDZonX1ZaFjEqNmqQFlbccNqlIDK6gZYho56EnL7cEW0UFHMp1
RWKDlKalo2fBhMmdjzneI4GZ8xFLF4VxpjiwW+tGBH+6XkaTOsPr5ireTvQ3UX31GgCNHXb0tCiP
r+H3iui1aH3tyWdjzIfgK3jr2AGNpQJ5YUjkiSfpY3SWTqEs62MZa9JRXvbABXX9C1duOmwKtFTz
NtpaET5GhLPkegkgp96yWpenpf1Q1zIGOATpKUM7Bov4MNuoSIni/mfZwv1Za+msb4BW0uK6XdGX
5VQFOiOpsy5PyOQmRLY8I825MTsfZw+7iJX4Wns/gFgJ1URzfAzcu+62n/ILGPhyymmzHVgswpdK
pPglCnnT3Rk4VBPbUsMvdYRT/GN1o3Gef64krto3rBgbAEyg6/OYww4o0cw0/FhYPPUrUixSBSXq
0g05GQ9+Qs4V7d9fd+JAuMxgw3Vez1f4r+iicuc5H7iK1737L/Fd6myR9mPKnj7rNRQMTDJ5yKdK
rWIlsStEIOlWdNy3AOCk3gJRfWDtoS7vJbi6gG2FOHIWABxAZkwGmNbygway1LtlY5ckwN+aw8j3
rdohviNKVVclts6Cf2xrp6P8sMlHKg6Z+Z48n+rGNGulOYtIRifhhBMuFs0uoijOoFGHsCEij+M1
iR0TMfnPGgYjkJT3scz82T25ay0tH+cMggXvn+c+orTnlL6V4p8dx0ZICac4osiWpNFZ7bT5L/Mv
x8+aitr3iaVwNfRjmVmPOMMJR8gxBqr66k8zNYjM5dkvRz8ack50NIUxS/cyz81e2GuXH4AIEpNV
Dqklx7VKKnGluQD8jMWM0Qqu67mqHvpmas++QEJF8kVwGX3A/vhm462C0ORGjHQVIzHke5zs0PU2
lhRgYSggwfC9D8OhipzdmwKzDp15efvpBJuZa59vuaZnKmFRDsWLm3taiHJuxk42HwB+Ldp0CV/V
wjsVTLPwh7cOl0px3XgLWcZoeCM3Yz542uK0nfJBzZEMtiCseSKUkGAxcYJIuZSYbf977L41Yp8o
o70r5+LV9B+CRlDTkT+G0Clk7njGfuyLyXkLVhMgesoJ8jvtuTmu4bsnuu/UwF6q074QAJAngfh9
FoBKdv6PYA0H6LRMoecEU7Tz3Zc7LPvxXVz6q3VhmGYO6azUOT/UvhMaFflGu6GYp7SAWbcfU5kK
8/qC86V1KEd3nuGd3mL5nCXHNDQ2scUSP74VhpYOig7YSK3cpkC5YA7NI9jts+9iTIFXe4ZcPgWc
3EnEQ0GyYVRGdYkr4zU6Myojp5HsYYykNxpbJi1+mMQVe+3C0qJT3BabtJaQh02m+d+l2rqzIHoO
zAA2XFFWb6T3HOabhbiLujZzvNkRzWktidnWroYPeC4VX3cgdS9lg7vZqpMtHIlCizGjsYXzNBBi
wQq+kWdkeywX2R/ltedOVmwLhiqg70LdKkxLFTR3UhTjXHvDoZ3j46l/Yt9juWKdwebssXDd9af+
EA48x3hp7rVbLAH0WsCBza/W3b/I579wH2gbE7977gGZOaTnlHwzOxF4EU43WCNSaQtfBnNKMSB7
lDtTxXmhnULez8SW+ZK23ZGB8eDGgZswXaQEwwlnpvBMbTGmM4WLjNOuEAW2tEFiBT6c0GgQoil9
B8mXQWfX07m5KjeoOTjZDLmOUFGUpNzHkBywhLnj0cfoQ6tcady6nc6PpYM5rni2GQ/jzBZyRWnO
ETb4ZLa3BPJSiB7LT2ApGb+ENudz6uj5yDdWm26ncjH7E+276DAIomnNsrTmWl0/iRrVTc0D8URu
jJc57n8ZdFHCDW+xuBpi9wAsVPin4c1Tk8tnYqxAuwQAurFPg4aPQKeW7OPwImXrcZc5I2+q6kxo
qVAN+PofNeDisUDCKFUak+ZRvhrK1QNDYqv3n9bctWDcorjaDakWeHDnY+kJYkuptDjBqRZgrQ+j
x/d2RN2NpXXeLnIZSmk948PdXRcUEAdICOc0ZFGE5O16KJSCcXn0nttf0IMsGAKUGSmv8G6erlHR
VbqirGHSb8yZ2B4RXg/PctGChGM25ZZZFHGpPSk5v8qUYFeT6Djhw4LOqlN8CIs8xll5fXKcU9mU
lo05cvfPCfMmTk50ctPbKpCjnXml4gdwakxYPMdCAnqBSvthwilPgY+01+Uat6icSipQZGnUIqaf
vhtl71ailiMC+R85rMeaBv8RY43KpvVIHxKs2hbFgLVqvuaHRMk21C/8YczqY+yHyUR8c1PuHw47
D2fAU/8UHnY/5w7LAv/co90hd0O0pVGxzHqES1DmoU3AEvVhteDVj1ClviVMxpU+VcERP0C7C2oW
X7EPf7tXA6mRliWnQAaho7/hEr6GjDWDwojM4icmI8zuB+1DasvkZ0+25fVJqmp7i0RU80o31iQX
VCb+C047BPkKiaGoTVQAmp88Bg0mK5lkY6i0/cgwaGukm/v69CNXU33utcxn5xkbBY91ZtaGEoaN
YaVKJ8dWa6OZKpEPbFOpFCT26HDkogAuFmmpvJfq7+Leu2ueHz6W+ZbjtbWkCOP9wMekmZIJN18x
y822kkhcIPjMzYGusUvtg+sP7tJyYUYd+zGXWPBJyWmXB408uC/r2IwS5XlzzI/lAgIzYfSwI5TU
WY6ww0Re4pPXmJlLQAYfsZFIb0gsQMEnartNIDrxla9ecNg/hGRKr5qzR7fkzvwcqCmlubWEB9D9
001N77S2Vg+GVIpkqvfzjaQxfFwWqh/jrB0cj8xTwsNT86E52qLfF53FHKGfW3qzBYEGoGnH8/z3
hqFvT24a+X0ke7DajCiZnLGJF0ENaVk4AdiBA6eiQy5JV2N/CqAKOrgRLxFIEfJYv7ic1SD753lx
um4VUDxnsdsFq5rU2fKKFqifUnHacn5a7rUXOLyE7FgYVBOcBaCUxFDHTyC8IMN4bF3BaNSOW9jF
osn8YxKvBuVcFa4GYvfJ0FtFmR2b7X7xUwJ77QyKMYUc/TEZvXEpegX3AtpBvaldLNFvsxUta1aI
V+FwRX/jB4oWRXyARKHsziIe9V0Z/+z2lhD/5GaZuZBnxhvO+TS+MPSaqLBrh++99KQFNRpz0iDL
9KrWKJ9D9y57KFmTY7oKeSjcwlAbqJR8aY6nI1udy+MP89STMN0bkkcV1co99p9JsVvECP/MvhIC
I9TB0Oyl0Naejy/rhleiOCSyiDYPFSijJNiZ3eiDiOZ6bZNZ2CXzH29oazNzvta61aCK10KHBEDb
bXElmWAZiELBFMSoslQhYEJoyPaXTDyTg/YAu3mT/RSTjlGg8GmB+6/Nvf8HtOOWCc98Ymt7AN4x
yonGtp+0Fgxf1/0rrIWTVPHPyE0XImpyD5Njfh17PbpDvjJwg9gV1KliVbCvSry4kryY9/xlt+jy
eKZbB1gTwmJ061BlpTd84FgrvOrLwnOJMUozxrPDuodKjnGoZiHF4HX0ypI2IzbE/Xc+MwwZnG/t
1m5GKRaJLwUYbkv9R7ajwdX802w1QA2miAKTvs0pcOGVZ5XRIsltYoOyVP4jdi7BsTQyYSm9CKLv
px79ou4D0vZBKAQtNY3N3/HpPS6lbRHUO/VVMmIGGnm+UsZfUtHnXKm9OavCL5qp3m7E2tj0sv3O
QblmpyQJLV+p3Ha469JyLQUF2BWC1jYmxG81dPOdN1Pv1QpKfAK7TiSyF+L2M4k+oAboHXF5U73p
mjCYlbjSdBlQq1h/zEJrEoK/tpkNQdP2dGAwEwwxrKo15rGM+iLU9imDMyvVGxWXUvAKXVvsPCoG
vHaa+i7crgfRXtDwVvIVqpq8/4k9OoGOTAlrUWLq0MwQyHGIIvNpE4YruLKxirub1cf/VL7gmqC+
7+wbJvUxTbxhtnBrPhYmh4oY8ZHPxRGNlLh4BMslmnJYvUqBVjPt3jizs4hqSDDVUUurq9K1Pujv
EBxxXz/OZagCuy4Wo378vVna6B7gRG2pqdxEEaY5rEeaq0HMZ9P28YwK1oTQMTgjtm5hBkyhqona
gjryBWNtToLceHlJUDSClohhGX0+md0swEdnj1Y5yKxt9O9aKM9Gogls3yu5s3d+dybkEg3kDOxD
28WYSqGlQIbOeXaKIPybC3MF1Z9rvy8lghGtMuJPJ4Z6BMRiiovB4s6wqgfIPjE1jq8gb0FhHf0Z
hlqGrPSQPugps2TwRB1FzNdqKK99PRBCx+nwLIBGjUsOv8djVBWLuLOBtLDdXFYUW1Ok4gwSbNEO
+otw09MArvEhLMdT7cqbAgwZqTKxAk4mu/zcTvhR1m9BFWEUr5foGoOJEfZSwWIGHp2kLfQ/XGxJ
tknwxM+d2gW17lyT2EvCNlIVql/5cB/NATZVNo8KE7ittB9DFDHEUF3RTdobTRNsW6ciu6zflIFv
+fW24zHZdG7mAJlNHfpz1AEmwdVAJyDdyg/mg+GG0W9L0augd9YVmjIZchoD2FYik9kdzgCW7wim
Imf9QLAe6pYswHHUT2If+o007m8nkF6Rnl5QpLjtHOKxnjmjnW4ZI5UhHn7vwDFaed2IzkqePg+K
AwXpVGWUFEMdzOKWhrkQdN/x3CxAQg/+wL3Y9n4jnidX82yfAawrZ6V717cOPUu8IuVQkVxaip4R
2iv1ODKwPz7ca+FiYTrjEMhjV1iYIL/srbofsH0dq3Fb/LWzlpGGzOQiSJsg8mZj9ldrd/LQeoXK
2HIEDlX7foy50MqGhReFZeYxFst/+bOfF1FWnJUPkgYZqcdt8UCioqSAjyoBAJA4lbpvIzyBoeC9
/qEV45EJmxpmIlaTQjx8zjkfGBX5jjC7Vf14PdGAu/G8rRD0xH2IDd9DJuO4tKIRe7e5cMLwWXqD
pgE+5dhz/9orSALFfWlqlCn+qX0F82awKs88abVv6jhuVkG83U/Clk+Dh8fTIvWitw6r4pwIT9QN
ZbcPiZG8C3aa/0WFwwc+DqhC2Z9d0r2YdMvSHnmJuVtuzVvxW3KCZWIC1x3pJ+HPp3EbFflFDX6F
A5slCWLsvcKLVat4eCsFj3w6vF97xmEMWXenHqBH3Qn1sGVq6JaFbh3ODnD90+/asIL5XFa7wXZG
/IsfeLjsu9XxtjDDsqpYXFDroh38D2nSmTD1YyiY76JJ4O9UpY0QiXlS26mlrq2byy7UQ1A12dER
5kOWuLRmvJnVcGDTnfeZvDpuTLNw3tdlYj/ObF5+wrG7iqDZ2rfCPokH1U7frtF/Is8XH6tC8TPL
fRNjdeIFmkHrb3ARxIlneiHEURW6h+zkQePZ2fVevaB/pQMSx+dNQkRpw3mgH+U27/J5Dd97g/0M
bQa4uKL4xi28NYRVWEGWnZxZDspYKfcuEqOZctnxYFbnxAf4Ls3QzUkgiqwhVMgyLttfXu0FNAfW
KYQaPWll8PTJqFyQ91i6aJVivq7F7MPJwaxaGGBd+4MCz6DKFuAyI/wquOQ8t6ojNSs5pTSjBZPs
pDDjSAv9g7fam8lIdCIsQy79vHjhKbtRIR3tBMsTx4rLKPPbEaT3aYFes97xJsLfPvefp3+Hf+3X
+cWntS6+x2uPY7yLv04Btne2WvmuBRh1CkBmvXj/0aVNRI0p3HvXXfOl8Yghwybec+uGAdYlqvyv
fCwwdOtpJxKhBXoEH+URcddBLTZe7Q1zJ1USWiDzMKHM7NGrQbFqJurYhYDZaziYsDAzRkcEXnbt
P41orM65DkiAKn9+KXglK+JUXwJo24nu6eO96Cy8BscJxKtzmdGXlMD8Oey+TgYFQHdXrNKj35eL
bVs9s9hPjRqySYo2jeKtIcq17b0SJAqJE8wlbhZnD28M0paTNjpXKJgSdJTSVD2yBZJuBotQwYPv
yK6YtpXSXlEZHZj8FcnEvLa2iUXhBB75jr6vjR8fFVrVeNEA+gImjYmag4e0bqHwQdkb+g9ytct6
FhyQnkoyowSGzRQZo8nNsGfi2b98bqu6BGWkHHAzpN+DJlO7rWfjvSv5rSaOVVMNcZXQuzpTnAJG
d9m1J50D5OPyB2BUubsJ/mNTVSTIvP1ORJELiUnBo6xMs5brIepdZ/HUh5ckBgBW7WX3nkogGi4m
gBayshormZ+EwCQcJfzPwUIYqQA3fx6Q/FIZgm9fClPLWv2NdDPyhIkeb+Q1gRArqg+w1f/5G85L
4/TCwmGZ+DUlxSKJnP66St151aZPTSbKgo/X3+nGUzFav4etRL8TVt7YvM+eAOPQgbPZc71XCI6d
hwr5UKYcx44ZUfQFp5LpWfyIYR8Vee8dlOm7LWqDJ+BgT9JijDfPU153a3+fa6ZkKPjyiCRrEQVK
OQb5Njl8L3oZPlU83OqZl/y865tKrGQnviOLpX0iSS+ZknzNsKFM/IIepR01KOB21Jf5D4xi2Ygk
RZ+os4K4Kgpt2KkCtrpZLNZI1jXYV6/jEvSTmUAJDK+PDlqmmnY/5fRC5XOD933QhzBX/CbgfW57
1ywWIVmKKwoF5+/W5zp124sXFoYprQOcyvkBZmWQ5gZVE8q/3HrWnuXRpxVZYoQIr16VZUiIg4Ot
QtDVSPZG1GKDOj3DQEsWoXZNc17jPs2xTLwmEekAAUWZ/6vifP/wDp+kWjJtEA0wwPZOcnAKdjqw
Tk7pu4yRM4YAcRaUvgTPgkHEISw4uhAllHrjaRM4r0fjOW2j7ya6tWUn4sReL5z6c4lTx3w7l5bg
2T46vZs7oUs6x2myhZZWFL6pVSaQfvg7WMp/LxsOL6R+eK2sblamSv5Iks9gxb5zz+YU9ZG3HX8X
Uy4/tCsa9THA5UtQILuOhd9Wa8W4gpsVvZ+HVG5ws+uc9yNdQDavze9DGAjQTAuoBUviOrq15G7H
aksymKuFWhvipJB/hGws6cyp4olMuoWTf3S7JW9325MOiODW2ZV0d65sVFsQnPgPSJ4AikwrFLfW
GGVagDQ0lBHhneMUEnmoIG9IwUXHGlOjqZnjjGUxdHRPptlzUeMENV10Op3fblModKse5+mTEav+
mX0h+H9VNEy1raEo71nhW7L/2rMefbEuMagjxcumqCMnWg322sfXR87psQuXqbP2kgW20mobrhP9
PvqLDuPYWCY9LFn6CJvbCWcKj6ExLtC1nhDAPIy5avb3VRgMvherGAYLIegidvYkhhUFYV/6Z4yn
k9ZV8EufTdbAgKouFRDW3jzNcxBJ1usX+DJ5kE4z1jaUiGi3Cb3pATi3i6y2kXz8szHPyImXI9ii
j1NHc7rWZZISfPUUGAXSizUdfUZUcjInMglrYLkCzoFVRgO9NSRrmO5fWutk1+cQle0zYmsKuCKA
VA3F+QtFkc7QNolVoQNWKzYiYDcD/Tl9KUzMMft02EFa9u7CUu3HrK9spNTDui92A49x9Ue3HQwI
hn0tJsEik2AnOrD4U9pReNJQprusnqrhtqNe1m6JPSTun0WUCJ/hvja1/N/x/pDYlIbPxEsvQyGQ
Qe/8xyUhiHpkpCHUiWlc26/T9HJhwYYxw6raG7uDd5S1b3kqLFyogEzRkjo8P1Mj2Uz6VljX1wB6
vb6sEONY7aygcuQnvs2niB2X/ii8Uo4Z/d7K5u7c3RC5R2dK4VUQwd7QPRgZtEV5F8Jroe5PSYIm
muyGmfE5wahNK3/Vt6LlmEE7rxWMs1NmUZfV32tPO3UBZJTpVPHKzDWd5QsBuOPIBJKYrH3uAA1X
gP6sgLC1gTQ5N1T5UJkgaZU3z7oJALMe8zKbIp1jdXTNpcReLQfUjgm/fJtpX65QiuCbSnOZQJkh
YITx2lc+Dsxq54L6Ww+9UVkzkQgliWhlvu+BaH/TKHu92XVbHcBd9IRL5bU9SozUKF+piYrKdqP1
Afrlbd5PBJWuCmi/AUpHw6w2DQK13FTejHtyhpX92a5iGa5AiuNQxVSTPnnZ9WyTliVUAK+4JzT7
3byv1xLvP2zagt66JtPXmw1A9BXUvbJd3K0DTkFFtc0ZW2tHje0VspkpaEZfQM5kSoDpKmn+A8P6
Fd/H79YzhsNipzi/Bd2faFCpeNrQ5HlNRz5cxfZXR7LSjvTiRzJOe1L6W2u7dprOtw0CbV/dzzfR
vPvlKgA33ZMQ/wgW1by0t0sdyRsJguYi/up17KhSMeT78bj/KGhb2Vqgh9etl9wpR/olCmyFZSau
4CZbj+hLG4g11P2AkAsJNGpqM/whan+FPV4DPDYEv5HDomYZd98kY4l4nubJhDH7Niv2jkMLIPzX
WhGSUHnT0fUlaDvWbMMKYNVG+gUlnjeSGsmLBkS9PKhNXawNVvZdoVxpBEsyW2DdntI7BrTYi801
DmD9f2wrStomlpjRlO+Up5HA493s8j0J3ACkHslGOTG5bUMh2TigXEBHOK9FzqtejPu1LEMAolCt
IyS1ZTZYWqQS3U5b643YZ0mAbZHrrIEwygIBWdbcgjpAH6xTW2kDtbp8fgE2oFTbIYa2gH6tRiCE
Z7ylzLJi/Ax7LJ/9M6FPPZptTCDvptcPUB4DfUw53ayIQ7WDismk6liaeQzLA4c/ZhHcXBLKryTR
8Zt+wVxcN1Ig8g/9/mNF9OawJib/2K50ARkAG7aUMgOjNCl2LJ/fHxJUKgjIm93Dil5ffCCtNvUO
PV1ZOfz550ZxcfJ/q5DD2ByuGLEHfwf4BzTnkSJz5aFt8V3gSVXHaurIC6k0Vg6KDuMIWe4YodeZ
VIAEcJ/gdEe2to3LQutgvhhne6GBH4aDp13dipbDc61DNoxrBy6sPteyMcrHKhJK+IHJZpKogH8N
hWTV3ipvAtj3nCEh6upzc2PybWoD8v7JUzKg+qOiARo0zTW9/sr7nEApnClZ4PaBqwL0R654/Bdn
KPy+HzeK1LgqZU8GGTnCDizFePY2U7GM7550HfDCNLWKfxuHY8ZDAi8zWFZX2FHVpdkigHcxId5P
yGwShU7YFoc13xQ64FMxm5GEK6r+Is2JyJPwtXFsVu+5MrFB9+MhRxqNU1fdyHRoH433VO0Ga20D
AusXrAYSEuxB4xUzPQmdNA1Q5WDJvWTOiaRasozC2DUTmeFskVnoCqf1jU2uip8OkThkdg16iRbv
GWz/bkZZyvQl78x0BUegJooQ72mv7xTsQeZGFe8KPOK60CHh45D/CzGTsLpi8cuhmBZUg2ayHrfn
2ec/z01Vo1dWUlawUlRGIksd9RsUo9kER42M79O4FDWEUbynm9vUC2vqVNpM1I8ga9Nwp/pXDQMk
olFCLtJpHr4FPP9Ou/0N2WrGFCTac394DU/Jyfjokw47eRO3pdj9dvyYT8GQ0c0oyV4nKGXAOwiO
GpZ1YkyawPXs8zHChOXEWFlgwXIAtKCAUmxYsz+qEPx6C8Y9csvaTxdzXKxW9MP8sb8JPtvuprK2
QPNzAivlmMl/2Iyseh4zQ3/MXilKNnJ/FaMnY+HrTy8bYfjyqRbBFGN0m33YTJnsb8dg1JnqfnVP
l9sE7dYIPgLrKtDp9m70TyFX21MkaXxyGwvLirUiBPnGRSTuP27DzjyM4M5F//RGtFu1csOsr/dn
swCiilLG4vWXwWtUGkkKMChE1sVASAMr0wzxw/TLrhlt42wZdu9l8dr7KDR1wmWqsFfu/W3aVxS0
uR5W70gOuXhpBNqBf6F2tOZDWtgutg3tRz4L44/4mJUuH4qecuCC5M7zByotfRgQO9fSAj11/rMH
RhPLxBDa27ZJqT9p+iMvoybxspduC8+1reTFQQfpk8kflkWy3vhoI2tlhBfB7dk23773a7PbNQsf
2A2/yXR3kPGSAGzFmtFHVfxiBICrrBcne1A2hRD5I2Asogny1wVxW+yn7Ot7+TPArqO9hWfZwwAo
aZX2qHOOW7x3C+zz7cfELu/rzVT8eKEYz9teENy+t0pkGmzhSyFsgqaL9h7qck9ZauZIe1QbSrOK
Q3ZaO0l6DB2bDqQUA865wVM9Fno01cDZ9dBc4ldtDjhLWmFJpEh4pwu1FB192g0SLjgymYDA3pMK
lGvFVR24kVA6j8JwNN1HLGfMEqeS4moy2WNo+eldURjkMb5imR9nPXqGmbG1Gv1NtwyWFtijNMxJ
eTEaUzlwRmuWFqi23I8a1C6naJz2AEyjmV7ESDY75BDTBNGXV8jV3aqfhiyh+uL96Nkf+KGt+H86
YMplGRF8z5nVkv22buMQg13WH96plmePyij5KonTVW8CZL+QHG80byfFqf0mZkB0YYOhcrQ1++2F
n7LP69lGgf8N7emTf+YN54ohqmAzGPgnd1XGLELv9sAcCTjgKPNWC3lrMGgZ0GbNpQkgtHm5VipH
SBzY791kzqGgnn+z6ZEp8CBAcejeT35BpZaRQd2Z9Zos0J6+w7f1lFu1lox6IQ/1iP44H1scauZq
TmC0lcHT67L20gJ5eTnrMzl3wTWFzJFjnPZ3WV2BH5bWAnrpJaITwBGiVAVW2yQN+EZSrrrhQPph
XgSZ9kGcfK+xt+nGbz58I8R9CTHfeWdZuCF1wvSLehMcqVtRQVt2sdTjhi/dy+sP4AnjcehPZejC
oH4UTyAkT+0kTCg+X7ma1l3c8rIt2KNKnxOXh9mJ1G1h31YQ7LXcqMc3CMjZVJZ8lrNl+PaPOEKa
xSiM45UvMKFYpfBqIGL261VobzQKhYICW1LUzrV8tOeCd701cQWMgnazlktbhqh2ppNPPLFtAD6w
KtR0v+lAQRwzJukV9STkNXGW39Y/jZNtrtnGaFr9xOx+q6YTrRShvS/rSxA04YS1UKVddQUztAh5
rT5AWENTgE/Cb+LXUNLGzatujniFrAoDWDsNvGQeIyPe+0EELUMgANY2/yVGGBaf0AUCXM6DLWg5
TCAzfPchmpGaRUUdv1yymHPOzIUYxnEikr4gA88M2TxGmMEHlbPbWPT3eN3JsRWQpheybeKKow0h
pbionQXI0z7mHi6W1zHV4dYx7MwEyP6fRb61VIsEaWdrTk6iBWm66BfgKRwDToNLVTjw7KU9hQvN
3Aoc9Gh16O52Y27vXx344F1Z6DXghY72NemGyKmubQMRx7qq5hW88noohCeMtkAfEZdOnqygsVKm
5x0DOhSCeRn5+57fG8n8mzSCe+ASYLhmiqT5wY6Lm5BwGTxuvFGnPE5zqMqGWqxO/0ft1Mybg8rN
M1hJ9limsSmVrUDYzJ8h0cEkuw018B3DlwaGFmp88Rh3MPlhPbY7SUfaf2CplkTx6GDjZxoOQICb
XK2W7cOUtfvHLgyEzY9TeoXZMHXypOYjT1FcQjymKc9TyDszA5U5fuQQfZWrqkZHY86nXrpq8GLO
4VPFF53asWaDxxlZD04VPUqhgVxyNE03d0ZM9oCLo3avIMjuiycXG/e0SRn7OVONKXOIqKU33xuM
ON9Jnyiobef7iKOha5YEqHY89CkuuMwUjb8jfQDB70+cgEEm8bSypzZGEkzd9CaXgwa8qub0slgv
tIuwYvqGn3uLHJoybs4bhxEBl6MemfxgotUv6HMNkYNWzwUw+IIRSoHv7tMsp/jtRklID1T3B4XI
0W7+AyGR/Cf4JW8uBILyeoUm2xXDc80tefR9tHLcSpSuG8TesXy7+tvsvTsvyf+tlNIxi01hiUck
qCl9a5Z+eOU7K8gozM6mvYzHSIO8ij6aEg/NDhMtMHDRHR/6VFrIYocX9FPOinicCkZYlH5Qg90I
c2Id8mxGL4sXLP/s5QeOs8BVIqFYxUS0+SludsGzGf24KJwQuX4P/fqxYWitk95+w5/sYey/qXj+
Zi0A8g+wxv2L2CWabdky+m+kg8cD3C9JstziXfM6ElWyFo7Nz/PxyWHD6ZKaNjAbVfhbvBnncSrd
rmT6omMuafi5xxPWeyabXbuBon6MgQXcToRujcx8Pjw18egGstvoVfe8I6xHEq+WZOiyUscoMHYy
9F5ysHefhVWwc9ix22YMHyawZ72VBuym2PSIWgcl80aybivr/vIEaKhHhOEQtu7omlDHTzv97/eR
VhKhHwHrzaDY3kixnzSbYnc4XSZ6LCgCMadpbpveqRGaYSL4hT+MA5l30fR66mDxyvixsQFb6048
9OheRsSO/x3YoD/mmPNAygig92NUXAeNba1yiWgkOdtSL6k4QiTP4IZPu9WInkrMekqWXH6NIQyi
/jERzxQYmRFRIplF9Z/LKjapjCdExkxZAY6lcef1LGZKgR5NZa3hQJgb347XGMYNhK+H8W0xaA==
`pragma protect end_protected
