`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12336)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NyunkX2COVNHsTptq9IGD/YE7blreTseiOs
sndrLY0vqRZzpaSCiofeWXfthV0BQw1m3JhQPmCCO3eV1C/GtahvgbJkVIO/WerHlFAxoFlOtinF
o6ugAklaQmiB+gM2md+LEkXEcl5RPShDJvZmaHRI0K042o9qsodlDD+eehunv0nlUTtbHHNn24ac
JlWIERFcSuD8DQV1zBf3ZsQBm+IX1OqSe16KUF+LCw1CXd3aQSws+AGLaxVonq6zqMc4mD15amGy
KpbZd8YN1uCPZ7C5w/8+LpSfJYEJzj9TJfRdJTt3EibgMb8BfULO2k8j7CB6ybqxvs0HPj7CjpDY
KPjRF9DQjYs86EuMKoYVHTG5gWFCeFpKV66piDjP3ZfZqZiMXDVC650mgiUU7tLVcFTcVTzsq0V4
x9smkCGyiaxzGgX1uQfn9VLweAy7AMrhoxiicDmFHryGk7hFIvhtZo53PCitHyjEoEhLIkiUyhqN
dc//ffeVCyRQiXO6HCQfNEsts7WlavNAUotJkqGUVgRqNY+n69MIL/IhIrVz5pfM2vwgRuHW5rjo
u5DN27GdMC4dE/UxoPFDZAvJ+3bE3Cy+PPu2ZiI236Y6wJKVbBl75lH3tKozhiWUAMWFrV7xt1G0
TlX8uJURvdFE6p1onfed+cC8CMAAeXWMXgHshfRHwCfiQeoJz/JbaMwVdYn298EEycJO4t7Nm9vD
DwNQ0K+vtxxjQHTx4BiZh3yzXtOVwD4Hqr2SsB9L0ncIflyIwWTtm/8KxiENvMf73YTxT91K8kOi
vn5h2/9ncRgZVfWJ+VbB8JzStJjGOus5vXWJM6ghVrkL7c7g8O6pGIyd2Z35Ghvi7YuIMXbv9P0j
KnoXOMsW2D3pDjeuYSdREpRRpvIHYB7kclFI3rq+kBmDNrXfWhiTlUTEjjfeJCzv8dErgI6TbWe3
9A7qP3NKn0xQE/Mh7QtpKENm+KU6fxLmS/FyPtkAiQqISZkZ9UsMx63+hKo09x+jkC79OB+W84s4
u8AZyaLxVLZCAlrPqkxCx8XTqDKG2h08crWQxT/SF6nOdRcH314vEc2uxpJkqtSbRTcN8wOiGifJ
vKD764nP5+MgkK7NgsdTykk71ZiyT0HBWICLf26SGHNGKlXEi0Q2HxFMBoMaZIHNc8wXhiXlubgo
tigmGR4iwwCpoCvSGK7C29kb9ftgc3pr2AICK3J0OX/GQv3Ub/yODbrhalE1+7Y0uXF47lzDKIX6
FdgAuxEMPDwFAxc1lIURhS56nMJzC59y7xJ95B0M6ownAwwUB//J43PPRY71rKmeuz57kLrpy5lW
sG+shmXpQ0qe/+ataOJsCXiSzpFQffixjtCTPznZihqELpLqoQ3RY8t+NkvbDamgL5yIYtdACi4P
B4PIlA0/q3BPX87NmsIoUPh4fi1flRH20t2HMZ8CPVnRCquB0R/JUFNDqmzE7Qa9EU1OK0d6eQF6
/aA7MIl5TaHqQ6bA+sprnw8RMu6kMPG9VqZAsfUxhTZlbeA1Xv29vBfMc4O5vH84zsZLSk09kHsw
JZtPWyP9lEeb2zRR0ZYMsTQF7viVT6CZfurkrDxKL0krMahNfv3LZpRihDgsV+HRCG2oQKFxrziH
Tisol1wVDUvsU/bFFLqCYRD+TaM9XbzlpFyBRcr8DzGFd5Q3wufjhw85NlZ+Pk/ZToZClIDukk2I
1B3qYSXryI4B6uOD1cS1VZsSkL5jV88gNMqJoL8WvaIBJqJOSpL3gQZt8WImL/DaW4Aq2wHiiI93
eVfXOZ44gwM0p+p1x9oDs3vHRkvdqwTwqz5oWrg8WdTlk3Gv9TVxOhqybABJ7eqUwe3T9ivNIhyj
zWrTL6xZBUzDhcNSzCWHxTvlUiQa3E47J0udjC8n9Dat65QEyqy4FNqqrblyvF0LMU6QE82YYZAe
MRSg/7zWzs/0Topj/T6iGmUHjRnH3bcIwf3gRbtxCcMAcvks/DS0DyEYN0kpR8Ku1qPjGvhRdlyi
MtOD9Hv3EYR9Bii1w3XBxhEt4kLdc17pnd1OXqGL2bav0IX11iSk7l5Ajj1i4Boz+3CZ/LY4jcZo
D7yAgTAVow5YjBEC77FSXkv4ZDP2V0uicg8PbmjFBjQrNnlTDlPgzeRo9wsoIkftM0Rk2kESKVXG
APtE19gXr+rz8Ewl9hkeaQS3GUGMbTMss4NsyL0DvwHXjT0EJhEGmfzUaarhaRFjAEC/YZ1nhfYQ
TgpYoZdWapomW5L3Xb6TJza169uKfSGZqkin+5BS3xMkqr5h1h4u/1amI3a/8HH6VOOqygW+kQ51
ovyeFmOBturloTZyMaLrUuRqarpO04n7dsXByZ3lvoNaWfVqf5hYQOajuzLoHCz+ghSMvdjWDVu+
NEqawDsyqxN9lrWua/9mEzaElr/yFBNELqYC2pxVBfDO2FC+eTerk4tjUNgH//bBbkB8etUpvpQf
clGseowDL+iY9JMAjMFjnZV8nTHfurkVwQ9oYnXs+cGQunC3MmfD4vlKxJ3hK36YDolAVDO/+vnN
LGJ4CGyyCd77SFSoiycksDIXZ7EiGGtHfdZym3ArmAW9duzGeo83rn5J9monWWmTDkrfqY68qWpW
+ei8TkutexnoPkG4GytMLkgThTnhXSwoPe4LizhWAVPKMhsl3vA6CRfOhE0FG+gKXutF6JRS/zUe
evwr7sj1ngZqqGSlecfgciV31HYScHCJyCTRtsLKrvw8PfKZFiFWis/7uH1cL072lwTZ1TkRXuhk
ANbmMjg9V/G4yriVvm5mwcdW9atAbfEozoe0cxxIG/VDVUurqGiYjzLjee8OOSFVImhWlS+j2dmb
jYQp9VmuC2UqUVPZ9eF+W45d/9h/i9wyxmENl7b+GfaFStx7Gf/zs31UQlfs1WAmvr720Z4k4KwG
MGKb9pz9NUTd82XLvgUZWRSyrMRK5bQVjr5RMjtLooJ1yC2IEWatk9ZFe6TqKpbxYLGmaYYCd3Eg
DoNYRmboQMO1u+E/6pCV1D2uALH9lSzw56/HD0QvQ4wPYvZrCAWQrqwCjgrFKrEQpSOL2UtVFsca
T2HrKzkfr5Jlx3lRU8xo8gmchcGV+EChcg5h9IQvH2vQPab69SRMjI2je7qZS3w/VvMg5DJHHmjv
mLS5KmvzoSeME7TlVxiz0m4TaNYr4d0iTvp8eyvxhpsCToWLxtHMd+D9X+RGZKs/LfV5eOsd3r02
yR27fHGkg+xvAuamcq+Xw40ILlQZBUkpp3tqRx0F9KpaXPT+g/ijobpVP3xUtD1DgmWbMhqsD6tc
zW+837UonGxDzioXLNlIcmzqx97BNxKmJulfSgKy7p2EMwykVXc/eB9RqAg5if7qxVbFCwRjLHSu
TVcFxalkBskYsl29pXOetrHIuiWia2sqlbCoRiH7JcEfn4L2kK9jrynf4BRm3Ai49cfBnRi5lwXn
1h4juOu9kil/hqjbX195YGI2ufP2ZLaLAfrNED0+r3vRrr/QFZ8JI7DKSSAaJKI5hRNtWHr76uFY
g+D1O3htMtuAdAdjRSvNhEldcNVMg/H7PWSP0gOgZpsJi03/L55XmeV3k4rv6rAYM8Bh5SjBQOP7
EPkcIoGFcSnLxYP8Ch/VbX/pCtNrDXakqOK15HXk9k+ZA/CKMjfGccbqjYm+h4wz/xgv1DYsgtSg
AA4MuvgMgFKcwulQ6ZNUTDJjtr+tglRN0HN5jzz+AkJxAMD7ho3e4M6daaAB5rwD+k1kra/qeA77
vf+gr0K6s+8aAyqJsFW92NeHBPWLmihCMWimNxmf6oHVQgoCb6dvFXbBEmNTXAXKiA4bzBMqFYe0
+sRBo4WKpEJRVy7qemT2mIGBe1jpbDrcagKB/dsrYkdLntEZ6C40TCegTJRsBSSlQVmEFrSspJyq
T2Pty5X1NFiso1cTZDPn8N2f7CE9iuiG4WbO1YZXkXuRYoj9EV95l43MA6Eh6hUFRn/NUlJKMFhT
lpIna2cSx31hOZO6eVOyv+gpD7kRKxFD294i+xJkvtBehTfmYGz+nQGW9/BWNenHCaXbEU8Ly2Q2
kdxeFvdzSqrogsAczNqKP7N2Hf/Uipj52Wl1ZHr5V1pJeDdK0sVdx8S6uXQNZA7oB5uvTjtDAOV0
qDW4ZRcj7e9h5F7NRARXgZV3K3Ivk5YFpBlnAZO1K2OFVtLz4VOFyOpew+/CqBcrfn34ZGCUWwWI
UICMGLs09Y0eRWuEWXkImgIbnszQ3MXOngLyxjXP3BT8El2Re/4hvMN0d/8wgq0UV/Ws2t4QNqEX
E6TXCYO7iIZcrnHjy+ynvap/AUw8M7eSy94E7Zs4CrQ2SVqDYGjiLC1OWsSJSfajn03UcAibTUa/
yLUFmZElzzYEjfcf+rmJOwGWbSyNnmONVkV0amlKsq+UCWMkacZdF1Vw64Jq+843P8U1fK7djJp6
PKq3QKFJBXPv127+PzENPZicjWAzjs4gjeljMJHxjE48122JSrgWsU2mdlsbBk/jjQO6cWPXmMxl
0PpKOnw3tVUJFwyg09gqgynXWM9okFbBEFGwQ/n2MOYqowwIv3F8RJR+CP/rxcSh04K9E5Trclzs
NOc4IlUDkSMbOHq9QNQ1NaGOIlCyS3k4Ctsv073513ktprk5Rkmwx7MHFkN7urUxiFlkxw16+CXS
PzjNDOzmQrebmKHBjl6pr7d+83aJ+WjDQdiOxOXD4yQGwbYo8b6iKfZJc9Mh958+/nKQuTjvXHvV
66wctkJxiwvzgqnmFk++hGePfprGKbArjQJ7a5Y+mXwtMiSTofYEznNYy04JUcwO3mC2sZzxldSW
ByvMqOtbioZb3B0P8n/llel8Ax4ZOU1bk8voFTVng0yzHmsW3aS5EotElFdxC3RelbGXa0jS/3hX
PjYSdtyClcbn+DcJc4DhRizcoVqzQuGv2o3i09tU65LpI/nSVPyI0+ol2v0zXAtKnZ8lzN4jMOh/
Rx3T0h253zcOl2ydMEfZ38Qdq4b8xWG3IzNcWsIGTNK4kkFoLnx0PODBLZ7rgm9SxwyrxyALr/oY
SfskNJ7ySYhXOdU4TZT1K8UXjA3pYRy1O8rtRFLWzoUMwosdnxWe5k7CJuNYWt/JDPoklqCQFKVC
1hE5/Em+0JM8AWIHUULceLjrKawqoKFTD2ehmY1jTPSAgsujD9KMYJE0yGJhmucWcmH//6Lxe3eJ
R61JeNj1pYaBhZFAk5lTvIwPyTxvOMdrv/xwXt7m4EzsFFU4Uq7bgkvqeK63XMP9PDdSicaa6PGB
gBIxpTAThACredpPGNNAJVZx9XCq33yHih08kgJOP0BIH0pbLJq0DEV4U+0l9ugc0QBXuN6HdJBi
FH3qjGryTfrAKNGPePoSkp5pmFIEnL4jDFcEl/fW3CggRkthZuWSAKQJD3/8lQYQT5v+Usg8yxKB
E1S/ZHFLLcgMcbPDqDtwHWqaQFmQRDIUpEbqeyVjzxBr8XlXkxdTDu2nK7tFCWNZBRgtnL1ccyYT
KW/KCKiefWWpIiU8kJq4wHgm0dxxh4K57H0U9HNX7x27fAleZufYAoMr0VAcBVtSKzhKjmRljEPg
ibaa+F1U2xF3Eyq4a1tDRTAt/xsSrSCJ8VSoQR4AfmSKd98IehSiqmKIUytI+9T3er4YQ0q0wZzn
50ppwMW32/juq1URpEXZtbZsviNQ8KWBXifL8lCA3maBre5Rzx09T3v4zisN6peOK2o6SiCUJIcE
0uH3VPKf863ubb5Xe7ShW8RAiMNcl/fJXogojj4PUvtL4wvEDuxdyFAbEJ6HnmPX7I0tZZVfsDL0
ONrHpTQsQFhy8VksgDAZ3QZxf3af9YGvBbAn1+GnRUxnrO0LYFtNT9Wzp2xqVml/yuOMmbbW2t03
ZMw8AOm8ZGshjDiqP0+R1CTBXf/IuJYCGGaslacqh9bdpw34vSFYlpnk4HXAenosl/wtW7rx0eAg
P4HMtcHwRNY4WOYJgRoEg9tfYFmh+PH3c5pWI5ECiGA5E8AwdSVIE4PkHCD2mAy18PasEnlrDLLF
ZM7AcgBxnXAjl5Kk/QxYwhor9InHmXPg8s4Ey43kQ0V5vhHB80TOvGxmhAi6BKeSyvRTUTDRXFwZ
Y6eMBdH5ccVz+z/dVcV2MtE/dWtEeK1fczKosLCmTrU+fB22RCNILnWp7NFCjV1417tnVWFPdhc8
9kAhwA7xReteh2YS94auLr+XobYfAIl1GkAB+q/ygk8HAk6gMnSzF3ukMsZ/5jvxDh498vlvJ0DD
LOuTveMTOOQ8gbbeZkdNn0G8g+sZUIY39bqoQi4hAP+koHvHw80Elcu5F+V5lZeQ/R5YUnL6PcYd
eSS49OJ/zRVGcv01m60J/Z12f82v8LVwPP93JKjrmmZvGeTaM+mc1FcZ4xPehbJHa7DIVf7N0PHr
f0BPckHkTjdIo1tVGsYM1qw5mVb8lznqLcdQxJmaUp9guhIIqkK8tHQpUduMvCslneN892gcyhuC
SdT3eJpLhOg5aNGfLiyPeH7jkI/bZ0HnuCZmYBmABciAKnMLFjY8GUCNKVUqbCNCsdvcq2q9vjCq
0R5CUQp0xO8YAEBgeOa8IWvlMOXKBs6QpeS6hiRsPa8mjRWyFE8RaJWBsbNonRTD7orjSClKy0Li
kE3dlUBbYGdCavhJr0qV1UmuPeqI4vVFjII6jChRCcbZTEGPYz0J/aP3aNyJsAjc/VygHYajzj/1
ifO3L0C3Zs9M/g0ZYnyDtuw03EcQ4kgTMcnvZdiFtM7jspIQcnb9lAcObtHda6F5iFLe5pxWpZHZ
vs46OxdjBxwOtrTtwfCJHInqBeSnMZsO05MKxEYk8MftIDpr79EF0aMTwHEiKVZDkm8ZKi94zETE
s9ClLRyCci5Y9olntqxnYKDL0EdENseB91glS1gdsIKtgRy/7GtYrRVadyI8AvLCe/3803Xcb0yG
BLin563cG616f6yGEFAxiGbsSRHX01ghSlsYchBqCNyVeD/AQz7jqJwnFGJ9LvjFsPjpPs+2q6N7
Ho7cGGeThBbFG2KTh1S8P6S9/UZQTQzTBZxNq3RGMnhwdGFkBb7LGFsmRT4VAeNEeYoL1n/gly1S
RmSB5zxkavm2cDQgIHRl+3G6KpHpDHlg7sNva15p2BEDemmDtZnczl+CU3vrf3qCFEUOCtq1+85N
hzjgqIim30PeB+tyYdCDPrbRBBqqplllTNTbVEz9EGxoEijUIf9OgO00nCK37sbMe1zecj/SvZoI
YLPMAPeT5HsnTICrPChumEaaxzc3Yr7uSwvqTWoiYjZl50gQZOpqx932N3KNxrru8yNcIWiUatll
f3GQ9H6oa0T1likequOn+2Z3zeu9lDpOM7PNQHT5Mw9zR0vRiCu56UAylceTxQn+5Y1xS2GuFTOf
ItFerTzeDynsTs+V1w8bnbVylmRPbhCfZL7UV63ybipV7LNv6O7VTm5BPvWpkYj97pLyNk0cH2j0
AO4mIXr7AXynI32wOAB9vvYnFuodepHP9dGMm/MhQsffFVtn9dvVMJTqnPhFqk/ao8SPRkicon6G
0a1eOeHMTfafEqtJRej0PgzJekl7l6u4uN0tvyJXRTWMj6aBvlo2VnyT5gl//Ca6WWGosR7mw7xP
GLpSgeKL/J0gSUQ1undcD+aFvfoSgpLZEs5PA4p1h1D03dEYK1h2/r4mZXotBttz1GeV7HqTwIt9
MCYnm2hgKnqmA/WByJy98W7UFRlF5PRJqp7+6qpHwoU3dr+pDHjKeMgubhrfGCpo202ORRguLNAY
hkcHOCW7XCMMitnqK8T+pVpyj7pkMBxLUGVnmyzDwXsUsKR6kV8YAIlpv01RZnlg9xW+wEexrezU
PfP0WaHTaVuAHzByIfFwwVvu4/dFlmT/bG4GktoxcLc/4K/KP7uNfWoSeBjSHD1kZLKVRbIdJKE/
6q7bWTFTxfPB6+gStAveQXJyuNmE3F8VKLYOLUvmfKw2Q2wQd/c2Go+QwWR+vbrZMfvkczwB/YOw
3O6oUWVoR/Qj6tdhyofZMso621baUlUfiyrrc1Cp/+OkSc3xLaiDsQUsEkCE5aMPdRtF4oM4Ge8q
A5t/civFv/9SYvuyINenmUmstripspYGC5gS+/je/ggtAv8EGVB8otUhEUT7HFG25LJyVCa/bMff
1ArbPRA6WQrjwAt0defmbO/PQCT3RVfknjWL2vwRJkno23vsaKhKhmKOD0LFQFhVNK+catDDtxkh
TucuGkz0rPdUUAHvJcltN+xG5ayfVs08LcoSi9pNLtByMqWSsY62I9kRKeP3dzzY7ZfgqDTMNPVK
WmoMzsl8BUOf44icrQ/6xH9fNNrB4IGy6gKozi30waBmV/IlPDsGGrLcEbCReOUfJ5fLQ3Uo9p5Q
/duGCkhBuoDMsaicuSc7xQGXh4GTzjTUXZzcrE0cjxws2QCpZTYxLKFqAIWAUGIWRM3FuIJPZ2Ys
kiaoLCPeHeC9KVWB3nPbrA05UhqrtojSmoZ0/I5hDPOLEDKOaL/e716V092SMVGRde3lua+S7se5
HboNaLAJq01Iugb3fn/LhjIdPOrGMIa+VluGFOYB2pls6zAd1nk2VQ43hCM2lOgEVbiAzbi1UmO0
gSqSg3OxVMX98eVqKpuG0nMa0w786PVi2dS+xONV+NBvf++T4KD6vl6wpCXTBbLKU8rToBbxj9ka
3wRJ+cbafjjKNIVwkOpwqYD5PpylQ5y71T/pE3r2ynboD8ga2ymreyHMDBzJNOtZLd/0jUK2C2g6
OlmtkNn1KNoE4FLgGYWm0kkNfkiJ4Q+SleAjnXF7E8E3RccwrHnOnWH699TCW9cjRwBzlEnyw6Sj
0g2eWDJL/BqpOitfG3R/Y7Az+iNBH/kJ9Ogcp8ohEmFbIpGxRblMjvpsfTX04++sdm0YlaFNGkX9
S+aqb+ii4UT4QMaNzD4a2a5wXH7PmMiuewbm5AMi+VVdFElNHU47lfIuPyRjyzmu1lYmv/lpuWMA
LimmKK2wR/FZpSO8KpgWujSL8WUfchWvTHZoqwcb050fF1ktPb3/UULR3wBVjOuOyr6vSCUH6R73
HlCPIL9LXhRj/nCSkev2/z5pCta7i9GygXRo4BQMhgXiffsKesC+dDcGJXsTs+jK38KN/2dTodXv
ApFVRa/dTndzg9DGpySNplH+YuH62rCOkh7oGbpxFNJoBxP6CC51B3NbVtBAaLm2pz6BftbhW74Z
QhXcqUqZlNLlXGhx7WZgMWhl2bFt611aA/0YtZAUzrIOAkVN55DXlYmVeEjnM1RFPn8gO8oryoIu
QlRRNJiWbg08DPY+duxDqBWo4mQAcz9/rxv3BgMFpkNDE+JsAgL0mIY/8vGPcoOjKWiD4yDdv2n7
bjE98Jv9r+ZhehEpeSWmQ4QFzlvh8THUCZ3aAshGwOMxIeXwrdhuZNgtitXMiXaanzSMKDIFFvfL
72TsKOzXqAad4zyD851+Uz3e3cZCV/K0u8ItVQvpwW9ubO8g22n42/mqNWfEKQ49Cf1Th17dF3pe
i2KYu1x54kTE7nO9oC59Kfkm4CKDYoYWuxeM/AiCBXL8AqrVXTo9zk1b3Kbtm506FfWG4D4ypiMf
AxunKmmmHJQ4er0pOp1d2S63crFPswa3A327jsrZNFGNcY+srPQgdZqnHWq3C+2kgDt+8ku+pR0T
8BuJe8WVTQjC15IQDIre3uwfcL+OF16lMLVAXMC9rysq+SZ9D8ZufB/Fjjb6qTYvr+IwukOUDRcs
cQ2qTtwE86zBViNigHbCtIc0Szm5GIYWOeOPz44zQ65Uq6C4gU5AyZJH9ikNjHkk9dcxHA3QhZmE
znX/V9xaqO9DU83oQhB8t3+l2WfyZvxN7MEXJIfgd8MMzuVr5wTrl6E/iL2LunpdjLSBvZM3F5CK
pADiXeZmHJucR3vAUcHzORwMrnGjo3CYYZwG2WcVKHXEWzj2j8DVofid0DeCfI1eB4RyRUylC/x3
VR+dhDBBy1aNDC/m+9GYIXnykpA9MLmB7gG97adAtfW2l9ZWliTHINvT8o9yHXpDvFESCVPIZL/K
JFd2+nkLzUC2MVovh63hRU9PTMay9aK7bnx7puxxpHieuG6XzIJe8TxllHt7aulDIYshMldln4oG
ahfuCvZ7VqaIjVUBUv+MXmo0BpeSjsyfLPtSfp51iGUFgSort8SH5O8sZISEH1QH7ZwNSZRocqpU
c1GS5IuJczt14bd7+46XrNV8oHFOI9eUHIciMTVrHZVZ1C+q9bbaGT+qg28xHJgEHgATHa6fTu7z
m7lUrw6rW14+JPAM4AoWLeJcrcW4K9bsl7jW49pHd5hdqahnmeCF1i92kydwarph7bc0//BYJ3+d
7R07ONpibkxAoLV8NRhSy5NFhRJVwy4FgDxVrcgsw0h/zKr8jCAIaHwmBU+R4DYeWwwMYW4Nvwl3
Oc/xbk05+gkW+p0eI+QVDe2hf7oSjBL9ouGTUBagweJVeICH/LgIXxHLWrzEn8fHYGHH3DkPOYOU
36p73lJzSG+QHLTsJHvUz2pSSaIR4YyoIR0KtPdEDZbgaE0BSN66V00F65Rrha7zUt96cwceD6rU
JVPKVdZ8wiVixGNRBDDcumSd/AgZpl4ZZT0vrp4RexRrMCfDfLVzpdBWsNG+is6ps64b8kSpqblC
AB6EXmR+CS4CIBe4fDlltPFFCkbxhXKUULHWHJ8rW2iftKWxL++p5vyEjop5VpcpkRJTP8DrGhPw
iyHM7Or5G7Jfs7DAi2Mitq0opjmfZMJkUm9M3wLgQ5hDBLIb3onj3XCn+WBTHPI3PnIVFDzfiP7t
2/RshuneI+Y5fH17K8/u55XPJEzHMePv9PckG2Sj6NMLzKQR5wb7p9tXDuQLP8W0fgW+IPFEV/Bw
ObkBurDRAFVE5eRXWANM5wjckxs1UaF3OwUpt4hWOwuDM70YuL72nueqnydlJVd+P+cbYV+o9z8n
cEFQ1BnI+wLfarqRN6cfV02YRlAI5l+8Co88xSNDfMi4QlM8GzSieKo7mtr8KKextFeQHytnKecO
VieMvtv/hTJBsAtY9uSAiFcdsSNoNdkgxwTHa4TgldyqDfTSWa1MW3yUsV6lMZAi7e1xpzl/rd1o
CxABSb+9ZmXNZy2AafOXJ71ADvo5ZM1QBnC74zBcSffMeq34kFjh2ktjtd87VsHHCbysaQEaM5KT
mzX8PXNtmeexs3dEkCPb2j4C0Dr0+d5qUEgaGSfRXx7KlPcf1v6Q4E/94RMTibnT41DtqFtYY+n4
qfSCFnlpeaynr9ulTzhd6n819BvIfaIAResLExqqLRadaJ2jFZVaawWEF0r4Baqkgs9lRnhRQD7Q
+7OY/3MSjWzztDCzzT1tX4Eyo+d5KfJZN1r9NuWGBxDiHp6JLi/5pSy2EcRP+cg9F8uNiWJJKS24
F/whY6kdxMg0BwqZEMFWGI14beI9TAo64miZ3ogGhhsW94lCMUSCpT3hTbXvCcQF89exJQRxN269
X/vIJz8D2QPnjFDtr3f5dyolJowcgvnDonkwUxravfVqbRe+m03KLr2im9viO2uSKiwYYiMQQNha
eswSXnq0vFDC5g/C09nubzIvbvw5UI5xWWuFehZFiHPckrzc/2XZhdv5DIUle6XhDrFz6VHPSpbQ
Mn5jHZKh6srsRbJhIIMTzqpFdPYb8BQghEIxFblarVJeSr5bBaORP6TKLj+NEGllNvBDsfbqw4Sn
vG0vsibtXNmrDbqsKfFMlx2l9dDSUC/3Fc2VCzR7YUblPLdNEGrXUg825ubFrKvKLiuBZdu7KYFZ
fyFkAKWBIB/mH2f/7er9BU4uRYXu5tFt3e0jtYUvWJmjXs5Apom4gw8FsI1PTZiZsgj8lo3Cbm9p
9FxvIssAaESbXCz1LaG4gcdM7Bv7vM6uFViwppsQK8Q/zZAvCFb/vjNVacBAr5dEHNhhHXAlTmj6
XIgGvI7L55n+7O4cy1AvP5pk8AgBmjDQGS4dmJ9BUQQaWlQy8GtqXPB0qfpEVI5lZaTwKvnVe7b5
80Q0jUcBgt+Esywq+i9Oq82wkrEdOOCN0Yt1UAEQeGhZ2UwE8QkcU4kirLlaxRpFO+aPl1Ocxnk3
OxmsQrkquy9ishQskPZsEybGhT56upvQvhWFWTL34r/2jxhpeY3yc+3EhaKglSWiCrx0OxCEE7S/
vtKvd8HxcXxV8xP26LQ0MkKI2izCLOBor5TqTCZzQX38EjChR2xEAkKBYVIX5h55aEocg6AKYAf2
UXqnTlQ0WkglnQkxBTNfoWW3pVOSUHhOCXIkSo9KcWB0z503wOPpbGY4ji2iwzbCCuesdW5KlOSj
37i43rNZJUuseggvlrALUmph9j6t/8CtVUjX52mjnGmzT/38tRT41kbran6m41JPxWhNJvCGr8+I
HZ1O4oazWg9vIu1PKFQFdysu6GnsHH//JLKUMVGG8T6iLXSZdY4kG6Is4wL5xQoXTtlVBias69Q9
xvMrwvN1HDmmo/Nouq5Imfs0vIK5Z4jNScs2wKA9jFvt0QztxXaFycRMJxD+tiJLm5MOH2Iwy6O2
4mchJjkHUs07J2bKW1UQzYAtJldsU9K3ImX707WP35s4x9y0bAH+7ipljuuletvXh7HTjG6vYP2T
6HuKYs3wPjYbtJPyiuwC9JF1eljl/hN4wqVru9mz6kl1pg7yJt8rHypwDgtA3GJsnTDJAR7mIDbT
gVtfCn0RYG6rL6fd6c25WeGWtSa+rDWXlL9Mfiuy6HyvQXHOucRKQ83HGE5BF/oKVoCMlGMv6uDl
EXrPSbUj87BOt8qxXXn4K9SdHTxMLZ1p+UpVdSGK0MfpbVZC9vZm9NRj8tbFyWTZfs4bxZ3LNSaC
fZEBZ5Wn4MWVW/q+uKERJjQmU0zUlRG7g80Z+/1w/Praaec8lAViD45eUWVW3x2qgyJN+P/2ULFo
+r15dlZ3axmhSKixKCW0jRox1FcQ3hllOhs4cJA3wT6qkD+gLesv97kDC8YKu0bXGkDw49JZHWjX
WTFJSQ/8+/OOCuMPrYC+w5RqR3+ra53TRWp1o6cWLenBXF5GpnZ1CGquAZTOYN+CP4bAXhYF5Dq7
LHJM6bAeq97t7+XPuJeIEEZZia4cX9/3ziZORZY6hU2IiSKEGOQN4LXbq2TlTPPPueQzAUzygPrD
qbtMORhVODm5erqlRgDo6aqwPBImnPohFex3b1zMiF0niZi2c0YEXRgOBR0YieENoH3DkLzH0BQ7
Obx2xlQynBWohvlvRpZct+HRJyXMt2AnoC5nixIXDkO7BxgZmXA7q0BSG5U8FgZzf5aKISRazLzA
yfyTHpmwdP8hbQg33SouUIIq0tipumdR7hgaVFJc6P6gsjLp1fW7UZIU90+2mR471XVL0kGHhWZJ
wGdx1XIumnpPxIBmPfwqdDEPFZi63EbvHjpbn8JW/Duz3yppowc9Zfc3XWyycdZ8WbzFErdZJx8b
FsFQ2Ivf+rzPOxvL+7Rr/qgZLpDlObzUw8voEGRjZ9dPF9gp7BWpamowUv9CqtYA2iJsszSuapb+
1p7zYw7lJCDfhRipU7fRsK88tD0Fjrtj+T1g5S0n2mHNa3YPzfJ5seZ0Hb2t6AoBDmRYioSH16a1
IZW0JHpstpI4M6b9T5htBwz6amJUm2CAl5FgjWZ43qnr7uTBVOczj8LSNeB/t+fALHGjgZ0yi9Q/
W/Ej+hWrLF/IMaAoNbCOz1CTNaTEEhTZ6Vxh8TVmNiwPhNdSZU9JOTSvCsZSRkJ+mp4Y2qrhPGbT
fHHW5yHtkh3aexVigArEFmDWrwVljMcXTpIS3O1tVyUeAUQJd6AWREejmRyXMnN22EA8vpAp1WN5
SJObIkNYC/85s5kf3UopxD0b80IYFaL5IK8FPd1Ga17OrPYF9NRZ6mnTfI4Zdkp6T9rvUsv9rE6a
OfE1K8I+cwjla2Bh2g+4c26MDf+4gkcb++PJOTWQ2cV+n7PuAlCsYF/TDaiqEDx6uQ5+20DLtWnf
z9pIdDAMnoJXUYJfXE+Wuvu4mrQAphCe//QUz8KqBgRI0e4N/DumzCxx3RrPB1Om5GSu0vgqCx1G
SoXDkqYuSY6MGg8FOQ640vDlbAX9WHHbUkjtp+8DCSXeBNN/PE9fyLzSchnzhyX6dRifXK86XgMF
iOv5G5RWC7RhoX7vx1sA8dLGa5god+50ht1/KvBqA/OxemcRADoBpzlhXa5KBOMx8JCZlRebPSVV
e9Vm9oW4TpklPmHjIiGzFA2igygej3tAlYJd6037v9gO20W4PTG270BX9IcBFHUASvGo4u/WTOhz
usjy/KYrTPqV01aJvAKx4/Zu6N8flxsrYZM0IJXBzlQWCVEDR/i8qkQw7maAS7/5vEuqPYX5JJR6
MI3gyS4FU1tijKMnaGuqzD3S5NmZtSWdTzi7gUTXwncLXkSBceava/yuK7byqB5EYgXhPC8NhGgy
hz2tNRuRVGFl1aChf2NKFYMDYU+2zTRbhjzV3Wqpv8ry8hqSxtqaUoRoI6as7jzAVSiI5N8D9Urh
Lo7Yq45jjO0TVKFoV6LQ18Go+5myUY5awGCTOvUAPwMNPdcA9BJQOWWlkOOViULYgEKhjd+7vF5L
4fOuis54Z/Ajz7iyJISxPYvoXnNzALKZ/04T4yEAJ2dKMunxATAE/+ywqW4LHOdBPo1gGSo/lZqa
Y4RNcBOz+fKmpd6dHpe1ubf5BWpfwizwH0e09Sj/iZ+F3Lqbg/pqUTiPT+BEoYnImIEdDo8fspJD
OlFycoLduj4J5/tHdHFwVo2h/59KXwyDvIAqswnXwrXFjL0G0OMHeIvGapq47ttUdMTC2kwkM2eY
1pGhnZB3D9+DFS8hCbIXCW1qVFt2UaYgdy8UCx2KhPlW4FHtrwQswZB0Xp9P9TBsOlHFWlG5GkL0
uM4UY6oHLHIBrmKwHdbqSIGskQ9m+XRoGXCABJRC8wo37+sbfu0VbQEA+XWjAsZZCw7GOmBhjwVJ
scbRePNg6wsuTquPaf9FdbxC1aOss/aoUH3PaGrlBu9XhhJ0f1fimW8Cjxwkk+OAM94KBLFbSdDl
n0G/UbESR7UbtQgEDNnah1kcoRI5SAJRqAJamW0kV1kBkD83dsHVqlNn2kpmwTEjDuW+Y8L8uP82
xVava/FE4iY2rCKhnuTCngLAbiFWK2iKjKN81RVglqqKphgfVCks0ICyd4gm2XLr3mGD+8s+LQIT
Rpj0FQY9jKNCDvY8FPX8AZFPG2UDNC7+NalhPMGcQlmJ5rcvSRAWf0DTytQDRw3cKhhyiqNH1I23
EpK5/HcRa/NGst5Q+5y/DAL+j5StNTJwHqSftLC+POJR3GKz/aWzbaz148ieqzIdj9vVfaDzsVwp
mpUZlUTTUqt+VbJlEFc0eJN5ahFzf1Md9zTamyRV8mBSAxEH8XLfmcuJRE7ofI2lOWH7QylaySOL
qdO07bGA7adgi0ih43NFpLtcByM2VKrwicdK9/gnOEoQxf3cNPg/yhWYZbNG6ktRJkpOVjxPn9mp
enclCLIvLLQPyx0Sjny8arCMJsXCjx2k9dJhioF6CmH6jTWQ4L7kawDZS3xDxRPUuq/s0MJ10AF7
HPkkSJzfCjAI+qJ6/wgRN9R9mS2U7qPI5gRUb5HKgM9QTSxUgetyq+vpN9dM57V/Jv9wGpEpnoWG
v44VLpYi6xuwcfcYKWiBOMHAGZJAM7ok6QRDhkP+32chRN07lOcy1I/6XUrG5sHINpP5b9EFwlWV
dcWsMDp1J/GLIyP+nsajTj8zDy6tkJNOBu3eoSGxhERiC8gO4zGAnEC+526zjTNX/HZ2xrFmKhEY
GoyZxakJYfgeQRh20ATIIbY/WWSF7NlmCYYRWOPolWnRa3kVlXjSGmsYqWoGUnrtAK7v751pENKm
s35W2nvH72MIdLPZwQ/klmoTx5KihwbswV8ngA/uYtNKo6D/mDOQd857fqgsJXd0grZBUqAFW0r8
vZSVpUxoVSb7dqIZL9vQ+q6sR7B4oWzHNwJmaaBhbJnvWDy3Q5wRqHxXnmANL3VqmfCGrTkI/mRs
KuxmkxCajYsPYt6Jt7LP1Yg1Z7/FQUA5Xt95mwsqqUYSE/40+gGgyGo8y3pifvH1P7FRzxW08sVh
3tWoQECR3/gSNH/XKrZ7NbFx9qqs9612VBpI3r27AIZ9VdtXgT7uXyL4qzX5LQQQ/k6dfQhBdtVM
kT+pmp3CIe+JbyrMzn7vOQ9nYkcH7DIvq84EvQG2pbKMDJD9zHIiNsOjTZcnYPNdGZKkyJ6LsHlP
MfwF5gg1/BEqmHrUxOUZO45Sc8kjBuNU9LrWsYhtQt097TDUdpEKJ0fcoa1uD7iQQWAfg7zicLv3
VD1lGCvhqLVDpEfZsRN9K9DtPhsmwX++
`pragma protect end_protected
