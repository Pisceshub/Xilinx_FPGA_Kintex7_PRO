`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
BCC9rc/UvLO+60OKG37h+5K6XVw9+xBlmGSPNNtCyHiGBNAs7uE+P7kAaWn27GhAeEpR/kFMWCax
az/GVqBT8w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KqqDQUWeBjbeC5Do4n6RoTO+nx+zDp05oc3Bq7j9aHdTCyJc3x0fyRiN85/GGjrUv39QuhEX8Yfc
PQieFCLLhIDiLcaO3g03QeMtoC4gucQf/+wx8FMN+etUNIAKvGSpHcDF3sE+QU2wR0z9UkcquWwd
T7s+2xbq6nw9IgjIn20=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ArQFRYMFjfIqnM01+3BErkf89TR7vHqh8+aVuOpf4ehtdLgHJ/5eVLEiyKB8J8p19WP3coK1LCXX
zKhiKuxxeGtbGwfm+yWYlBx9ENRZgRCMJMCvUsDVN2so7XdAPwkjqSnh0W76/Lhaf+d+pvRWlgkW
9DQk2DdXzM4eoYWj8692SXfxs2GVr/LFsjE70VNgWii3g4b6hbt8arRzcBGb7WdSP01/Vrfupwes
wvc5UsRUnFw41z3BPXfnJG4S7TLMUaKkpXt4XkwlgjRwtf/TFvPay2nUHGQKbMhpn3k11OWjCVq/
je5H9c1eGYvQsLZXkrE0A7BXPj2zxOkaxG0eew==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D+ZRBE6u1yF80QejORI2YlK5RectTc5Hc3ZGgcNzOnHuwsKdRLXxgO2EwzuQORFrUAcI2O1GShfJ
cDaxaqcC2RUD7RA3O2LsbI/gqaNLWKfE2cPM5kyY4LL3UpWPM0Uo5ak/GypCYQ+UOf0Kv83mOrCw
gTGIytvAqr7oSLY9s9w5ayy04DJKSe0dAiinfq3BJ0yg/LnSWrLQBOBrA4Wdb3lM1weRawy6ucLs
RISAq5pL8KX5nYwI6yisEb3R/a68Gt9JyNzCGetfTfKa/ZmZFgr4Mj4aSY4hNGRM3OGia7fX8MI2
J9WLaNV+MP1mjqAewxP7QuQOtPQpJ7jXaieBRg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ntat/Y12i+xTz2OshnCjcnc8y9zrqQygo70X+7SJQZtc4rY0Zflni9gN8Z4mJ875xuUjX+lsIH9Q
3xBNfK+u4PKka3FGIKhp3P9okYAJ4aQHDoQHPys7ay3p9o+QjpDu+LoKsYOvKcQvSTT5h4JB/ADm
8cRL+CJAT0lnMoC1oD+FzJaGD6rbUe/m+ozDAZO3EXBxQhmIERbrgUps+YqPcCfIPBOirPKyo36x
gPacfOHCAyEnDGqsYlZ8/OKD+fUUWGYGW1h+tcsLksdUksFOzpwjaG/aylVqeGnpGGdju9YCZsxR
FTDPxHHSYbWz1IdEVen5mJ4AEFHyNM1FWcDu+w==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iooVi2sFmNJOwue8KHSUPRW3tf4tB3uu74gs8Z6LDvu2knYgcu9jq++JPYpGEqao7R4n5XlVPf2c
k4alUHvp6Q50up5xf2+TM6YAlKOh56q9Kx06TJnkavZHpzcVUxjTO8lhG7ZWXd4Gx6jTrcXay9Lh
hZnVvqIrYIf7F2M9BVU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TKJ0HbePLQGnDE6xQ2nS66ju3E7NpHUMIS0eN5TmIrTiavo1ur6LEw91l2unykROGHhJ6ADO8P3+
+vp5WK18tY3bqWh/q6bhiVRnEA2oMtztFhG2JpSy3iPMMzKWi7QDcZAMQdJjnf/G2+bGK0FCj+pn
IcyQWYXOLQCp2MP5UnYVxp/1/Rseo1YZ2mplACxSxS0C9v44JZ0uWfMD6EGmpBALrJusrcpykUXD
E/ZZoTwRUL3BWG4AsvhqsJUYITtSPAjRUg6DenJjWOgD37PK6P1nngWyf9Jjbs53XYO39akVpu/l
Uewa4cLxL6R5/kYVDFXX0OuYcl7BxOYxaBLIeQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2976)
`pragma protect data_block
eAOL/opCDzBH1z0QvPCIvObuiNpobtG5rcN34aR+DO/8ElPVY3cRSK52vKD0YkvUlwDW9pBK4nvF
176bUQ2NUvNhuZsbZ3ma/PagFYpRY+tJhPpr+NOx+Z3albQYobwzzimEX9n3oSQg17l1+RF2QSWe
KpCIYnr+F9e09/5n7vDnNdNi2lbmfyEmf12ejIuyAgwOW8/ciNo7ApUgP4n/rKDzcPO8jG31mDhK
Ylo4cNAzZ4XpTLDJ2mYrFj1n5s/ayiqecCDPQ8fL9cror3qyk7uzvszvTW5mCEDh8Li99G/OZxdc
H2UIGqMnSye40bWy71RZf5M5D7+IuAZgke0wc3kOuj6Iip9wQni6dNpAZdpb7zpP3q1D8h+JGUgF
PU3GpUCpSRz8ZFFUSN2TyqZV1+4wVAelzu08lnQymNzIJ3y6TW4/SvJ6KWfTiOp4a2/LtsQgVNJm
xKK1dpnqDPbfUPPhil32vBWc1lX7hkCuRcqCujL0dr5aeGjVYgzY8+Mgk1gmEmJ7oOWBUqLbeY8s
AldPrlN74FppfbpK72l5UC4n/k19L76Rl8zlTx29AEsq9bgEXwcSvr6ePSG0wIeCkWs5f55p2s49
chyG3m1IE458/s7+C6D56muwfQuO/W8lBN7LYPOyIOhj4RpxiBq2WIyNAheiOmIqYwuk/Xt7SjtN
TQJr/82HfThPAxCrflOCLbKFTDOEUaHpKHFoFYG4IFVs3QIZksSeZVHzlgaFDmU+pgmH8a55rjwG
i/FW19ISqD9H1nwNW/+350l5owyHpfrvckTmcB5OS0TusYQWTcAXxdABJznjANGlrCjVJVlA5bsV
P9g+xuUBMBUkSCOi8YDQJkOr4sobp8aIrZ1H0CfeAlqj8YE26w5UK5GbzJj9fzzuMlk5K7ttSTs7
TEwHjzHb5uzbw1CUWocUz4VwVhwOZBEVFw6STA38pEiaFdjrYFDQ1+4rh/SwxWerBno6E3/4Huhv
4hY3hitaekV+wVcv38ICSQk1Z//Qc6qqwmlljPWYkZXIc5zC/RGbAakblMtCq8+qUKnCP7wYTV3u
nMFx1mlSJ99RZDcoNd4T2vOOvB66yBOennkob9qYTGVQFLli5k1k+/sD7YMLL1MdBbeWTfWP/Bsb
HVDoRbEnYLbxobWikeVPTHoyrnx6DCFxYBypEBnJ06cxm0h4kg34QdbqWnQsXZah6spipLP1YyrR
s+astWhh2iZH36s0WTbH8FOlzWhNhik/qh5Vmt2uCYfW3seBl6z6BG4Oo/Cb/fn/fnHH0FxfVhqA
dAwFUhVMSTgTcCh2O1CJn5aXuzdJlq5ZcWXqgLrZAJ6zXbZHZYgtM68SSXlWjka4LnDLtLN4L2xZ
WuvGB8Kj6iBN4GWs7hfLo/0x8NWvEiyPVj7evawGZnxfnTWIUAcM6y/2z3hjB54kUNrsHfS5Rqzb
rNnd7jXdWV4ytpq6fbZxykzSlrkIqxFqhEzMjq+0nsUvqC7inDeAQ9drYzcAkcwm232ZYGyqnnBw
VzNnCjGuCYEiJxXagUm5oKC7FsvLWJvwS3WfTxL/Uwkndr8UCmXOSSIaeL7tP+QY+0cAe3VqGuwK
6C9kf6I6/Z1N+/hc3ZbI4FaJsPbKAXweIGY/EfEH636fjdSDAXV1x/JdoQGEIZH0d72uriP++2+d
mwPhH2Q1tVNANpX+t8bv0v4d+Ok7rW57/k3IQIjHbVhK8ouIsh3T7sj39HAwPUD6FvnTawMc/f8p
RH/k+2268ENBdq7JBicGUHWRR6qRBHsAgXpFAxjzFv9NomswDSUlbLAG4dKZUCzkC95R6u54h4KM
2MF6j09ivccn8tQS5iRzuDbbmUH6LTCw/sXLhwYosDnIAo5P98k+TnntP0q9dhQ9B8FEH5XrWa+D
gC9zDIP+LYqgJSztnpC72vnLuWAAwHzBJA15yTR5kd52/VZNfaJCp/nRsc8hqq1HdFJADKBIUxVG
LY+eqwenzZowoKBLP/q3tYl5Mo0dviaIOvWAHOTFft0A+gmfDXS3kdObUXVClYqnQMOuLltVBBDY
OQ7RL2XvGQno/VTGOcTlob1sRJXjKTzOiP4bw6Ajx5C7cHtBHL4KLD9lZwlKi6Hzhk33YwEna/w2
qgclqeqcn67nFm8WKjsxNEvw4BjIHw6zkF8jyVrxsZvIzjKIl1w798JSmNPOoIm5v2VAq9WcwoRO
/u1taecvSYtK6xugaXq/vJspHIeGzl3zc7zdiokdjUDBCA+9InprV7a1jjpN50z/zJyYrjVDQFEn
RZVNpkCsvHd9yX7H39VWBTwdlSjPC/UrB0BwiDgnHX7Riga5/fbs1N6+J2lQdUI1eB2owfCnhyOt
XSSD/kXaIL18b8XMHZaDJ/Fc0qnalbkfK11l1N7WzrlET2/mvYF2lZtjlZsj2ZwBq7ywaFPCnktZ
P1coc7+fJ1XEQ57hq1/ygTkG5JM13E0G0F+0UX39W0T99+KznNMxpwD5w12BVgqgoJF7HEohZZY1
hn+1DyZOZxzokXjYpnhlHwc8EFXeYx7DteMPiPz7bXTEvabquG2lECHHLnucHZwpdOJr4qtt8bme
xAoEGLOFsLhv+Eo7yRylfxDC8I/zny/A3kz83D4HeWtbG8zEkpibCX7zjqoQG8VBc2MSx/ubsVGT
SrnwFghR8PPzUv1yr3Rjv0DnzpqmrenM8PWEcbwmlP1bFr/6yc0n1mcg0WSIPdw7YnhhCImBvW6i
peFTXy8wSPlvLdkbuKMY9tXcPuDd1lzZ9HjT1DxUVXCLJoE4V+2e9c55kIuObd8lNtQNydWrOQ77
Z3ktZgD5IrlEXrv2TRj9yBtCMmLDiyfX2gVnUQ3HqVEEfwMST5222J0ummwRtKRXjLXxR8fUQ0Iu
Hfn48ttK2Tfq2nGRK7avcEg/yFWcncj8Sfvvelf5unfOznGr+aneVsvaflUUY9Rzl71W1AIHku+v
9Er3lbGVm4hBgCcM0vkzjPuk2mC+rWhmFZYlv0QcUUqlp1cDtMDl+pn8SKH517aJ+asLCAmuqAD7
OvYuI6NsxcHKRvxXFxijwEK9qxXDf1TkPs23L46Hgp6WxURTyX66mcMUMQ+BVG46N54kms8o20fY
ne8+dZlq3Bm9oPmRc241lRUhK0mJ2L2w6wYoE+Bwq63n2Jf7hVHGDgN60SvnXjojeaMkm6jHbocX
PbGlMS367pWeZbnSM2sWovDc2cKgnnbwJHDp5w3RXiiRR9t3o8DYBqUSgIilsiKKP0e9EWj6p3Gi
CSG5C5Vaw/untS85AuDO3ZFT+x/VKuJgkcuJ7jP/yzGrR4Iyx7KshE+2vS/mLXxbDmjEEH7PBFrT
2NGqJUWffJ4IA1+mBAingg5Ei9sCqJ9LRjFgLSFh7ANoftt+9NLctkiuQHbLt+M1Lqs5bTcnCFaD
YXB4rAzXnrZzPr2OuUvLHPYoo+qhN0tn6fY7qukRWHR2Pn94zppM+lz9ntAo6p4FudisA+bHgv0t
7dNk0wiieo+vfa5OXxCJ5R2hu/76qWUJV4HrVVKGBvbDngqfTQcrqoHhmW7/qT9mJGr2/BwtojTg
uwlD2H28a9XDV/qqrkF3Lgb/bOdLvnmvxCSjhVY/CyQjBZ9LASpmdiU3FHalTvx6S4oeyQ2y5ypq
6yDppfS2MSohS+fccq7BaBPToc0T2PsVk+hJpOoeyAHTrpiljMrSjtOOCy3fb+HcoPJO0LOsIHBX
s757mz7fBenzRBdSAmWkihBpziGuvQ53z3NXqpmauV8BGWtLYtlmCq8EX1lMHcGmjllMNnTDgZZ+
FOk7Qp/Z2JKy1BLwB/djIk28W0Ye7eLkTmKRLp13gpUmbgYU/Zxihfc0Irat//LYmAhZEkCyWDYf
ETHSrblGoRMHVdyHxz9Xnrtn7Ct6RC8tdqnJxUtDY2BIaDcrdEpA0Ml5KKtioHLUpw3vY6o9gmZQ
L0mN61nnBD1jS62h
`pragma protect end_protected
