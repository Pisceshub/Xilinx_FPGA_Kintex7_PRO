`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16736)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qBDm5wrrT7e8nIMgL+m2k+Ml+2MAhdJkcDGrDQ9kWXhIAYArPBlVRX+6
vgdhrU7IfKIdZHNQ9/hDG32BYzrlRV7vzFDgmbWV4Oam5naZLndgM4v6WdAE/T8fcz4IbeXlCelW
Bf+1MzP+z8yTZExk/HUF5FfBhTHNaVfwhBJfZF0S6kq6hljlCZ1CDwlQeFAcVu1v87Th+H8Z8Kep
ensB7kj4ri9pVZ29eVrp9LGU0BnEazmb/9TC3xadmCci2Va9ZtpNF5z/DxhqAqNGIjuhmBF6PLmo
JzXF8SHcWcRA9ZDdh+CkYn8jl3PBUFX8azmCyUpyq5jjN/BE66ee369AyROh040dzvEp+h1ujXKJ
vBqrr9/gYIq/7Ib4Cg5QekptNh+1VnftjonhYekEd2Ra5y9yHiwhHTm+dvWq+NYe8yWTuwfYIylX
dCQrLd2ch0wHHf42sJGJHQJ+jIDAUcAHUxiQjVUtWgRSJ6JppDvm12KYmMpjWZa/l7c6ZWZyBsZ/
4SzZw+qegILy0Wy0B+42krWLi8cw2WKq9FWR4mc7IwNnMZY5Toh3f/U9i1sCHtNV7QVItDIoYwSJ
Ja4BmTZMLVSR2EOhZxqfpqxAfYNPwQR+eGZNT7BCt9TkFuM/k3xEq+70Z81PizCDn9PYMRpdpk9Y
GS74GcJ8uaSXCKVAdJfpVGQWI4nn+JPeeI2J0oSDfDOJPIw4dWETief2GYMNBL+zZHJRFIXD9+Hr
03+Spg0yZVbBGshTWIE6+QTUEE3uH0f2LoeHeHJWiPxI5Bx7rNxEpMgOhEGJcMCe0RRbdAzWASjG
EaxEsvruA6+JCfzX4P0SYAzk9Y+yQRjfF5K/Rv16OTGsXJXvYOiHCOn2QCukHubPETlN1isTuvZv
Sk7HAk7o09+sjRfBrJp/vWoKs+Qb6/ZIvJ5uBV7P708qiajVFOiwQVQIritbymER6QEcztCj3G8i
Vwhsq59dxTRaccJxoQewVGclBhJyMR4V+tB2SStTc38vQjYdF6YN953gX3Xdn5IuxY2K1w528i46
5wAyWvvFnrOKPUJP4uzU1ztOxc0NifWkC3iBc+PQJnmWNQd6kUMuNJtyjrOGnAhb0smTWXWZiZiD
nKEM8r5xcLL7IkozAT9mJqJ9u46h+Pq3eqpuYG3zdM7T50P5TltS6795ApnsSxHvTVkvA7os5fDc
RUe9pukAvzAQfWl0qPybglFjov4fH5a8Ot6zg4FSKwXbUTA7UD+mX70SHISSQDtJwjOWlQ4ZdZ7p
DxJ3ZgVWMKesrRYQ5fvZKofhxLJyr/Vtnra2ghE0Q7yWCVdMzQJt++arOHeQlKkBku3MgTOZhXET
E+Bo4POhiZYKKhKA2KxtLdoSUNH/Jr+1G12BFOYwM1L++gvPWNdAuPnWUp0MZA3QSLxbK7UPNtv2
4nqcPj9WIkLDP41VImYg4stnTHYFCH+Ml347UXVp5r6nGtgNfDC1fyEPsxZDr+Ln4KqqPDiA+r8j
updzvdPCgSqakq61nQixMo4BJT9IUe+c+iP4b7MOEiBbMzWuzizGajxkQRkpfBLxxQvRhlwT5BZ5
15aSu1LbzpjcJRmtSvzrtIa+VqgDAkCIr4brsCT7qgeo6JKutXyD1SwK3oCEGJS07vSniYI/x7hC
+bXixAn2VfcyjEjkGel/cp/Yg+KG7r+OBgokyzWUSBG9NPyqCHImLOinl6OVNkSEevrlRwfM0mtR
Wp5eDBSmu1AYNVDoB5+rDx/jxWAkPp5Uy6ZN9x/BrXD6sLz25mm8Lh4tf1JEwpy5WpTW56ZaHdwH
nFHHYuvKifHvrS7JI7V7vZdnag5kOdLHt8s/4LkfpFpkk6xYlm/jau2duF4HOjgvXUss569sXkqR
kCVS4QIJE1+J+r7PNXrTiIIbcHoCSeKsob0NDHC9GbtnOhS5+/GsX+VbhyCFlRHsf21z1AklfM3a
xoL8ClzDzuTjjO3wK/pFP6PwOdrecE0WL9EDdyOMdloe7COI/Atx4cTO7vIsqgiIqhb46raC9ENj
oG/G3xwPSWB89/cCfMV4HdStbu7bZZVsqWkXzJNB5q6Yz2L/ma8+sj0xTgIPz2jEMtzf8RIQnE8n
zUZzZMWoOYv/d9HJ1oLYpiUuBtNI078IEcCk4FbI2sJOe8mtvGLeO/OoP8qajvwQt0Q/chXT9kXW
xL4TFc9nBFFsHv7IC40cBI3RCi6BW2N6aOrI9q27a4RfMWZHDEVnb/cleUq4RRC5twaLtc5gkd1+
KEd7v3b9zhKChsL2RWwDwWVxg9tNM7+Z2tSYTZIEV7eiXu1mQe28sd1o3v2U0XP/et2BsLZvScl2
h+fwLFMiWWa/Io1mFs0hbwZ8hoqhSbDpzezAkctefDo7qtFCut8B7NIRC60stxSegBmyZzS7WZKu
8NFNZCdwTmbTdODXJVM66WBEJMjIJKxSCIRcrfs2yMuP3L05HsI9jhy032373bk2+AoJ7woRU+ZN
jZ/QmCFI2ZYlUP1YC2sz9nfmOLisXcCUYISFz1Bpnqt307ExkJgRk3fPLy2nk6pAQxtSwkCbSdKq
SLg1uYkbSQDgnHNWa9PsLeNCtOJl720AXb4mh5I9RJW1dEWmCJ4iKkvLpkVU/Yrdd1jtiTyIrLX6
WBY1Ze2Nj3do64HaKSDJ/9neDyWq8IwFuF9CVksKq5P2dmcoQLPh91duHw2OFFcBFMBXQ240H4b8
kEau3usc/w1DCnIJ8WaIYCNevHYSygWQhD0i1UCeB4B3l9I8KALmlO0H+9bt/C9kl1iQyjSK5E0u
CMN1HKdUVGwYOHyxn4J+uSFKSNOsFQkTj1sUsFt4YPvtnoa8wRCEug6P7+YHRcndXXBfBRtGs8RR
iJEXwdTjnuMFIwVYX693Kf64mmM4IXwNacZbqNeqCyLmjIitCwjPT0RBR1gEtw7QzKLyGmpFa1Mn
7d/N2wNL58Gz9aHt9QQXFvU7K41utqeeC790zmtAD35cs8uzOUxOd3hDHYsHF0iUvlNPLpHW3xIM
tReaw+l3jD04FX7LXwxjMG6SiegDRLL+FtZsKAPwigWsSzO7fcrOaoTFMToSNM+vFVx55tkz3tSZ
bZfVenLdL6lNd1/pL+aIHL2ZwqFpPL5pq9Lz7GyHTEkbA/ta6XQUay+g/aHBRibS82JQuLfvKaHt
KpW4iqzunDwZPX2oQwCQd5btAiCcIUyaHrQf8h8v3IR4zu2fO5Qsi7HRpbjQqQj2I3EHkBf/ZoMn
K6W/1jwhQZWpbDBxLAosqgGWxyz2mBDv2ZJyTMDOwfjkJobjeCB5/LlkSGKOPHCNrerZESUhqTme
OJrTgZtjOrps1rgUf9eYJ2hsOM/kjgRXyiytYevXP6g8WDvAV4zIq5W5R5yEwNXHZ8DeTD+Gl/pB
EuPZ5MHazDMYKiQ0JzyAXenGU4fH5ppeCpY3G/0tpu2tg6UTnN5zb0xytJ9PxCXM0cQO7Sfrsz56
MVxkOLhVUGKTlXT6fSy1RawJiV2JM2W0MloHh0XBr+J7WtzWFzWne3TwXlBFPz2CwRnN4RQRQGfR
v95d74tZRjJgyozlimUOFMfoYL2gYKTo0uIcO+gdCSHsO3b9/wE9Y7mFlgxTtWoxGaMHkiQ9aOrG
tuMoQEIqsQgiRaqKVw7KtnhTh4yOAFTICtfI0kjdsSKjcuWxSfwMuthIyHlY7Ft1Pd/et/IIet5A
8Wqho/vOpowwJQQ4klEuv0n9FK2QGp0ltNJyqwI5+yIPIc0qwD96q5kYmAYhatXM0ttrAlHNJzRW
L8cIkq8cyDYype09eW+dpUrT5i/3DOzUkUuUT5lkC8K0vDIMCvLcTwWAh0wS/II2pPr3RWhlXP1z
ExmJUjdUdMA38I65VrTDpHVsfoYF+WY0WUJP/2HjnK2QrdhpwMY5l5eaGc9ZjGWvibVbqNfZsduc
nYpdcUTkS2qqXyNtl9dKL+dnwW2sasD91rmOcnpbroocIfjLfr2z0i/pVVhPXpOrms1Kd4Bb2Vx9
zdB6CaLpYC6l1juX4oCOIgrzFVyW1hWrP049soOF3b2KcuAKwb8pv580hJ1PprzBQEUGmrR+46JD
qQPK5GQydF5mbRWmHpWmwP1kZWwz7c7QseLnXMJVWPsrnbWzCR/F/aKGrA+WFPFSB2ToDfbevk0M
K4IxCSdYqnL+23RHGVBolS+rc3efVT1kYfkj5EZ4XRw3NgPwqCdIxD/250CKxVFqghMQ/fwqDPgN
QCToITYKrHNfY0L59G/uymVLLZurBgHEL64xCyfY4hp3YjdkrdPh0pY86d3ZZ0Hnn4f6QRpJPa//
xkq3Cs4og/6UXOwypwsC81h76fveEI2udT2CcoAMFjT8KKJmMO2MnTXDcicMo1kuue9I06oXwLnk
kbWSvC5f+LNIvb3/VE8pcmgnWmocuGj+bb2s9dJEYKiUdWR1PQ0TK8dd0/atP9k8hLh8Q5LntuTE
M5/Yk1LaBIvgIpFUMp9AY6x2uy9rHckMUzkk0Nc+o8tmMj97toXmMo64o7KLSqy0VyWwQvDfYk8H
bnCPj4myiMc18ZNRxCuDW4LrwmpZ/APXebQCv2bR+MuLPmjjwgw8AF3Nrr/aey/9D3ybMqoAMiQg
zctHGKgyhlaBAJqrOLpiErmfsP4JpNLfakpXmGLk6tth+pco++LhfPzqVAyQmUUElNKQ/C2H8w/k
s6AnoYfHFFkp0VPQ+LZ7kEFcxvVRYLFr6Mnij5Rn61if4v1LZ0j3CW6Y8myVso7HGjShxDVsZ34K
vHYHTB8P3mNGFi1lia5YZemVOBpYIxDH8ncHXxCL+oSGDQ97OsMtjoZn6dCYblNk/nB7CdK8X1Go
mJMRhA7HSUNr8zcjHuU1tGmhxfGched0p1WCfTMyNmmiO5r2P46NxMieMrxbUYeauK7ocIkidbxp
D8oiqYwt+UETRhgD3EPCXp0x8SowHukaDR/6iGHyMCf0rc7SEZld44WC3NMOkFpzmyPx5ACjRzn9
x0xhoY5KrpaUVVsazxDv2TalhRW7Izp3hs7hTYGhn5tihOzjeHwhHJ/1zAA/efi1UsCnwvJuPj1X
FADbmCpZGSRUD0hSdy7SbT76mZR3NojnYfFBjd1XwlsTi/7UnH2UYp5yaRwJTk6XXIGqWeCpWM+m
ZZ8zxyMMCQpFZV1G1yiYhp+7KjTlbj7EAMu3QQRep3UqyPDUIxWK9qVXGBmHzPlJJzlNQzXC+JHf
vokB32dORFZrNUQ3jSV3cjguDpThplUN3tRe/lm1pWgqVeGpTRGE25xVU2n3OURlN7LIhdoF5/6F
6D1qiZ/H0xGMoJ3SUyzubeqJStZ+f8E7u7C1lIiwoSEXDicsW0a1z45j4LkrTxTW5bOill46o39J
09Bpc18+mWBKyl6L2L8RNauYFMtfJjUitFfGbwtytO3ZyOP9zkHiJdyvoAJL/rIlRfVD51QVRpwb
xmqjq9rKDAs+vWBuLTZ+cOI8RoxjMC0hnae1emVhzchQbpgYypDVppLYbglr0uweaSOvV+7e/VEW
421Mtz3/Fcpu78HFs5FLJeb9nf+LVk5h9L3aTdPuB0x2l3TDCxa8uSG7p3fURG/8DVyHLPwVI6OB
gzIC1LjzViSYJVwvjyxMQaUpWIROpfO0O4BJdlmqsGdNpLWQGtGRzdIh7nWuDNslDkGa9Vq2dBIx
XB8VsJBXmBBngXf7CL4rbZtw0cVNU7b1TPr4DkhMtxn/kfxpoi1r/9EYnXjQqxLGoNdBcOQWtKj6
px6+X75TWsjxjk2YJlcdcopVT5eY+fLOq63yMxguVbid1aMeELTuyarIry+9UwGpbN59tRVPiGIp
VbBJYA//+bysdP29kgq9SMUjJW39TRg9pDkyEJ1HkXIhbPXOsaWWl46Kh+mzDBRmHi8+hnutJZte
wSuMha1Y6bODW2+830fl+a3pJxElP2C9Dx2O35aVrqpMwikupV71Anpiq/oTCVxbWJIIQbTWcAPO
6Pfklyr7tNJE6JtIlZ+NfGX56KAsOVO7fsrG41h9ttDCYnL513KSJ2y6UYRGvx4FMu4PIKNcwDCZ
URTq5USR74vhP2Y36gS6WTxQ4H0K+JtzoMzNT04BLDEQhKt/fe2HVPkbaS489EAVOHtx07OtgaM/
hQ4Pgu+WT5jsAK7qf1K0+PApEnXPqguXKnCOzFMhFsdBer3xTKYDmpfh4Z2VrrLkIDX0ykgijNuC
+TZufYcnc2gnUgeDgZ00kYqcpQ/dkvgUGSEhIKtEDYR/Yta1hvtmtlmPQsKDPeXkzu00GTKtrHrX
+ZAH84T5D82F+kVU0dPgqPPSm3yH2nxKo+T4rxvOUo4E0WGFgVrh13dhRG9jwMSirK3SChwp5w+S
rFVQJbci0htl1tvPMjpe60Rkv9IBndQOiKuK1D9vGa+lKeJpkQqGCcyGkGdgbCN5bl+NoPNXvMj+
9mTdW3++jA1IQxwH/LqMrRUmW1T4q9MgwqucK3UBMk+vcjZLNrdvqGRwUldElUBxh5ZlpzsnH21c
Ycnx5uo4jqRh0gBp/HlmQ+oz3GGA3Q3FpwSVqX57eu/aE6J1Ue2K9fZD3za35GoEVComUIOwT/J3
8dJAl2j2RUjNSgQOlfHWMcq+o52UVKCOu80cgmdrTUf7E33kMRsACzCv+BpnQZ9XcuJVgmEspSkt
fJK6ACjg1Mw84dzLRcEy/Svq+yBq2z7TtGi+aIPQDOIZrwT8auw2KNOZlJDesqOh5fyt8XnYdQJp
SB4y+/sKSuGHeqrMf8PP6pV9d7Qn5T/1PYhdTy6p8pXVA8pLowfsmsaOQTph8o31ThNj1N8S1QYj
NCv7AIUdgQVggZZnLmHOM3fl2f5Ygxt2MPM/egokjqdyFc08jaWDqTIkerX/Pfi8g2bJD6/X00m9
ey1tBwO33aKiqXt1LfgpVzy6f/vLDKZu5Mls565ie74d48OmIG73Y8fQSkfi7WHmmvcwyYwN5J2W
dPTbWx0T5tadyFfOuHLb1tkvo4fccFyqCJ5qks8er8FTWit4BSNjxmk0Ug3WJfILegEwx+PRJcp5
VwxLkGFs8kvwxlJqDKv016xLePfM+LFAV7w83hummWPPaSu5oLcxkcTsi7bXIan922yI//cmOjgX
QrlYOfyCTNLkHMoQYixUF9ryiAUBLhT1bCtjfWgc7G1dHnRTf2upUg8TaTNmNhOAe7mM4EZGy87i
SNoWp7AoZVWfPbnljxiguNg4WwhFGGsD8vk3ILPSm6eNYgOipzWj5fTIqe55wg5Gs5FHzWqXPWBm
PkeHedcy/tYvd7ioMC7AwP6Hvvz588WEZ59kcxxkklYSdkzrx2Abr2NaRfibo1z2aaWCxIZYN8nK
kC4ohJq/e5fm3VOTl8ozBS73k4BOlu3labYhQGbQJy4HR1COSCqPTPskfs3vF8CnSjOTLwlJQcZN
3fnL7KggK1Wu5UTiD5EE8uoUme9ZzgMJva6CQEb2eb2r9ZoBNIG4WdyHsKNxyrCkevmLLFDGp83T
/MbmjshVy1+jDsxfwF4ghnytouAAltMZi4IntF/a/vcGHMLxqzRVW7AUCvnGJVo/p33xg4pqKLLx
WbtkQ3gbraPaxWZC2GNyofmAGAEfvUlfYkZmTIM5NRmc9rc2Np+4UIRTeNjUXdc4faoBiCIYxMRO
KQ3Jxm36RIxIrSaRRXH41Y7CfL9G2YxCsy83STl9kjDK1qqo82fA5A6KIGZhlQapcAdG+4JuBzet
CO723bJAqzOLI3081/v1YeNhswpM1toXwIqZU14xbanCf95ZY57SIS/WaqMM+MvEbJG9f2RH8xXi
Uz5q4WMJpUVG8tg/L/QvwOAvhJafl6YW6AsAP3U22Rc3p5aOWfR4UmFBUTnwmdr9LW3bECfGclYa
wontKPpDhFaDT2pJ8jgOqtdi8mGNShaEjbYwYnVRtpSzkVqRYj+GDGhZqT0dn9ViElzDYvHu3ODT
w3CfCYMnqAZaqkidBA0DjqHIQtZC5c4j8WtxAfnTb+4Sj6E/zh2y+FDmp1y54D/Z/T2CmrjeoBLI
FUthbe7MykQmK0Hu8sfTwowtTfffrIupRtNEjXgLqQoWVROwF3Vcz7xWl82qWTAdNwoxogVHWRyq
v0Wr7bEeV4/M7RiWVOfA0/U71yEvAxQKpUtkyOAIYIuL/ukGnpBM6HaGVoqoREEF7YcdwwyQKMAR
PxuYpMuN37i8XWI5bzVSmpaG7tqAIlwMad+jOOkm16GeTOk8dKt6iEQPQ4Ork8mMqCKrMTzz5xGk
kkaOnw7FNTc6ZPoOvRNQ560sfMsOxBT7K78Xn94DwkYqQ/lyccWt8wkJneQ45Ock3tSHtNh30CLA
ezNE5rs11D5zrFUiZvgZTUqC2LhLKt9AvTu5AtzS6YyJImVmLduU2Bdvf6SWBMXhkUKZsTYbMeQu
qhymppd76GSiBuAEO0CR6Lm/G7r/gwSiW8v+HYiPi4qqWmgYACjukrarO2r1EwVCUl35JBRXIdXK
6zu6VB7oaN/FuuL9cZ9dXgjzchtwoZqnh0si8hddnPiRj7QbMfuIhlgHWEmGgpDZWKP7mYzKcqwr
UR1JPyTpwUZ4QFawGY/P3qseXfDdZkSJJ6XCOqQmidVi8v+t9jhIy7o2OWKPnLGlnPN2hj6j/0fX
uPEf7/uNVXggbhaZVjfV5q0//pU7I3vXd2bG33QDZ27tez8S3n7nZJpZMB7UeOqObx5IwGEDWXy6
qM7trcpXieHM9GcPY14h/j0kP+bInxfxc1OZ6I9uST2y7IYWfl2D7NUX2FLEs1qP92PAWVLFhGLP
oPnUoR4uNMhZ19/fASxZGjqgfdko4cc45rMSYtHj2rM9+mhx5zAvfh60bIJmtakuOAID75LDtfC9
4TUOvhN9a9N5aej4whWAnaatvYJ35xIrgzU4aZ7eVtlLr4dxmCY2L6hXvi9N7Xp2ucKf7H+eFtD1
PwUTFFvbTQTsbrswbD3zcQKNubotD/gxecc/1l+n4+A4cGXTcfHVJ86BnQ/DxiTqc1l6KmPXiIRd
ncPWaQGDj3dRPIfa9Na+8HqV+oSKRSRDfZgNrazC5eIycg7+hR3yFXRHx8Yx10m4bMWbCkcCAbkH
8qwu4noC5i7wKlVlvw5DW0Uh+urTKLdpK8HXwVYJUyUjPtNItEXb83I6Ox5k38GmyqdX7fc3hlBb
c+mpccl5HJaDnAyQLvEFPvrqUh6BvCIUJV5YbxUGvo2O5xJK0ucfol6BLVAVdMgd5pHAmwdKf4uG
3iaIUOdrTqS5yHFxnkb9jMsomeRqkRVjjOBLejuz8KU30ptSO/rxvNMz+qGzEuZ+ZO4yCU+7S3wV
azTWAIKyFzJD6vsWCf45KJNOoxugt6l4CVTuHaqAsQsxjYWsKADCV7fz4bB1dMqYKaZpRwvqs4sd
dbqP3ua014TpQt+O3RGLu3OHMRSLHVQ+FZyz/0WViK51aq/Epovty3iyG1nVPNhCew752Lq6Ru1N
RZ5llcExNq0G/097Tk8xuZtbT8Nz9CAXjHvBdFWfY+Lb1LTdQeNaz4iBneoT9aRMrEscfkPO1sMj
vATGy39/upj0nm9lJJsoajsgWfIl/W6N2698IZAv6mGMZoUswKjZiL7FWed7wUtZeZLJnWqLYaVr
iGuW5TdVtvPmOd/yDqENwNe/4AZQ76/xgTklqBOAaEwrlYRC01Yz+dyPl+Evihryf/msTv1iNwDq
jX7d3C/uVAfTHwuG7FK7PzokNL6eHKClwxdG7R4YVODV4zu2GNizXzqzbc/W0PSRvagM/qi07taH
NUCaUV7TPoKzUDMkhaR3lQ4zw4rnPUqQO1cIp0mVdnjWXo33zcDzYNLEHXdkEECT1UVfzQ+4SLTZ
YANqvQUG9XzHHTqwxnGKghYBNMvXpkHTlrtE1xqYpZvdF9f6HdDy5iTudFsdAEGbAIDV2qP+nVDd
J3lizFjbS98SiQkU4BGN7XXoPrBiwzLf0HM26dpJajp/tEi9rrXs1o4oUcDSHbJaV2Ed+TH6kJrQ
17gxWamex7TjFNidQLnDsEZg1eXuNmkDJdre1tQfzW8vAQIihTMIaftcnb+gUVzIinnHnyZZUyMo
T+RDtAZW+lr+2/yx4qpRzfQkcAVipe4xfsA4vJ6BxSQl5Yra1xldyvVWFgK5Cqmy+kAsE6zoJvGr
VX4KqxrZHy0dyB2BkEpBCpUtUPlSgl7t1M+iGLOiIinCWcMhDgxrhFP0AdYX+4h8d1xuM8I5Egh6
NQExG0O/TjoJgFi9lTSFo+1ArL+Js53zuBPuH2Q9wCcSOljkCE2D7AW4NJgAGR+IQVKaG0DJqfAJ
lEzk8rw8EyQYVaNB2JTDgmfvTzOmYTJuzsDvOhUNwou4o+ROpAHm5T2XN71P+nIwFJGtl0Va5yVx
+1eBmGnZ5YAIJSDboKkKP7QBUCil1IRcKrddmaL6H2lRSPMMOM28fGK82hP4VMr7DSsdYn6QQn20
YVfFoRWdw/QR6DZYCcdrg/NQMInMZF+Dwu72Yoi+3bMfjKr2/FOoOrhZVRLkY5KqtH/G6M/Z2G5h
omo6Fi7Z6WeSUT0SJpT2xxuZrBOV3SJysfLbSjR+N3ugsTKceRKTx3v2mHEO/eG4Y10XhwoSiLp5
KC/tz/Vv9p6Qghxa7deHjAoRiT1Mo8L0bglptKgf0u0JG8LiIzNn4SxU9PUaOGYa7M+t0v2LR/kH
sEpA0I2hY7smym06VrNlo34KjoCuFvSOeJyGva8sutNwq9AEedW8UQO9e4RiPVsQlsrEiCCBJhv2
dm7Hmi8jvr3Pf5X8pVedusUnm0a5nT3dULajcq5oJFF9nx2Q00riys+5e18IPVaq9g6u1+B5IKVY
HATVGfHgTMBLeYTPPJ5l2HhOty1HtBMPFftgwBChIiVh/TBdvC35H4yGDshDDjHRbTvz3hMBDWsa
P9Jj+GQZZjHgvXYUq+IuxcPIDaevDOS8SywTR01jbX6zClJDaAs8pOnzH+IHK3qjU42ofXponzwH
6zOl9oGM0qUpmtKX7INI1drIgR5EM1RL3LgMREw6gylMrao8FAiHNrXGipKmwvlAXNASuiZAZKom
gLZN3o92RrKGRpSJKJw6z8lC2PM/uNznd2qmPnC3jwyblgshnhSe6EeaiySfJpuaG0+kcRrkt/mn
L198LgWHENlT4GVaQ3WuPx1Ae29kmtQzak2PV54BKIObzZ7py0alJqg9bQ2LwPKIlZf7iGQUAcPx
CgsYiCBUHMi5nu5nYxUmcECO9VHoHeJ+PqYRuJN/d1i8tcG2MCFO0E7JT+dUsFOBvxPEl+a8eKy9
17NFeiV7W2pHcavataZktN/C6GpKbolWwhP2WENWr5dBD7ripWzhi2ljivbhPFDFSj4AiROb/jgO
bj9ktbyxxtVADZlUQWyAP5nqfZwn/ldGGVaf5bsqOAkNoj6a3lRI3WpN3CNNj9tre2VtJKKDrQPb
I/K0ZKNPqxcYAJiTvmJZpoVkIJXB+12Ko+FfRV8SQGGxFUpuMEl6dnUp1VJGCceq+9IZ3IR14p7I
XgdUbc1lMuu2NZAV71WJKTh4YP0IvU8nVtnDZLVdOsihXCAcSFIHoca35ejBx8/RJACXM0NcPJXP
URDLfcINN4OovGYAp3klm7WwyR9B3Y+Ubthj9fr3788U70MeB+ZwD0DzBeMddo5aBL4CEDIOP3sy
cOswR+bLk1eREghZfEvSYcG54+PuteaCVfxnc65nkQyv4NfcXVsbDb63D2359jO68EaThPbpadAN
3VpKDu3xET6HAzr5iSmvWwHq6gysWsc4aFBoI9+95PzUqMHk6qVLvcJIgX8whWHiJAiqnJdl+GNP
F9GxM32mofclxk7Tjp1GYH4SY6QBRfCUWkR6rUVlGX/V7JK5Ng7CTeQsZLFgc8dzJndZdz68Ric0
67Cb8WrbcyXuWuvkgld546uIOLT/hp1G1yU66wdxd2XF95MOQda6yUQ4vfmz3b50U6Ouf3xNRzqQ
oCgqmJCzF5XXUTinEE5Ya7xGmuyP7IVakIhwmsiHnDUOxWPa7Sy5hSgMe2cixM201qDxM3Ehzu5d
D0WWC6ZCwDbutsvnDZlF576BKgCtQb+y03bXI1WEF1ZdZh5yoHpPLvQXSeVrmqJuyGL/dZu6gZmx
DYWMr7c38I3h8MpnbA9lqFxNFCwI7/759C3j8/l3UuGfzIJ2ttpwFZcMYYn+hc5XuQ2jnyf3Cva3
rnb+9bUfz/5c5dmTz/lD8zn1pO2L0mDhMVhugQD7NaBd4QtGvE41l5k1LnNh5P+xWbi1i5VjL+YN
phJZX6BhJr0FhxWB87tXpmH1GyU9+ObW63Go8JwnVcpRiv84Uy4DjcoFtw+EVHYPorjn5/6hk1n2
KPN1TBvXvaMoRXa3ouF6AccxPcpT0/o3+4+Tm45AhChvmo88vAbMMCeLuwqqPj89Xf8b+0ss/KzH
xMvdZ0QIqtkidtezKP9RFwjhtQftRPRvrt1SuHVZv4GGwWLKsKpaJmJG1rRsQwt5p48TdqQ3L1bJ
+ozluyEMHd1sE0BPjCS13yk0wPBD8XrazRw7W3CbAoMZIIExuokQzjtwYdHgP4uthkkBnkTwz0To
WFkXcVBedWnFpsqaAzylAziz5f/8m5ueirx7PMW5GRWoOlH8D3n+24xNPqSHcpPIw4AGYIXrio7/
b/rvth5g9O26P4OOIbBAX6WhuKPkyAU8VmzuOMktHOM0nGC0VXFTlQbtCJxS/xSCBEc3uEBcpTKv
6AKAZB+8t6wtyfcCWpU1KGxy6y8MMeAzpyZVJX9aNTEpEJWXdsSBmBQoF4C0b+I96Of+3JOXrXvS
wN1UhhNIzapxcXedyC65FNWv1RiQ3tO3zT61hXIPIlLDLDkogX5K9A1uzyCgn9wUP1bbI6h4GsmH
4fJMbYq4ZHV1YUVdMBAyVqfRe00iwg+ggque20CRSxI/YhkB2tPHTT6JmLFdyzhzwCrVObKhBZ4w
VlmVI3jRXBXWbF8u9tj3YpixjAUOqA0azQH8Ap80qBon+qhPBaZXuPQUTfIQBsBT41rkCrzk6CS5
Vu+RlMG1EwMO/QiWLFbbywi/5UzsLUN8Vj9fD5tzzuJgTZN83n5u3rpkpWayw1OkRy2OACAqmVhJ
6Cf0pmgGLt3nxFEzNZZ+Hi4IaLHq+mu7sKNPcyvUhLp4LCNpl9K5rNO17XnGYCJmmYGF5nlaR7lz
AoiM0iRpWe+pUtkRsxskblgvEv+/iqHDGhCQGWigUw72x/4+9hIyBJo1xOJk1+arVRo+CljyS03W
mjRpD36uy4OM1k7Fjx8rFpyCMr8A2JD7UWiNUZ9+0tWqFFtd3njPtIPUVi9Zh0cRp/tMLS4Dn49F
LSAJwWjEp6KwoKDzmOU8rWOt2RSaew52G2eLRR7QNYhSL6kgRgnsbeTnJHiuMariS9Mx/AdvIlwt
zkniAgDBcGD/PBiykQWQfv2X+dWHYmJLBV0QJr4A7FKcfVtW6wlI13r5IseeUBft3rO7/kfEGA5F
rrUsRwtNFJBSVZsioPPfuNITFAzpNvzz/b4aqeeJOeMzjOOEsYdrRGpQItdQlaCK48hawa/fU12L
7vnopar8bX4avKsMhPx0R3mGrYJ2SADHx7fgNSqubE2faz+AjhHCKxf0+fj+vM9qCfXTRUkc6PT5
QqPkFVRud1dy95sC1E5olQlKsv9FuAgylw0i6JHoHYeioQ6UfI8/1d25uJnfFziF8hKWMzQUJBxn
SJ7sQCemtBlkhEZtVmVrVeTs4HwQmhKHGfImuAKcVr8SxH8J/Yd7shBh6DRvOkaBjZb40RIwuJcm
7CD4xgbW0HxRvrvDXLoFuBbfNd7VGD70MabuY4oleCrzQQieMK1OEx/PsvJqnkHZQ49q3AWCSrm5
O/xemP+3uviqqaqB35GDYBGrd9oKEnhnIcrIf0uUY2SEOm2MERqxly1F7HKbD2F1b6m6avFDHvS5
TCB30t8wQYcmwf3AUwdRN6d6mINFarbc8MSRkya5v2O88NvNOUcEZ+C0fFonrysHuiVFhVRNdfsv
AvO7CGV2NYPf67TUOG0gxdeIPRNYHpquqj2g87jy76KV7BBQTxQVs6HkhYElmSo4mnz/PJuzmRUl
M2oluaOFHbpGy0G8hjoajT+u3RFL667hUdzOy8EOU3bGiQ53g4Pw8updbgM0FSOmrHMhPTh/6YY8
+w/H1hcvkLbMqZfGCY/T8E7XgAPxlB3UiEOdbiycc2Ohlj3xqLxdQYxIMxh1qmSgoYR7zvR3f+1R
j2lezUhqjQ41fJPbbe2DtTgVL+Bve1w2uRvXdQAcifRu+WU5WqNEQ4mokKry1VqKW95+g0/iqvVO
eJEHyF4U9MguPnhIGQFEt0M267YVXT+X5mOCxf0SmPRV9gZrvKKDlPnMSF/Le0n+V24wOq/uvmXL
9DswZNZBFyaKs08CLxMv6a9RLrgc7DIYapLVfOq5NlAWJdrBHiPev19TajfAnLFNeSVWIGphrzcz
oNrKKRh13usx1CJl0zSnCgyhmiKM3Av4o1jQh6VCOyD6KHgZx6Jhk2S/FCOgjWgdfSTfKsCP2xiH
yK38qoDxAHSP8mCbAhP/g1Ybv8KHJJ8MLIcBvSezbhXvSdmrD4XbEL2Mu9SkaiB7RMrPqqTDw/cP
i/0Z7+9z73GCd4B0uovSVoVT3QkUNkzChQdk0t+0Q+sBq5pF6jjVOnwCwkRVdLU9G7bvhMYDqxmJ
KHaJMs2Bh+lPr5RS0s+3xoGCGFscEfffoGfcwZKl5k33TmO5MczWoYmWCR38UBrR0k5UlVAtk6fp
en51IiNhXxTZAQJPwUaidTw+hHhVCOyVukmoqtfzP2QkqhnZCjdtxWmmA+viG0ooVKnLjScmb3Hm
SNUKWm5rgYeANks9TDtPsJJM/FBDWi+GBfFoCo90tnKmG38CQhLd+qNyqxI/DJFuKM95u/dBZO1h
NYnEk2gyGhwbolbtWkhI1oQwsvCDK/dvAgVVbzxuDK/DnuNjRnAdHmu3pCgY4tlbeZkKw/se7b2d
ZWAOkmMBdMeozMx1+Wl/4K14gmybWu0DpqdgouNTYJV3H1UbEH8GqNXkyiuDFG/J7k2WpVuP5+yC
kab1l3AQVr7CQg58hMci2QZo0o6tIuzWAILSS5dhfG5iFMEI2WQQl+ewAQhiMPStEMjVQnYxuCR3
Jkff4iu3UY3l9z0ZhlWU8QJwCNcnKrBREC9vfkE22wXewvBxad1bqbHSx1wJVYlXZehFjmMrj+Zo
A2iNIwAp9+V1OqsfLbMKCrtOcN8Ij36r8uUImCeu/V5fCs8/rQRCyGP7ateUi39EIh/DmC2hMQYV
v+LaqmUzMM/MI5TYQ4+pK8VuNgDtnDPPHa3XADAgiC9oXik18K24UP1kN0FNqGQWaFbk6vGp42Ji
gBLULDsZs7SOsWVvTVTUpaOl56zglMV5kkCmp8XknEetXfLf+3nWW3zhQf5B8ZiLEjOpgdBGU2ak
cTx4OIPOtUoY6arFYIBsdLpLa9RnL3NmbxwofqD6fVQkZ0J41pyV5y+RmSmr9ze2uvLUzJw8J1WT
ydvUqZ29h4mBNzdmd6zVA7WzVr3fdMEUWLEBln8o2HulDuDhynSONmHjG8RRGA/efaUHa1APBNlv
SX3XOo4IG/SGf3VimtuEDa9s243/EIc2o/jSGvo2ITz/LI9afrHqTNd8BFK6dcUFPKPeqFb1g6os
Salj4VNHw9F4OjbT3JWHCVVyNTArjMXjsbExSl3CzdW9EXShZpDmz4AvIqhK3Am0wqhx1b5xDpzj
gLEfOE6xUOx0ZqjP1wJ9iHeEHJj91JYfswRd05qgSpA2RNWQKkMT/fFSavrLSqeT4NwHFoez18bX
LiNbbKQUQfswBeQvhciTx8QYdA5bcz4c4Yr+TVYElqGq92x1SHcJBTIW/9Lxco6i5ufnTgYz/TDh
SL5T3AQ58oEP4g+gpc/nSKZ14K9cZU5No2QpXvxQn0Vkh0AVDAy+u1zDIrPb/BZAUweHJVfRv4Vt
v5z75UgKyr0vpNRXPPtEnes1pSu3cwsSgccXmoCUTc2n3DjZXWDWpTpU++JKMYInKsMdeRcViegB
fbooVW1rDhleh726Ehio1Hbq688Jx9oCLhk8zFtXHkEzESl5uRPzXRbuq4AWY/99X8rfQ0aW6VK2
iwpoMfwaSdUl+M1hX1HBQ4m4LRtv9bPnQBBTx3iZB9vXCKG6val5wwPVuZ9Rfv9x00A4uDdA95GW
+pKLqjWxtgsQclaTi5m7PDg1P3WWS/bqfAcSV9U0QqkJZQ9YTr8/t47ir1/eZCTzRnvRxJV2GO+0
TJddXKOaJBRYTvW+AMyQShJFa+s/DN0a6kKV7efiiWbO5oaHARc+BE8D607lT6DEcrDYl0w1iHpa
MWciUntlx+aWjRo8IbDJFjqCOlWvCJHwIp/5FatQfUghmAWboHb9ruVM5VMjnRD1Wj84zUro2zBh
p6kD5P6cjVORO7y2b8EwJOz65s7B9FpnrxUvyRWr3dadC4PlwtucrhhJ4A7Z0KyFEoDg3JwMrpCl
2BMXVl2TTpP8u306Un2LmZfCXvwwpE+vN2lMCZpdWXeQ4Xx368+r6qTyx1GtMk2azso5w5/v9XJG
s9psWeagXXJ6Wdy+9UCV4oEP+b2BGdayhjS//mSnjaMDko+V53CtEq6BUKY4E3uWpOrN6w+VAUDP
TJq/UnfiU1ZAMgAif8beJhkgDFx5dj29rESwLEWDG6BhQtIyrFn3ebxa8AnkhXx9mp+RLDiX0NTQ
cinLsFtTXm72WI28QDXe/CEnmjl7wwfkH9ajUaxWH59MxWnD5RbxugUNW/nXNR2sBTwAeV02RYsX
8nHjJBakCLBM+Ft3aVnYnZLXbcz+TJ0nFlVDPOzoOpZX0J44zbtzoHulEoIIxU5AFHZQ/xNVHZ/v
Wd8u0eonc0SLsehNgSD6jrGoX7E8eBr8STRrkSpHenpTMKNiZ7o/+AfyTix3HNFkUYzvw/H7xt7K
sArNDSzXtn0fxDqHf3wpvjuYZu9norjl+eo0och0fONpeX03oa0FFyVxP/twT8Cwwanf5TpvC7Ku
tMkVhxXglLfD+xwT02T984mgi3qPfg5fhtIWsl+54G/ElWIruaH4BN3nTIxiQbVSiMUhc9TwAfIQ
hPgVei//zLevW0EVZ3GmxSM/b5oaTvP35Kc8miVQsfQZt2S9U9RyC3FKwMOZfZIzU+LgGeZdLFu4
h9gC9Ckjx5z50TMPYzu7iXydYubxkXtf22aWta+Jeki9lCXaJOfoMwkw/U4rlyMgzihfMSVWLXCz
nNeKqo7jgDyF+SUdk1jMrppGdvZwORr6QiO0wNYjidNtr9rxDp0Lzm4TFv2f/IgEIhmYO71oefPZ
TL39usJueyM1SrTMRzk6FyLo4AczOQf39e/NjfSh+RJNahCNwQcHctZlGimm0Bg4yUWm7ELUr6n5
u6XbxOyDLxkc2aP28Qm5C8bbKpEkjlAEsq67sVl4d9nW1o+TvJ/8X6xtvxvWvU31PMlkEHCwd0wF
TSF1ats85iCBPcYJxp5UaOHs4q4V0cKZgdcy0nrDEw2Z8KjItlGGk2tlvnQkGIoLh0KevVhzkMp4
y6yo/tb8HA0gWmvlksWCFl9miiu2VAw2+/pzT7frlG64ngj8xsPxxKXTtvYHwzMvFpU3RBZqv9Pg
iFe2g5+YoMbEpdcetWrhDc5prWnVqRSLvWWwP6btKl1aew64f8sica4nii1SEieD7qZ4IELQ8koR
m0NOzifVVNKytS7rAJaSdAtaJoVu9kWtfCrqSPx2Pgyv77zKCi28yKzRICzp6w4XwOl988vhE70z
2D9mpWsHMeO0knopCyED7IpyOdpyiFZDv5VyPIm5VSG4t6eEg51zUqr5FpLAC1R/JCRkwKKSOMPP
yAR0mTQScRTlIU64Tth8ZFRV8kevDg+2ETeV9A+om3Nc8P66BZgmzAdnthXEtGLz12pAEBaSTF9k
zSynVAJ70WggD5BShFhbqsuX8pX7ZyoJ2mYe6K01fLXmSgwCnnDX01fe8T1fZZxUlKjGgIj6D642
G/elR3E4Bt8etOWiav4KFd4/HjtvV9TzAOXn4ZoRTQjirmdUProV9t5KmpfzfS6Sk7PraxxPIBi2
IcsJA/vZxQTKfDwTY5Jd4xWZluyi/62RsDtA0naT8PEpUMi5WA/aoCt3FYopbyoCa4zOxF96WlYW
c/bwrFamLmN78n4KQMHFgMDLPuyvYgAgAkjWH6gnOdZwFjY97//NyUNMOQwBfjM3YMqbSpA72b8I
SXQHkiZCwwCgF0h1nx/sgIqxp0wcS8vbaGbPKOetPZRgrHSQCrxgB201tuFlYhNBik/y05eflr9O
G12MNQpkUNoQCpPGi0PQVzc6nCnh866Ktsa2YOJnWgDVp+P/vvPLJ5pQGOpu4YuMX0jPi8u4iezL
oPqCAaem1rHp04uK7FptmhjHMos/2WG2D4JwvT4dhKaA+LyOA8GN/2e7rAPLlJDWKkm9Bn5KgaLn
0em5G16esZpvnWwwEdfebwFdrmoQyBnhafQyFQnJEWt8UAcZn30h33Y5zjUU+oWjZ9LBiEwehl9I
sqvN/9gB7nHUi1rzG0MRV3KbArdeB1MLIktHzFDj8ha2fFn9C+AKlH2HLxO6i9vSx1pKf1e7yrLV
9fZXl+802O+P7+0/KtTA50T6Sy7gSxnFhM7uvJqnwy89wamdrdn5n7fSEr+kPLoh3sgl1jPRKHvw
TaD0GYPmDmOBRGsiXYRUhc49NFFMgCx/d0WZf0yIzmis/RE+6XVl2KIGdjJXfyYRCTqnPKP2Vea5
cmJeCi/EfG711QGKZ5wDX75Sw60sFcBaHMBefRvIXdHjkBUX23+BktJyMcqgpN1dP4MWflSj/e3I
FDDzzScwpdCqaLmTTo6TOxT4eUTaZQkHIou839qYeiK6x6ou+Sq3LM86EVFhnDyDTQ28c2CreWuw
WUPz5jug3RNwo+CSEtGVLgxcwBsjldKr7dwctD/7KLrlkDeXTcXHrrJp79Uk++VfIdG3V5fGiP1q
BYRQRXj5qkuP8o3zkQ/62roKua/s1MA1KHa1LWEIVdfpHzF1QRlrIyVEVxnyKYYsmLgW8pSbueKp
x0YcaG2167i3VsXfWcdfviwakdXtKGXYi/XzTA9kPf3Wod8kh/42cF3yaA0r9wW7F09WrnH4/nZd
2PW0uO8rDUiU0mmZJP7GvGLRJWSn8KqWyEdESfeToruZTwAuEEyTCNBw/G2xXyZvsm/3ZSTn6CbB
rsSOgWaFqnK1R9/1Rvs2OF+un/pcIZHXgxG09QYUoGXkQOhwJYbBRV8Y8SO9Wcqv0EsetuubRs9P
EO8Kv/QXnDBpcrONLBZQ4dmug085Zm4+RSSqx90nRoz9XsS60eBI3p9xFiGEhhoLtVddVd/J4cSG
yt/C0P+d/jRTV+QValdQ0C1lHxhRbgUFgpJNj2d/b9E/StEwEEFZlXbA/e8Qgkhl1/84ta08Liiu
jKYc260cySHJWhAjl8h/Y0Y7/M1nqCr+65oL64SYaFsEGiriBJZaFkLEZ85L9rJZ7TpeLLiZLjYw
24xeOZzjxvKVmmtqgM/BhqeEspcvJ6o0qM+0+s/Fe2C+9Z9V4as7gKuR/1hyBMxi+xD1zbgyPmKZ
qP0wQbAX+tKaKJKlhUs/IDpc3m+UMDYT8SyrYLlvb1dmOtG6Ut7UN+kwKd7tnZ7Xez1dBGUs0Ix+
9h51oTMlTcotmjHTScGW759a3kAjRiEovEq1iuXUsrTAi59L0MNVJtKK7SDok8gCasmaCilue3WT
UzqcFZQp2XrgOoNfnXTBe5nqu9Q5kx8G4WJbdWxkzFjAUw97VF8w7F7KrGYQTHemMjzUzcLe0jTf
G91h1HNkGwreSsvH7ZoQ2P3csUwejCbJVrcEK6ri3VcAMKNRo1nx2rnQQud/7NGlpSxblvfNey+m
IR1hEJyfg5xOGx4zT+5LyzKV5TAIBGJxTGdxM6pb4Zw3RwqoMUttg8ISs0rGDlKBDE+kor2sLQ/D
4b41vP6lJuFwsfBKtx84mRglJ2stc6YFI0gW15sUKx5ojFn16YHajyn0uAnlA7+4jCuvPXIex5bW
xB9tfrAdwZtgkTyuKnuDgrFHhSM2dX0lKPexsnTseBvlZvaIWrPd7z6WwdS+j5F1+d2l/Wd+bwuL
w6vfd/X4oWcvAU+E7RMpjbSx6cNZGbjp8kYZ3bAEu8SbiWZGnQIeeSbL5985T5koKx6EwV9nFw7q
pJUB4Z/NXLt4ywyZ6zbmWQmzuZhkaKrqP278D10NacMUGiHgMrhEUTvyE2wVNqKA8AV1hyt8HQOz
eyi2+FuiwO6z6wnFARUtpZnoMtLFUdFxMwRN2m+wiWIkvjZMJ7j5dCwIiiUpedz16nZWutFoucCp
ze15hHN+TaqjOIG2DqwbXK0ptoSSJ1O7YwhPQSWpKX8eTT+fPthFd2YNNuYWqpBczkVbHS9YfNXn
bFy6D86KlHzcSST2/PP/cHOZjrmLF3+qwQ6iZQE5xSnruLZLVQDIUEWrHXwH9wGYyd90+0boEnMn
BM2stk+3quI+QJglymhE+3OmTlZAKWyPVezpfXYLjjySY8kfL26ySb1m//j2qDmnh6aC4VdeGclc
bWAlwZLiVQ4/AeqkfacJ3rT1olvNeU8bvXzOxfnB0XMOO+wpgo3n6uWciJ41edy9yJr2lket8LT9
F+7+kTrHUNJWC/3RqgE9Bbej4lTXbkfnghySKGudx4WSILkfjpr4Ua4tXaJdHPBSPLYLcgfnu/Wr
MKb8FD/wIwVeJRO6csvmB0gY/DH9XYNa/t8vKb5oA7P2hS5HVfVp+H/eyjOIbyWlEjamQZ8iJBEA
udeT7pxuWXq2s4T+sOrlug+eNkUAyxiAo/lKGGlSY3sv89jNW2rGJJjmyiDeIFMedlXG0ckmCkl+
L744Kl81/mehqUY//PF+Cvkfkc2oRT9aOfOe2PL84wsZ85/nPn1WvLcicHY+qA3hyREohVAtQ5OT
4/+wLo9WA10Xw+5VPeWsbM1xHNlFz/vZL0JvjtRP4QyOC5ZJY4XHOZkCP1Dl3Yjpr/NUZbLERr6E
971peiu1L83QkmEw3rNEB/mXrC6o483+dHpBBw9nG3mgl9doeq2G6JkfVHkvEhGW0o/RJoUXUSc7
7GEuKKhgKUxfgsbBHy44dEkGe+vOfFHjEyspcUrMlTJp0RXCwekbflakSBr+O/JGa9GE0qriDH4c
jX290XFtQc68Xi8JE2Yyh0N4oY8qWHdNG0X+KJuJZiMfcn1494ZDcssyv8A9F5kGqqRUMfzHhFfE
yKwKprO/m4H8wffMOmFafY/DDL0lVqOqUYF+Y2zNoadnBq7nODP9erES7qWXyXVOLwsz2s/odIZv
cC0/Rm44mjC/t+wa7mGYA4DucWLAq+2nCDxNO/rbhwS8++OR2aCy+WRSaI2mliKT+0vtLyIhmC5y
lx8v64Vr38VkUO6H79zVaCAcQOKbMYIUKgg4PVa8dp7oMyTLqqhgcDDS3iOZgDm0Yl9yN4+ddha7
fJ7D8YryWXNNdFmvOpBsG4Nwp8f7hmNZ+UE8RI9IL4XnzpeLFxlFgjxdHFseWhe/Bx4f0KpxoGD1
PFJNx3dQ/c0Z5brvus6XsQi6lo2MB5+JHhzSP5oB2bAEr43CXLc3Zy/dRpHXySuE+IicC9z9UpHL
jgnS01ITCI4KodpCAV0qs0W/usq9RjFQvNS7ocezVuaxfBSpoLgW0rVidLA7N+p30Vznf8VQq40N
62Qc9sQa6hwx761ABo2FzAoYhEPmrc0sAQVJDy6fYP7yDpB6vkny3Y4Rx2dHNy25xe6ZbjKsWMfr
RCokGuPReWBQu/EuCe9RTLwd3eHzN8BMxqCzZ5A0Ul1plesdLWzekfsN02IKiVFG3LxhhikL6UYt
n4g8BDn46i7OjZ0Xib/ja1hGVqPdl87VwINEzcbws+3mW4gn6Op5F0N8vAop3pStCzTocPZN3dE1
wiedQG5YAj/Sr9GGpzdSuBI+JgodPTx6Av4eVet7NRsW2JDVydmTeI1yZ1jzm70wUowSzfCIch6f
D6am4i2b5WRgGncNNqnxSE2kcKXxAxXTAUv1OjQyjqGWhD3TVy0P7KXHSYQDtO7RFG0Cxa0batf2
PjSLqXXEYzCRbFqryGY13/9y4oQOPjoAh+m4VlHr9wFwA77jV2Ns/9YDTphdFUaM08i3kb846gd3
h3rJ7IWya5FfNHjHdyOvn4JPZqL8D51CiyygFYHU4p6xFGA=
`pragma protect end_protected
