`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10432)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NxONQpWmaioFGzw5JY31JROvens7IFn54ap
yaJP8qMhwIH3nvmxbnaOWWS9cSyuihnoXtbpDTUBcBJ7255T/yd5TiyVcKhKvZDP5YbWc12b44Gj
u3n9PxEmBSOY5V2ZVKsJv3Wc5dLFNc9nq+M5DBZvu3uUGEny/THFKRhx3uMMlnqJGvXz+/L8UQmm
oKise2uaQCO1PSmDvRyxiQyOl8uuAW2SDdMYa+kGFwajQfQfpb111roUc1FXWeSLKwL3OBz+x0Me
ywGVUPwDMX26bPUsOY7YuJtYzQg2hgfhCTpJrsepH86MPjNaMqcHQPM0Kq/FuMw9ZFpqUa64QyXT
UMoUJi82pPt9F2U5afLcpVTjTvjAjQPYa7y0Y3Dh4A9awAXmBQi6oclqFZ8TZIf5ZZ9Njc+uymPi
CT/dbTUUm6njQT9D/mrjAqn+DBemp7tFMPZQB+9kuNc7xwdsRP/sPnFjwPXvlUcmV0Ll9mhyOD8p
jVtnMtiIBdtVZuHpLJWLzSJwh/a+t8iYvNu1/UXqw99ApQylvXP75WEyeA1Fe1lD+hwElUTqU9rI
qoE/SWwcIDXXSbsrUxH0UZqhi7ZIquNMG2xz3iAwYGZYyY8QmYm++tYBlJ7btrdbG0ZgCo51fqqQ
WLAilcEzJjZeDgIe5KuaF8UWeigEwtYaNePjfkwXJg7Gh4WcDIWHFJ5id3lcwNKKmI03vYlEBQqA
zRP9asI4QG3XRXcdcrM5+H5ZAAkbbs77XRx4q7TM2uRL8NnItLFiHphg8UDzED0lTU5G1Mx7pb2r
MAQDsCVxZXZR4XEIqAy7WPn2luqpqGaoKNLeI+rqL4dt/sC8rnP9T+ES+jv2U/bQ8/4Cxhw9fg4E
oHi+X0/eS3dvP9ws7432fM3K2OCcC2aD086POX/cIbpi8FImfZ6k9AKeaP5+fCr5LvMz3anlnVrl
Mv07kMFDBUV7SVc9AmSvhR/f45j/jrHnhzOCFC3AzCtTDgRUukq5+KqmnnH1BRaxxski8MjMwNl8
TCqQFUMeG1cVRyNKboawLjPySt/aFEjHgoAPLk165wr6Rxm0in3FTWqi04YxI7R2FuTc/nNhU+HP
poWyjIW+e0tV8IjJF2SMNfHRLLAmFngbd9KFosBRl8C4+vxDQkEURxhdFegdBw7k1Kgnpu8Pjk1f
bTkhXWZFDNIRatcnHLzwj3tjkg+cagoyLICmUHpk2H0oTgtxuwR7WSaP5WJvotHlJVKcAbeJtNLS
aTD55vHk5EanEoVF+TRiwrBNJi2wOYNnW4igGebiymzlihTWDVHBK3v2DjU1xwWKY3mW1S5R3Va2
fOEY5miSsq2WdRPLLT+SR2VaTCw5qs12o5fzbyU7/Ua1dFk8MAaONUbrjQXziRpe3Bdei5rrpycI
05YZpcWwRNe1xgJqJskYcg+TPmARHkRbcOChUjAQvzt/CLB3gtNRkmk2n3Dc9UwNMs/WlqDVPNmG
nLdCzUbnN/BxbYJObOr66c9JuUHkyvueZ/7abzMPQ8ayRHmX1fN4hTSLFBqKeySQ0e3xSlW/V1bD
0dSiLwaAUgGpZ6/8uS0FsGvNe16NlA/K1YjYzzl7S6uaoxywNUsZUwOrxkAz2yNr98j8/5xDoe1p
x2bQDo5oT6HCTLEvOdhM4fQr61Q0sOUQMXFf6ZNNfq6wHydac3QPRzUUH4z/s1FzabUgw6rYgEZf
EmwVmrS1MEcFdaBmmuN4k1ZkP/U1sBY0DHDTu4TRXE4ZgK2vPDNV3MsIHx4Nlz4gVdDEgaiZzpk7
kl+tIHESW0fihv9mlRr9FbohQzoXI8txlCZDaU2U0nroBz1MFqD9WB7Br867JqOgP7u+ZaJZMN/E
b7l3WoZPajwprPIwJlkNuTVczEjaj1ooRfwpmFQWS55UrKnQ6Xto7rrSJHcp88OwMnpz6bvI+7io
MSkyh//N7o37BCjZlRoqyx6PpTL+70hbQwZoq6osZKGMEVzo+ef3ki7eTOTjZAK0178XKq38PxDD
7Dm541vbYxNTVzWo483jYqUDaEeR6y0n7vtHdsAZDAwNURgMlmpQDkfASv9oAvpnCPeJ6eH7GTJM
RJveN3aGTXLFKIlSPG55go8wbUGPd9nlF/yKK/rBknkqm0PoQttF68D2JIbMTpFYdk/R1gFmeBL6
/e5CdI/XqvBZxekcytnL92PhtyDdBldlMIFscsC5cFCJQtaUyT3FDK1FYtvg3eD4rcrcM3xl79qV
L5XUmHvkdBjTlUzODC98uRVutC4pQPO1Lvy35Ndg+kTTB0haLnvhWmfpTNrtl43GZlXIn5MT6WDY
YyCBfj/rZdTyQWk16q+zVMqQ59DMjrnbtwvXN+s4pof3UUPI7z9r/v33/KSEqxOVK970QjuAxbLz
ChoXs/ffu4J5pKJKHGVfjnbiyOzso09A4bywHpdMCAERCLW5hBfFO2DXBIIWuYUgtrSzAIo5EbeO
ss24MTYWBP52Wy6hmJUinvujvCOteqKRIYQjMnRk6kYNdhDPMymXh7T1ECqf+JUHp1dGrqDqxvXv
0ZP4jS/YuPMjqD/P0Y+L2Dv9z2sooVXaOHGwYEnglUpVtuMlIybefWd21zm2l7nhxUafvde4EGdP
zuddv2f4EhYhxjCovehmh0zEaVu3EPgBABXwhGjHuy16sOn/uPOEPMARyeBVelT+Z7jpDRvLVDyu
tFpzPiNS+vaa9CuaiavXCoDHojuYKB2ADz+qh5mvXQqJM3mHAQm7kf48ys/9ujqLUQfZj8hEOj1L
LuL0aRYF+4P7bV2FITWSM5IVY2k7HebCluxXfXCpvqz4zSfRbYfKWBFxpbZZ26Dl4BYoc9pue8yN
1ikhSxNaS56W5nq9cojZ4BsdWXEhjMYBNAUW6Q9+b3WxDydJkipe6rbJCxnbG2FXr8351uMewaLe
FCCC3Gm32X1ojwW75wZdKA+ztDrSVpY9dC7JJiT2L9qUyk5dO6U8gcmAj17SOWOWb/eFCx9zN+T3
ongDhoMVsuk/h/dCsdZsDXswVT3nTv4EjIOfvSEFJEk8i6dB5ZeQ7hM3FBPaNpgLaLZenRbIoUkJ
NemZSKVnXYbk3dsnJ0la80O9s7UmxaHDermelE8KPBH7J/RYLvkApxz5owt3M80/k3tIsNL49/z0
kgkoyrMvdjlljLpbwrn6p0EzCpyXbeb6igVhic8hTTdxg8WIsSUdhQDB46hupsicvSpv10wh6MiE
44qihjlB2o0SJPdh1W/9elG6sR2M03GmL0llfbTMEuctptvnaprcmMxJ+A64ZuzXvje5gDKfRZHx
efNOxCmlCB+ZjT1pV3VEevlGKuWElKDAHEJ/Ppom32zVsCyNU4aofmI284I5zPg6AW2lo0D/qn0e
TJb6IcLGx67o35kHzoKbGV5inUem4RudhuFlB7JT0jPrDlHgqMmVEarxa0aymuxAjr3g0emLmOsZ
qCAGtUYas1IZSp50Wzlfv8FH407Z7uftxBIc9TI9AvCOEa6J5OEgaorEChNzPVMb/28EG0VtO7L3
x5sB/1JF7Th44oHGVuhesjRwVDB9BeS30sEG6yCsjVpeo2+nVPeTQGs4rTZSOyfKX6ru24Q1tqYW
fjoswM4tJjHEo5RkqxjC8PeDz6s9L62HQ9yl0df+3VBbuuwrlfEn33pfEm0rU6GceDKsx8aHJ6/S
Gg0MdGBmjOEHeWzHJC5pqYsbePeIAsWeH0AzEdrkZ0QMq6gsuc5wdMX6tYdxqWMYm/SQlRUbUT5P
+Q/gFpYgOr1hU/iCj3gPtreagm8yu8vyCmn+SWL/xhLQowvKYRfEFGLmjtZZx/RRIrOLFyekZOpQ
l1HKciQJY5EM0AWZIVBjwMuzXnGGJOsDVlP3qA/AQXmGQyi0ctTsAaj+3DrbMp61+k45KJ7v8mIB
5llAzHweb7VJt/bRwo+DoWnM6fZ1+e2bz6JkqHFaFylkFD0w9YHKud8DTNu9S9qyogSKU927wPKI
lDglJ9aLXE2fYL9Al41/+7DSyrkpbhs1cHPPVRd5v1fTPfkGRNxdHjwpdfxP+22S1meW7M8Qzw6G
z3rZF5tk2DeBLh0rdJe1zQF7bvuLfwwVwNDFZkGTDwkvsNMUnaYQKooBEIc/MXbaB0gI9T7QaEQ2
jRl5X9C6ueUmjH2JqZzeRMk2Ilbu6c675wj2PnTEFmVAz/BvAxU8xpQt6mJaCl9Wc2SwzWbXzlFE
ozjcRfny2MR+XRn3QHRM2Um2wccpnVj2VKF0YNtJnCDqNlQGSGsqWbX5YFIUDSkoo6jxTPPpsXM2
4jZvjNepItpydTW8AL4ZrsuUdvNbsOq9H30bVOZP5ks9al66tXoi2igc5xAE+V9mZDAPptHwy9EU
l2S7phWFqC5YWrWYukWDlFZ658x5fCovZ3uGWgM6kCJmLHHaAnFgEqqq3yznAT1iaIou33jMBtGd
CFulPZ7htMKHAL4vgu41HYVgzyCBUUWWMJW+eLOQ5FJb70LXwFBA9kTJpppSXgE7ObCaqfzt/7iQ
7dPE2FLjeitbJVweZDT62rIfl7Ga6JQH9AWv/B8jUaF32JC6z1l/JQxZ75DJc0Lt2GpGI8zyHuAZ
R8+vHp5WQR6qlDtLBb2ddqishiLglTE9VbsNfl+Po1N1r1tcTrG3k5s0623zjft3W0W8lY3+V2Rn
lVN6hBwNEAwFJvv8wtYFWXaLn88/9pzQG4oT5ldVCxBlhlVR0EAOP1Zx05n1hKWNIvsqvhn8QUiJ
kaGOOI7NSJl6BCQbquHjyKzJv9YmnLLjdDkyqU2DwDbJVa2ZCv4NpwSPy+4HKUmJ7F3bT4UXAUfJ
7tK0tDRVnYKAUVr3m6WzU0v+UAetDrm2t27Jt9xUYmBJGN014z8EaSfg57si/gR280QodKh68jBl
20xAFn1ZbpwO0xcHLVpvaHa/kUXkbIAkmCxvmRpHD6JN8Tlvvtg9PP/7KZ+Cd6+wNdyx+gOKwPbK
2SnnAzID4N0y6CI+SoeUtVjCYudX6QSziO+9U34BOxhvS42ZmMF2z8AfunQ+CHdhk/40i84r3eqq
T3fRdfMASRwFf/uYtqIOaudenGzimKZ+hMpgegQOYb/RKPnFVah1b6jkTHH/wx7HPRLE2CRlfEMI
V7vdIVq0p+CiO//EGJlVS417+/4eLwmC6g+C5Q79p/uau0NuxSnpmyaJdk5ulBElOC8ENqjBfhZ9
ANawYJGUCW3hjgZGzGmLJ80pXcwOp6TK1G4UE0VDbcGxj7Qkp9L8Xi2iH6oDigMPMFHTOTH65TCp
3kzxYru6w+UYpOFHzLrpLhGMvzQfsPDuUCR+x1xZJBCkh/ZOoCUtxumMqVwk1qHBKqHMX6hGfTkx
UsC0fz/nA41JKW8t9WGPcbOqtRa0u3b+N47DlVaiZKMX+0uVb0cUju9xiZSVzZwwTQzZPO8oNFtd
qVsCOObooJDkcpZn7r08Uq4UvfCtDgmFuHT8EaVdu17orsAR+NcD4J/xOspL79g9rsiT+R04YpIm
qtCR0tp/waVhNUwiZJcWwA9aiKeLEwnoE2t+sANXzpEHn44kEzDlvMMIaZXYUoY5vsSNLrCZfnqR
ctqVUc/Nr6hdH1IcBkIvNrcClCqp46wn0ZiikxuPXWbflaoE1lYWofXoLmLQyShMtcogma1SaN2t
2LCyxvyLFAOqf9KJTM3FKhziy05MTgVLjwcoI9XlNwuDIsDvFvhXGYeBj2V+foXAnT+PQivwMRth
J/cWnzF/L0G2GKXD6tUcKWwnTtKsz2cpLhwp8zrIHXGuz6mmqhYvpR2u6imBr4Hf9cKyVFlWhZpq
2GvKiLGIqVPThOeFI8H1FFBj+lnLZvymMCn1yTAg6L5KgfUYFheWMFv9r2w+gC5L6h2Klnut7uCs
qZ3id/KBCxF7CrRuCjo5/FgXBmLdJQ2hAW6uO4lf6G+hf2Wc7S7A2Zd2iz6p0hmMVuCKzalNUlNV
Fryhd3tKn8540VbrEn6BLLARuSDHHsfWLh3sNTCO3U/wb1fFbQ94homhuLq5NU3P7u+iJczn4EMT
ZxnrQFUHSERuf/mdPiBHAq8puXOfEQrZYhHB5ZaH9Q/7TZDhqEy8PAWykQDJahiN6ko1pIoMvFmx
G1JQnJZQ4tLqOo9ypqppZe0S9eZNtMcfWlX0A053Py4SExuHmJDhWq8fftdftm1zV7y80k8OMmFx
ei2GEZSaNOZMjJm1GxNrBF148OFAAwncl7c0c1sOdlb+ut7vQXTm/rzyqskeTG7osGxH4irL8V7b
wM0eqzI7ejjr/g2d+/VK7VposbR2b9iNL7vDlbPVJHu/fpUY2SYVfwNW17THPRRUdd27PdH5bw6v
9jzWje/nx2xajgShlXtP8rszjVqsDjlGo/iFgk8t/ARPt4XezLKn5nm3mJh90fKfRQp287VKCdWA
MPhD+Lid91Zx/j/JlqLep5s0Su2teLPTtOtTj9qurTqpxvmDPLWM373bZQ7JldHB95gZg5wGirEk
OwCwuLP6yext1zpAUArismWRms41L0JyCUMqYXQQPNAbdB++dyTvk/m1jt/Bjlei6BJWLYXuvFR1
KuwYWsTkr9KgtVwa+Y41m5iOwA2YShGCYfdsTmqYwxFmr82hkC74m/B1imLVVmVr6dH1o4+zJ/Fv
PzYi9KzrIswHh3RRhIUDuyV7KzIEIaoWWcBTlF+eaiIO04XMLYuW3Q0KeIe29mULYgxK1xF490L4
lVwdkIPqPSBYoFo1jFXbuz/TL6i41wOzsLKQBC4mujQA7ZYn7LpOqUHw/OdrjHr7Q1d9ZTSRKJQu
QlISSSw13JRMfqsBrXCEGylP7j3rDfCyU7uKzBznZO+DGXy2mqXSmC+mMc/SDwqpQd7nB31Ilok2
54dZcVVfGRYX+UCdD/n6luks0TDRwi0yLfZpfJP14rynOQxlUGDdGhUgeQci0QxeT5ZpMKM2Ok5O
L1c4TIaaNdPYBHwLJNCWpjk4NWlOzNdXDCTVfQ6vhuZi5DAmr/69VXXGM1merGTE983Mf040QxAm
Y57Off5T5rmoT5qMlhcdiJLgb/+uuGuFSMhqmYTyKysOzTzRYQsXSEtv1ZpAXMMq6GTiDdBES1iJ
HYXV4KjwlALIxm3uJzQ3oK2alKSYl+bZlHPzqXIt/UC3RWvBjuH4YpCymzzOLC07xhnuzfXLi62p
ylrJ8w08l44YSTKlBrXukFphWqPhAiTMQGaadxEj5Qv4gGTD+RYn2EMDVegzEwxd5uDOHrEjA8vK
CUN3ntFIaRQzuMK7AJnCoxOjpuA+bnDjmVwsrO3V1uIfW6zPR4i/QJep2Q+DfFl9I11pPFEUYZ0B
V3TQIhgZVH2IuHfSdZtUGFBipWzT4Rw5vO7kt448vhaLFUQLIKO5QiHebMygce6c+mQi+P5yx2vK
EMJgPMXCp+QiERhebjGdXEvOF+IQ/qybrq7HWciQtup8ArNrc9UxwK3MHBpGqUL1vzeim9sS9AaN
pEPT1JsIXatnXbafOLON6FQt7N/8g9hIGd5X9yJi/M65mIR45iUYWzrkN2vkFI5rXQktl/LRLXq4
Cxx7Kjt5cq21eAwS7cwPBV0VFdz2/86L02sgBXjVm+ngYtaM/5O1senpOXJhT14rT0WEpCslmSZ5
WpLR3pUFd5v841JCTC06J7KjqaDOK0wV1b86JD9kku6Xj0+v2RUfEo8fRN+foJCsG7TZrn2pmxiw
mMHsRfNdRgsVQxhjXVcoXSKE/jrj0bt3N/MEaIK75Yn92Ynk9IvqwGDEKRxI3kmdHzVIvqQYRQU8
ZISRXW40BMicQYcn8xMkPzgabLnmtxPStLssg7aqPRmbSeaZul/wHe4W9gHCz7KIZSdOShN47PlV
FHDz3iCatKWXy7xJ0wMkHzNn2EjM9DCKAoJnB5HsrZlrZcvW4wxRbFcca4fHtu95rQ24g0LKIU5e
4iMNjJzSCEuWoZdur2euGh/7adlkKmHU+2VsvRaYv3CbrXrfJ0Fvts83pnFkI91UA8zuDFEXm7pW
Ifhvmk1WAhQKkZLmg95LGwVHbLLmKEpKQgbzMh5NeuN/EcYRuk7hzWjUtFrK6Y5sBupOTP1D0wdy
pzZFoF57Dcs6fzP3yLcHnVC8P4l32RA1zlXgTu41PIilnkEtS/9uyscXqLYm5rxaK6gscukB8I6y
uJPSuWjmvVq515hsDsdNGkIczvpjSewrsclcxjH3/Gsg8Mcjuf+S2XWs1QhHCL2UU/MDWQNyvKHp
3ugRAeF3p1STU/q96+GEKFD/6Qe/3y/KhUq6pl1j+/E1RXUlm/NNChsalQlXzW6mIvKbsOn7p6Kx
Uig1csYTIpcIW4dfXEFpxy81LIyvCHiM50Emax9rK8tFWgi337JYam3GhPlxsAXzSyUPmImgg/uP
v/A5d3T1NWl+uU29CGu3N77Bm8+iG0nH/2qEoz6yrhIuTZuv355cMpcFdlSp/g8htho6UQAYZmN+
upuIQxzWhYXbtcl9waCV+XeVo2CQqhofBolj8VcyJR3QtlbMBovC6RpTj0UEWAyRiFFN/h86afdY
3r1V9Fw22WGhy3DA11JiNVHgMYZB/opm1ufB/A0y0xixQtemw7IBWbD1/RTq15Y3+s+oqPBFZKu8
Dr0Kbm7nLnnJ3Ate5jOD9zR468ADrK61CRnyP8MdQwYj68QHV/gE1i+kRN+TpoyIP1VkD9r72Qx+
LqMByOiBKw2VAf5tzTr4oOgLdrXAvTUUABavcewShHnlxwKB0LgB/1c2TKUhCD7CoxG6HQMBIcln
BtvK78q0BBwqgEmAne3FP/4iDsmWhZnTzeJAweeDI99rgC3dkL3+1Lt5UX2dFGjY6LsGBgQWl0P+
Z6PS3d7OnRIVki/jfH1bL5wERp8l/+77bVPZh6szBfGXbllgTw3t64allzyaRdEN8FnQ+PJ+U72w
nacDV+ZixBLA3KqN5J6y8PBKr+L7tz2/TVZhjYelPQw0ASpoTHpOrpJRe4oNGI7aluV/u6VU5SaX
h9FwTEJhowhkyvfaLZBFOWXN3GRvQt6BGnPrVg4pkjVP/og+ln+jDIRBJZNp7BSCDsZul8ApySye
iBrG9Qj5pN4tJJ/f4LHEEwmcKIL83k/uxB69G6l81RD0sqfDYFM28k+O6UzAG9hdTIyFtO7h3ZxR
k8YUXJvwv2o4FVMdE3o63WN8Skh269LK2KPSxpklFeMbtsXuvUMTV5+Rm10fh9pQOwHBvtaLodtI
eYZ+C0nCQwIsS4dFnjNeHSnj23tm4LOuwzDZPR21lb5ershTLhDVcOHCmqcZHYTBd1EmOsQOAU0P
+ZZHqexWCqN4csQJgtyZznxWWSqstyujjwPQu4eQ5Zvibftqo1mbLhlBD2da/GvbPmEWUYk11fwV
+W79VxKk/S9CB3JlfPfP6CEEVgTGoHKrOTsYbkBxwcGPJmMWk/0qcH8UODwsrUBhXOJBE/KR30gh
DJZiA14eXqFGSRyp95Nt7/9CYNPD6418VPM3ACpwGJvnjDbIsZzPKWFedXCwGcYLUZN7Gzh6o6Xq
HI8hldOu6zePRLoF0ICWlYUVg84j821AI/Z6dPtfSbFrMrYL9jSl/+0RLeiZPOAmNVm+xARu0XcQ
ZGkMPMWqGW4omE95bZP345OXDXb+TQ9E5iCzv8uGkvj9qUC0/TVGxYWorOhyaeWSQsNsau+O984i
nD6JmDpScB4YRGn0DZNiA3S+dH6fTx0V78N3by7ycJjrCpi9GuQWkGC3vnqueA7TDkU06l53aAjg
VJrfhB+JBDd7w8Grlw+iN/XmLUYzRbhfgkqx31D4f5ZduOQRXGax+UURjAppHj0eWR4UDG4ERHiF
fSlnfPAYsfrhNBIpQqEDQEr6gZijdt8af1DuqaON/HC4Vp42BXJ9+ZT0r2KQn18o2kf1x3eKbojX
pkEdN5ImSyJq4m80XOqspz58cDNhSfJoEOr6RlNki/hG1QtaHOVnMSvlK0y4/2fhZnOUhMcghoH6
g6cWXPcPsBfKZc8WDkN90we89wbs6/6sgKmPTmWUiwW4kVlqjW6TcwfajjspxUycEskK7ZiORBbq
PbR1rWa4Do0XlX2MDSan/B3woAT2hl5wWOC/c5ovmzB3W3EV/raAceef5ELIDkNgtctbEsmE0wdM
NCgiQsSdffsV3LySOw0aD/xFrv4u5kIqaMWHfNAXePV08x0c0q709oTGCbGKoBofi/v+68n7ulie
bX4El/20sc1THFc8SPhEVa4rMCwRqvjB9yTdz4/E9InEkYXYbqI0Gd+H0STws0Wet7ZCo43/mqNF
zj9mnAI9Ajiy59peRwg1dGWcvxQ1h79v6fMcjAP5fh7m1MSIGHokE/rOtsq3mrLNygAuJ3sWxwAn
28180f/wDgF9F01afRCIk32tXw5pjh18J+PbwEIZkRZB/9nQ8TSw5PBfY0WflFgP5nuoAlUO0C7b
28lTF8lqYXu4qp6Dt3S1iVahz8pWgRsDCCk40EkWqSaC2rlYy5613AJaqCLonFQgv6VwyaRnceHq
PCOkg7vbQCD/Eoq8/YKjaOaTGYv9Y8Eh3RL6sppBe4rz9g+WlqXZTm44n6ZEMeameBwnbtg3v5jW
XJN32bvyBxVs6d9rW09BR/QoKqiCiN5N6NSUNf5BWEXjfWDMEgMDFvZQ330IgvFxY0ZgTgEUrMZ/
+oCCXDAKXdJMxaGu9GnMXM+ZwS/X1c90B7+lce1XvvBbSYnOKRp09jyUiOr3uZnGM4EFZsWEllB8
F6MMgi+avP3QhjRvdHlG6mAgA8DjNhsHDrAbDOO1eJqt3JMIb0iTC6Wu57CLhFJWbYuLF3BNpnWW
LQMwLzUqYFWoovJGIB6rfbZbkyjOiZ+pultecooRW5NLRokW7gzBfntdeYK41fRsVvYLDBs1ABl5
rieyhyA5qyYFFVB4rQGz9UlnIt6vcvbBKUKx7w+S7fmN4vOvyqK9v+W+DAbwqaQOZbEVPXo/NxC6
DQJl5l+J+Xf0YIwfXlpStDPcLhjY/vccq5EkCwAXlSreCxCK9JhJvy2XPI7SLowKGLuWQa9etUUy
G7yJWySdowT5CgmpiiMTS5TpaJS34XcT6fqWr3N0RxX0tQ0X/7wq2hT1Sn6BvLq/DosLcJX8Pbvk
IQ7pz9cschaaAkyaJMQ/Pvk0mX+tRkYnTww++hYEcFWXBZgY2AHEdSo3JUMJ60kLD3ZSFtFdOt5i
qpl+RCx03yJzTAbcKoq/Ns/8TcgFN6hczm5QzUk6tl0TJbbrF4y/u21FsQMmFtco1+x+niBqPxkW
N0+3YdTvZia2ta8itO7VcJMCCncp++eT1QixZdPJg6c79xaZkUu6NK6WDXP5LPiqqKFadWvtUIIf
wkY3nrKaKCft4E54tY4H0WmCkdCVKvkYtLJu+DWS1pRj22MZzN6HPhjMULzd0b86AMqGEX7qpqZS
72nGtvJSrrOe2lV3ghLVLfVYICooLBzLfsyK2MZ6q2RNkvmo0l93vF2m56PQ9bzGMBsyxUJ5u4CN
Eb/2cjqLv/Kw0had/TkJgoazk0YFuuTitkANrRteb3dFB+C64Fl68VCapHVDX5Ss7sYF7M/dWrGh
q0850X+uBY4CdT0ANQ4GNk9bkRqEDTLGB6MuzOqoCZlY6TPgz0hiw4H6oFuYX8IPgR5a6iqKCKGi
Lre/+kFrAe/klbP1glKtnP7N/RWz9Uh16CS3OlfMPmNQXvniMZ+3N632gMoZKIEgQTVGeQli8iHQ
R5NGRGZQsbDZ9nj41763vg8gEJHwQVWk+jH+L1LWrRliYGOEwhqXhr2kBH0KDc7SLyvAHzbWhyK2
7Lit6GcxVDfXX8CVUp6cAMJuq+oLocS+iVif8JH5dIqsoS76rHGpbNdKnQiCSYaJ5a0RNXLa1+Xn
aeD87ToU43HOmqGDpKQzmVmM8FYA8tAgmEZVky0ec89bhaa6DlIcjzurQ6jm4guE4oF0Xuh4ijPI
MTpZDgUkq63lkSlBTZqcz22o4fr8tP2PD8KMWEXQNkGrO/1xS/woXlvJAvJw6vlBI6Y9ypbsRYWl
1yZNQahLuEx+gcC3Ei03KrKeVFPx010SJu+/cZuefuEtI07GwRnaVxp2jx/QwNemkyH1KEQCPdps
tArGzQGtIvWwHuT9FBwcQituuTvubCRl9+6QIMDOpE0FK5XIlZyNXkCB04skmBMuwk5kEvIOv7+8
bt9p4UCIFwD7d5gNyZLSibpZA/WF5FF6RyXhAh+WmkoPTJKq4Uim+jKS92ZdvmSNwq8aFrJsY1fg
ksHNc0umDIxG7Qc6LNMCpynODWgN8LDXK+f+yUTsZJigiMQzAxuBSlrYM7lcujoGTGq+eOcJdsyr
Q+Dvk2IDheWKHC4wTHmXdHASWongmFy1l6f+hye6dgaDHpsIssI1SSe8ychdD0VB1pmxsTOrEe/D
cOW6aVixrmyHxOdH1DWBb2oZqQ3ypG6cRfHy+pnj7cIoz7nFt2n+mJMQiA8bB6mqmqIKkcYDMGXq
zw6963uRD5LswtK+peZEqGX/U4wDZzPsyxv5xKO1/DSa44bMly++eHgm1dLFYArmKuW5/bAH79R8
4BtamCMDlGBRJjE1ssC0XZ1c2kBwhPenXGjVXJI7ERbhU2bCyLp18Hyq6iXY3GKXDfnj3++9rAdP
bRQDrq4Kgu0MpZRof0xI+yHg2r2LawNbZvZ/Jufo8g3jtwtNrhwegXzDf3g9wQwQPPQUAEpq5lFV
RQsUCvH3AvMrj3rLq3+O75xTQuqoTrDgZxQ2ZhnimcxatFvYGbMdultYQsLOrAjtx612aJCgZfmR
3QcH066uaI//eAti0DvQs2voKdH4rtUhl/IcpwDWUfFbk0GM1aMTOVM5N99G6OdrVNDk4jkdAckL
3IneW1wbaZ49NmbXh5lPjgr38LhOTWFBIWuMx6YsSSlxJDJjHo6UjW8lE95sOqjBuU0g1Qi2LhtD
8mbagPguhBzTi5MeBtZGDC6R+q468Fyji03bQogCGsvuTD2tMpni1MPTZngOQ6BG3gMyu6DAV3OD
LE2ebca6r/jCMh0YToAMkDtND20M/s6EsxFr1ZoPyKoojtJ4AC8VpKARyJvje5W11ZMwGEAdukH0
7Pev1okI2dIqBVr5JCxuKAPBxrAjopOyHZDB2axERe8PirtFp4iJj/TgogG8U7mjpOBZKJad4qmO
IP7dR5I7XPOQpV+fb1U3pn6EC3uuqUgBfZFyYpCCEQ5dW2FkEzTsI1AmcH31hE1LDmdVkKwm1S4l
rqwwvCb59BK7eKg3c3WiKTDCXFTU1phRPWzyMuzl9h27yc99ITwefQd/ZI5r21tE6V03IUgeAVgr
VCWu6v1xK6I4P3alZpAnnRDilMVSE34X7KponPy1qd6yYGRE1GN7hZetL+9okyfcLrPboYxAssYW
h2Od6vfPYJP1IAM15CBUaY63if5bGE0ZHMQzE/0txYbBOrYLyquSBFcBTPiz6sQt/cX7GpiP5fm2
7Wa4xh6fhe67Aq4gGpt1AfwiIKzjhPhbbpUKskAA6h+FAb8/OHfQQaROQ6k29XrCTik5PinQM1wq
fdiEWRT2Mz2att48Kl8e7pfmharxfojaHkNzdK5KBiURi44Qs9Y3W9rrlbmaBRfJtT+BPHqVquDC
j2xPaW1ylgVklyct2fUGMpcCX5Esd3OtFjv5ax5NRHhIfQi7yRHcI+hc1ftjPbLpr5bpjCj6tKU9
/9HONIS+jcdYdb3omaOVoE/WxlhvMxgNH1FJA6+u/Z6ct3h53yxUGAn6/GQoh87rwVHQif1nxy08
jdjda/TesHr8m8UBSwRmMqUvPRI3My1j9MqpGC2m+J51Sg3FcdlzLY7P6MXDehcqiXykpqyGL7GU
KQ==
`pragma protect end_protected
