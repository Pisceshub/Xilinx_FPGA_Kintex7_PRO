`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEOa6Sm2SiU3ShE3uln+ugCMHKaKEmeXw1AArbatnZDHT06dfes0ekJS5
Gy2/u6kY/SFoN9M74zMYSo7t6VvNi2WI9N0F5fWt4b4Cn7cqBo1UwRiYeBukcbkFxIzqNVtlcINg
LjC6sCUiTXJyhJN8ZKmlSxut/gejQWg7FlpvnM9byMGHqQmTwlwvC+8eAgQP5O7oOpZ/STxTxAAg
tkkzoNBOet4ZsuLigA4RXsF6GL4SRAFYAWgyf43WNhI5TEOHxaES9c3S2ozFxd6Y5uRL8WK55I57
LV5/PrfX3xmIb/jgSiJgGlshEoLzg7DCswgILmFZpnLC5wV3Hgc20XSHTNeT7jnVDxoVjCQME9+Y
V1P6zDfZFb0s2TUpo8yRXeE7iDw3bub+wYv5iLV8xFi55SRsnBmKhFFbjUcAwy09m86AzgTSJgpP
lSlqBejKUDOLIbMXuuT+whCqq2Ncg1voCvZgMlgqEClbr81T86KYrhrtf560Tkt49t9uAoo0w//S
Zcq2SUGkRfthUNT7Q7nGrIcCqtMmR8tCeE+3IvXHrQX+i0CJCvbfOc7Z7RjEXUDzXGOco2Lo82aw
0eR5yVSUJ8tnL6rPjfKsDSOnmGkt1OiaLFOKeHzADKZ2BKS/khr1/P4qNUsUXd8bTEDl0pL2EoxA
MG1fB1nFIj9RqpqQYyAEenf3L4UeYuVtrKdz10BXb7IlCmumEzYX8XdEG3xgSE0XHS2/qYFRJXMc
NrNHRAfZ2uHQh/no9Q2pp6yyvQim6YtU2uUWO/31EWkb8QCFG9yxfXvknK5oPJT4DJG7UzI+3Zi/
8ohsU1W7GuzqV4pusGPgcFgvhOZrYWhAHpZlC/7mVuk0Bi8lnNZW0NYpqI5XiJPfz6FHw4Cp8AzB
cLfN7wV7dbh2iro2eI2S/EHRHq9Ogv8tZZWMO0R4pRJA19Egy6XBinqShzNFpvU/gkeAtCqeLFgi
l9S27y/2/52k4Gnr2ffthnhBHWipZqXnnEmkKLKqKZQOAS0jeayog0xCNpskeSeKcbcbpIXhxrGP
Shd768tREAeXLwHVdBTf1lBPNIgLL4wQNO+jAvR2AYl3JGTbHSExjyif8IZdpza+Xr0KuMKqbVk7
sfO+yySLUnl7j/9diUW7fBKai94dgxBjnxphqaR1GnQb3WJv6kM4a2LETmy+TQJhTnGwVwMy4vaa
Jws0NddOXK0VkGSZp1R7J4fawn7u0eUtPNVn+EmMwmqPC18DQoqYZ62VeKqw0le8zOWMm7onMMgS
krPhKYDh8q/8HD4lfghBs52zbuxPXWnZxZqVco99P2nMzd1iAGWvr3EIH4GyQiHl0fePyEbgCB1z
X4Sx0nFD1jBTKxzWthuS9bjLOvNjXe+lh3c6eCu0Ke7fNC2f4VOCTh4A8GQXuA5Cxy2NFc+PreHy
BZdP21pldNrOdt8yodQo3tRk54FNi7ALZCu4R3rIxpPqe36iLDC2IAKlwxmPYZcc1aMNmurOKze5
lvhj09ogIPIRtU3+aFLfJaz/kxQrfQvj7LuROo27Z5vwaHAPkvn26cceOAN2apyjDBUpqKR6EHK8
kUdzbQwRWi56V6wJ/QxVN8dbhg9gQw2Tvu3SJoYe1I9NP0stEvjIc5seIA6x7hGM/ukvRDNUPeRn
Kj6ZElw5Oy/rI330hCFmoZQnEKTLPcIB5XaMwT+rpzsMiRA3QPF7iUv6v4/EnDYuZyzc6RlBpq5z
ILFYoOnhLx4fgoqjuuiYvKJOpIGWkG6YRGtAPtVkJtkK5RF0cnXKc38YLc+VqEe0blWweYpqgwxQ
yn5tY+yYDJIvLFRj/0MfIcORrgNZTG8e7jxEVq99YEvz47jUEjI6Roym/qmJa4XMDMVWAt5vgek/
vSRGfJFm3JV2WdBOGV7jbVP0PwT0I4BSyIkO7xYAZDwiENgJPqYgLoskp8E9AedmdugFHLsd4UHh
P60H57pwJLgd9kMKD8utrV3/dqy+TUrVPYEnb6fAtizsBpvfS7SMZY2kcAoSV1xNCAd8b+k/nd8K
g4+BzDFMMjFv7CE2p5Ce+x4wLxhprozsRhTFVX5WcAyMfCwjxr/a3ODL7UgR
`pragma protect end_protected
