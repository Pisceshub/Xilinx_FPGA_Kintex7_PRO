`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
OYGjrUgyGyjPSvxk0BDAPOf3ruUMkwgusjVTsRN9qseST4k7tSFqdKGk6fL8K3Gk4hv9IOZXVNMY
1p1L1fNriw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tm+rMBIktME8gs5mMkBxD7/nRTfCT92Wdiaw4EuYdiCMUP1q01oLk0s1uSFtD0CuNbK5xIQo5JMF
E0FVaLZcjqCuXXr0YljhZLQhSE3oaeum2eW4FiCLQeJo15t/PbK4gXIGTXNLc+VU+/RoRcftv+Ab
D7/BNM8naSzC2vQJsgE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
syt0OqKWoepxTu4mqmNDW8IgYKQ5tGGtJsGemtK0DKH4ipGLUJwNd1F8WcolX2RFlb/OjHXabGU1
PmfWJw+vu4aNUkFdL3Tf49x7JjEUmn6i2rhq5dHvvDTYdSNp42SX2vwwiJOz99zjchVAtU/Uynd/
1wL10tqaY34j7+K2PRGrvQeoA/fNjnQfoZnwEBIZozsHcJrYLteANZMNBc8OA06stl0HEDt0D5Q9
KwzEltJSNb4fCBp4Eh3paIuopGUI9UOv74IOR89VV+K0W5FkC7a8C44wkv5xgqBKKncqjMNTygte
xWVmzWVVjwZWr3DULVJm3G4zleBEStI4DJrf0g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lVYg2jC/rfuGSHQ3B2wXyheo9r2eE8emNGsZva+ZuwRSnlhk1GtNpqt7QxDBPD1iTlt4cayp+6d8
umBX0Yl+SxAlmmpnDt5GDVCGpOFXUl4hN44du0AfrejtrTUdvn1ZwhcWeRwUggie7mEz5mWel6Iu
zoEAU+h9sWw//anSDt2E8hPzYvAKv5RwuGQRe5aFL38AxEMCWolaViPrgv1pS9rtD+M5E4OyWFYM
Aw2YTY5gwV3aXR7/9v+7s/q/LfHWrO8MkoBADQEgVU5z8hJWiBkoau2zGoobshb02Fh8e8Pnb8uL
1sELBT+K8O5PcSk8rBrGFDtTAO9m3/b7ainU+g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bIhVqHY7XX/9422GMAtp5hmL8V3AbZU8txtMziArtQXImRdh5df70Ask9mhJ5vUCRtYA2gyyvbHz
BEI31PfdEWHB/eNsRSebOEDUNlZrTYimsUJQa+uthgost55lt9sJsL9q0tt0GeGE7kQdQzUnaYQ3
Eu1Do/fkLDMCYgKUr7L4wgQrf9Xl84uTg1RVyy3qCXF3BcBS5WQD5V/T2VqsOexbw9dGk2YQGVPI
oGiKkCZlZDz30uhC42JBiBe49sA3vRYv+nR1U+Obfa58bhWeGQLDNVE8aB3nWGbJIKtJg9U2KVIb
7I2X6dCOXkXUL/xtWvdhiH7SzFqMyQ+sa+dnyw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XQMBqtIU3RLKQTvL4Z8YyqgJ9fCE4u6vK/h8HCodHF3vQceapjD3GXSyzSORcbbLtsgPEVeV7Qj+
iy6sbNdwnkmDk2psNagzyUndpESKtQZ56hNPOGBPs5plpWzqfXgFkmaOFDGba0WnIirRYPXWvs2w
1jACr9H7QhJ1Myul4iA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
i6aj4AtQZlOTKakuKkFoRjWDeJifU0Vt18E4rwVTbRF/Vkkd2YvlJ1IfE0gv7QNk54NUX5Yyt4Nn
7IAASXaIl8LrIK34pHRoneed9qq1qYKdyw6JITLwa+Qe/2b23PAD3dtagneaVcwEV6o6m+MeYroH
2DwK1txCld/WFT6pFaUMZ0zJBeg0KOkHDfqepvbgq2STLB6NtMzF4RbQ6jDvteBTAFJXKSRDP5yk
pL4ZKFrpoOeRl6kWf3wGjyG4ooJhibtARFlt32nlyV30ChfbzGvZv5/sQPIl/kY/8DNRYoaJFOJ8
WpUBESOzd2LYd57EAW/Fr8bdX1D4NkXF6fPk2g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 160960)
`pragma protect data_block
apSnHH7lCVxFNSXYvaA+qLm6gVsw4Lb/VtodeB28LJAKNdlqAfli4DrzDwGVP4tjmB29DfN4QoGd
ncLnllQXogn3COI7CP9QxjV6PYDJQrPWpa41BOMQ/rr/CD5I9ETdCixa4A+SO9Emq2SS3urIge/v
+uNb1B9/PNs4tDsZU98EwvJeXw+vLefr6f1gpw5FNhtJVkKDS1wDElOFsmgTgmKfL74j0fQBgqLl
jR/wLfNvm20ayWCiTiMDKwEai4Ef/8+kNPZ3EK3AEVq/L2sAismf/t0lNt3dHvI7c+15IP4SjfTc
6l50KjU9djOgBhK7lNSZbmMdz4Pxez0W769sS3Xg9twHHglzrZ98tiYr7bcBdaZaQT72Xby07jfq
alGXYYc+8pqnlGaT6e+oe3q+tgI1ZCz+5fzogp9M25S3X1BfpddFV/11pVIceTGCmsl/DB2EnCid
pEiVpJoO/DD/sscm2jCr8dS+goCyBR3b5yk5+EpwOiSyRBhWqnorFlIQ1N+LmU4sFWLCE4nSnkeK
y1SU43lU5dSUhCxhA4c6tacHp3MBSuS6zUTh0eKF/V48aUrhaezmQt+5/IvTkPe328RFSLoLCFQj
ngifgu+D//Z7ee6GyAFUbjNUipmfNhJ65yu45a2SLlXWC3JOYpkpTJxwFOXUhX3Lg0HXMOAFk4Qi
DfGCBAK0f7d8NehpGcTMOkilcQ3u2KsN4QtC6WsfRnfWRZeGkfLjH+CD1hHGMoiuS/8NxnaCKPpZ
boz0/r+6UXNFbXxQioW2Sz9x3lv6NfZQf/wDdgDnNmJ5L0DvFJ7evZdAQmhfBTATNSUYDRhfQE43
QMTCgkcn/I2WgHJz9uueSWTA4a85Er5ohDG8Uazw/qp1EvmRkcBGdP6lbOJTDSmq53p5kro0JJ5R
s+ij81OfBgah80DCi9FqxXgfVkRyyhDMrfA4X1fq03vU+nvwDC3MaZ0jJEY0XVLRVofk5qQ+AYi/
X7OwdLqHfBUywT+Ca14C/2FvBj4sSDSbEOG0jjyKqUiWOoQSNXFn/q6YHK04bPpU8RcJXz0WaTbp
fOQH8xGEHx4D1G8FdEb4q5aSEeRBkKpG++BiEpjffdOsteY2TSwpppwsa34JrV3gEUNWJFR6LBBs
eSQU/8KvAc6DThtIBrH46sd5jxBUnj/s1osYizvsR+6RgDiD8uUgiJijVpEgyw0HFy20O8LLbb5m
f1iMTksvzfLQwBaiY811KT+QTJLTV5p79Bvu4Mwozpjrq2jil1krNxu2YUDa8FAWa7GLYaJgZNep
Nlm1AhSKFCeC/23Ei/BIp2BSSSk784LTa/UtcygmxzrGGBlX/GyEyjEKflNBjfV67do4jNYqC7mx
OTaNY1c2fFIRgOah1VAVLj5JkIYyfLy64hFnZLSwgCpIKybO/PdxrzJciufTbfYQZSfoxLWjPBuK
wpNHbEvLSYX4fybv8iGbhec3HhWT2Sj+OvTKNMQ9KkGkqPMNrjKtuk7dXRY9RziuHbUm6AtAua6A
et7qYp35BdZ1P7PJuYGaDZ10+3oceQYEepq0DNBpbNFecQa4etTu4SRPxPNgPmzJb4ayKNsApSf/
LiW003YmupEV10JqsAF8cZbp3NOcpjcn457TvWHHNrFF5PE5E2LhHqEMPsEdoedf4dFSVPq/KicH
Uzg4+Jea3MoZZ3xhDJWGxMKNdR00I2NOTuM4EPXXecd54GeOHePzX17e++8oexD29K3l0gEbg76Q
xHGhgQGoqD/JJdSDjPY8fMI+HBQV6F5W1p/kfNPr9Moooh8RJmH+ztLIXCUZKDVlLJr9LTbmp+b3
Lc7jPxWuMGLd3VL2uDLVu9x9+/H6N3tvXeygLPs97yyCjx5ObqCEDp6C3p9Ju6XVXre/g46xqNKn
sbw0YGxcWCwmiRNzcLsEJ/wFL8sWmtUroT9AdiM48d/EWL9VxED4RPOtkia9XicRUPM/81PizS6n
EmhQXHgbtG5eazXDItL1vxlhrgKvQ/p0AQp1U0N3hIG0vjJeUOmwUyNBIXbKpb2TE//w2Yk6qA67
7M6iu9uVfzIOjXqqtP3lN7A8w6EFiv9sU8q0zQ5eo8YaB3Iqs4etWe7AyjkxX1bg0pppYlc/PSCf
EFBmdwUgGwPPerRYjz12NHsUsmQhQ728MrFiI2/WZ6BndBr6ewYBdOEhfUk3D39/aDo/MJjrlBt1
XZ++U6UXR/fqwTvBlpsZSYiUuOJ3Jt8bmJX86RY1Ad5/vwXCUWfxBopSLwGghu2KXrAJZgWztGgd
O4CQ6NBuCV0TFGBuYfX9vxU+bNhyLowSkRDyCeeeI03FAzydUM5SAEvaPNrcL4d4jMe3XkxuaKs6
0aSKkxNWhdHgcDOWJY63Q2wQncSAa89Su1LEWMp3pqtESMPTqzhEI5yhMh5ZBNszDYvKAgSTTvYL
9At2b+bTTpE6A3AM/xb1rJqDwt1WdlhOdkX+ciSq9TCtbB0hKZwpCZ8j3UykG+LHKYH51mLX+CxX
SAVr6/iXvRHBQ0s9OP/M/e7hAxBLWMw3pVnq4AOTvMT9LX6Zx7iIfZ2cuNyVtN+WqCAhjFD70HTd
VypYBjmQyV2hmncNvYoUyL7rIEdVau2+DxTEIvubMIORCUxFhvcuFwEaBXggeqxpVERcyd+heKbQ
mRkF50oY7/Y3pBSw1O84CMb/H9TpRWUoI2BAPcRLdQjtGD6DNiNHgsn8eyXoVb4f0c+DEYSko7xC
lRmbMsnqG9BjQkFUZZza4+tBC/kNB33EzV9/RJ5mbDorXxIsvaJ1JxmS5q+8Hd8ESpXIL5QHoHem
I6G8eZEhvLGYKxtyISUlVddJEImkIauLgA1FwlGJpp35Kwc+UUHgMMhYha004YNUE3K1g1+qL8aW
7d6zY49HgAFJYKFNDzBU0os6Ucu//ZCvm8359t9oB41lOFsBmRd1ulSLnlHVZYLsZMuO40g9qzzP
eqFG9iPLo4uc2tIES7pbi0Y+lJctkdYDnQLHWNB6WsOZT+/2ZCU4M3TI9usAd4vcWBFSm2n57rFt
EFTA56BOBXDxYqis1JzUHhbFdBZOLNWzDd3uO/6ksNkomSfVBhmuthmOd1NDuz/XmvxlKzP+0lBc
2tsWnM+6SyGyN0Mjx9v8L+PPDIlvN8DX1RURPqCqHxvpWQN/Exqw00RxYMMLtNAUk7spnQE032QQ
BTw1Cn4K/EMyJqbE7ifVDXQf6/vb0i+7ZrDeZtJmTvlL/v1TNKWSVK6Gi89IcQW9O2wIiD1AYFbR
z75GFm+6CVDuyYoCLFsd2gBVcFwsK4GcMlzy42hq+xzXPBR2IHh19Gfi5EvrkADVOW6HLWfJdSBs
9uHA5ei84Mu3tF9LLj11ZBuzmzI8OzTZM4S2iPN3N/z+YKNQgHwFnF9zMnhwahe+Hjo6+cpi+xjl
WgSBf0gRrRsHTExXnkxiJKgnb6wwVhau38UL3/6qUx3K0zwUM73NAIspmTiZFdF6ct3jdz59zsne
5cb8KRTAIYkgdC5CwaZfqfQRMa1+5oLIyH92gz2Rfs/68Olc4Tgmow3W8DG4yOr9KwqfiYFHcnyw
20J1a2t2fvDQiHFK7gfo5FvqKfcanfnTts3i1OkfOrJ8BSBfFSo7yKksFNTS4CbhfLl/HEhNM6Cr
VXLK7+vbP03DAL3M8HuMaVdJth8EWF3niDzu/3g77xjIplXYZhWDaEFxvDYyl4uIpTzkNIGqknkK
GcS8e7kfYKbDI8c+zH0Ihy2TRO4MLK+O3beaevpXMpIVnpoNQ3oCPY7DkM5GK+twL0C/B0myG0dP
GskKgEZoAbp/Rwk3dYLKS/Njg/KtJyRuOzceUNBUwB5WDoGRGYSUHgfp7uDTZxkZIMshtY6sf5x+
ORvHv3Z8wfvbvIy5SI5qtPO7iaBZ/U+hpw4hBKSlXrv1zMbmMeznjIfVXe+Ll0LTxoDTAP4hcS88
wIwoNeaON6/nBiFfUcx71pBTSFUmpkv8yWKCBLjZgdRl1epS3Y9q1gIZ5bxbgOZjUgEsw1bbKKJU
79XsDdXoENBYeh83R6Bg39/vGIUaKXD6Vtdcw9RqP1d3ju/5lCKtfB+48bcB3vPuo69M8bNYGOUT
U5NeOZ+/hQSliw4oyBsP2SpjMnndyojRRqYvoJz5p1HXaWjwW9ZYgte8+ddKJ/I5lH4H8bE9pK5d
RLYhZK3oXFxvDf4a9LCkEu6wdXihmgeKeDmnUi3Q8+kR3YitYQEnEtxVfAVGYcKCKMpGL8So5d79
4pXCKhZcp+IxHQ7O6eW1clFx3kCP1nuc/H0eOzF5ROl4k2HLKH190NG3N65k/zqxGdlM78FBosjH
NraJfKpMj9n9NCRe5WVWUowM+PCMeAi9aekNZdp0/UdeaNLbZAyS94lrbFrfPSmkpuuGli+3eKsJ
FnTjSDdx2nTMrQ5uhc6UgkcE33v4JLseX2TCA5W3kg6dz01vhVP8XEeUgiyIoxHq/yfoUk8Il5gu
r6C3ouV0SZWPdc6ylAbSfcEaLqklI4qFa3+lkDDjuclfKfDfooOCDnS+qgA2etBd5y8rZIFUveyl
sg8t7wJlRsNs4Z3CF8fsqoAFLQ3Z8Hj3z8J7ry7V/OjzrH1q5sWsei9/wBz8w8QD/KiTo3xp/g8N
5TgJqI9jMip7gg3jVDJlmTlBrSeECrQTdpqXPmjvRGaJBuF0pEUivYksAVvSdxOeDZ+Mg0jwD9DQ
jh98ZsH6sXzX3uZaDyRqGCcDi5T6cx+T9Mk8ca7srYTWHI2FSxLfR2ltQ3o92QMEsfxEtzIPn097
9vL4e+K89AU7SptjgcBQchZDklQ8H6vovr0zi4cQvwop9Wgl4UTuFPf2AkqpG6X8WmL0l5+s0v9U
Gu/OwaFUe3gGf+qv9jc1N4S2XTesZUWBUdZqa9Mgxx7IwntikqAY595hvxj/caj81/bRlvyDCuuk
v+IapypjnlK25bryZ+DHk00sOUzZXVXKm4K8YSZcCf9Yr6iIhDzV2cB8gbLXhxP4EBU6TjC5sqqY
EInHcQRVijNny4u4wCm5rdpzsgnSiN1/F9UY7joqbkQcanIZOWoWcVyaEzGKI9hIaG/YorX8ZJ2C
B/j/T17I1uY375wa71iLNHYgDyASFsYAKpvtNCH/sIJq9Eq6SI/62gaEyMiHzDbBL14bPdLUWdxm
T8IUlUp1kxgkwDDoU3zPhFD/8wUpfVSzzCYEQayfJJZHw9q8fqtNzhFJjrGp/YfBZLlbK8PAePR2
ckl/cORco4zLmUqTmomz1/BOI7tuZ6cf4fe4GnSwUdAMn1w5e50fE6K4N70jjj8B/bN476iowAXp
HM6IdDfvwhR2pcaF2IZOT/Roihn7wz7emSsX7vKKRcbm9HOGp2lhVXskd1g6idjaJEAZpwZQ1mox
5L9hdB9BwLumdOJIEeNU+/L0PuirwGbDQdUzyrEqA2r3CHB+WEdWQiEFuv+mYxzWhsvyMRUUQm7j
XjMbXhbR0mlExRuTwu1cVV2O853DNIxtiMfFTBnm3qoKtqMnPRgOrHNiqMobN9Ru+AaiSV32JJnh
P0rMyLsLgHvajwrVrK+mg6gtOVWoY32K/atJyiX4n3r+totBk4nE2EtdMRCJrgtUH4tyS+73hTpa
iZTUXRYpR6XMD0npmHif8vt6RpEAvtSVwCIEiL9lCOC9VnKc9D9CV8qsMUgWoJ2l7Kg+BhV8b4Uo
gDdYGorYl9UMrYQsoUHhpzu8SREEjK+LsiKMzQWHdcZBmEdKsH6EJluerxXk+Zip91xKrJQe8uEb
BWqmSKqk7eSEL7s2w1B6VvJWrYHylsuYq3YpR+Ex/1BBYImUdIrB4Qn4AMMtumlBqqOK4rcuBMj3
az5f8DuJPLpcTLjjo2gmVXTEu+xqqODg92iD+YgSDXq3Md0Ev7GxjuFnCLSGbe8EAWF9bS6V4WOj
41vKjcwewXQ/fwQWfpELERhStWEFrzcqt5HaHKQutFPm6/AWbA44vJluahmRvbRQpG3RxY5h0xSR
UJPLRdTSDtnDSeiq5MFU9uaNhl229qOf5eHgzv0jrH/KaVgQa1uhchgx2aLFciaDSwiUNuc+WYIV
kgPMrJs/8Uw3206gI0r0kTM/GRX4cQPMJrTQl2SIDIhY0UBIXVCbr2rjh5AAhQ6U07isGlTb1fOT
aM/NOQ73TN0DMPqtJGGztglCPPdaDawPIB/gHrsYg/yb7SPJxNVr0O4mPQ2VKHksf0dFHUptcvFp
4q4GpS2n9L+4TefDwoMgobB1BGeq0hIw64iYV+XjbdOPIC9wj55mDkmYZhC3H6ZKP8qIIt0Xm8GM
wihr7IVhALAy4+EV3z18Ap4HOSeLnmHEQb+SIYGrcUzY7f58FDXbL/fTzsTc8f7arFdtsM1rknOv
xa/1AxmjDv650ulQQGjO0fMgXWtqckGaV5s6sMS6TFUXUJauBhMHg9P96R0VrhH9/lcVyrODXfKH
X4aBYTg+W6azoVwfT183ObmjwIchgAGRH8DXjW0kU+tFoZUWft3fBSUJt8Y6DJPOc4rSQaixsfWx
DOyE01r2FGhCDF+9hhy/0XiWzl7CtR8TowtSy67uDTBVmeZS2sd+p7ItKc1/vcNM6iH8vm561UVX
1ydIIf2kgS8hc7unkWD25VsZZ8WPrCFwKV/6dl34X08MJfJg0eBUXESTt6adjP69F7aMegMx6Z0I
feRvxUVT7JcFL1hiLD+M82448dB8+DkgL8enaP3CaxmbxNTEFAG96dTjc6KYC+ws5eToc8VRii1b
me0offoqnal80LQ01pfSIGJcUOtZ5UilGlSzAiHVWhbkOE0/w+hKEimBWJoXlY4cdNdrQ+sN7hQH
37qv3i1IPgyjDjw2Nvafi0Z3fwJW1JbfJZqOxbrMKCx5+ObVGeoJBYx7H4qUu5mfBsOnmfTMlj1D
Sin1u0OqJ3XupDWH4xRdTC2rWUBprdBnJSp25UezguUzS2KCIdCpInFPbP+6Yo8rhFvdgrFUW0+7
G7GCm+UtfaL07atDISTHRt+v8YIXjHfsS2+ajcv5TSha+Q3mnr/HLQJi9Z8I8xBmoDMpS8fyjkMw
qg3R1p04WN+zWs1wZJhA4x71ZsjEYBaTnCJVN8hmMtQ602jH7hgSCmhXMTiyfoDxTHQwWd1X6Qmi
sQ3nQrf+5U9I2tDbwZicuEqoEgwhUxjd0s8IsnUR3hqHej4xtE1P6h1E3hTN4Lh7T7cG73oL5Yhm
kjHmvs51rJcAgzuDFQsq90P9UmaC20cRUfM8ZPRfzZ6q2AcdqGWOOamO3M+2A5/lijNK+smH5yYt
sBXxtQtxLR11+rwKjH3TE5ZZxsftj54t0sol0HffhtKbn5NxICDIr8FUJN40zAHF4RIFcLrPnL41
JUBXUOOW6trIVCXPd670h27mTiQYUn2EJDos9ny6nIrkf6VxnXfLEXsLbEkp3sOnq6AvwZPfRhua
Mhw+AA9GCRjsjqSnDQ+PpNivez93k1FnWXn5em3prxXsrY/2sefKQCcDaTpp1Xt36jYPXJyaXoR/
S9HnufOvFH/aTaBz11agRd6zg+E5swZJjpwjU89DhobzhYBBdDSogKOOoqtl1NnnYIBKybfale+m
77d8KQeB/lMFGJjYGg7FL+und/ywIfbawgPpOpdYhtngks/47LO7ir02kQb58TcEoRhNls51A8u/
gE8wcGIRADGzc5rrbwgXIIK8sAWm/eCh8CZ36MOk5ZnGumcCeSmGf9HIxxULWW7QB3k3ShtqdgyN
Glkh273Ka9MmK/pcEVJGZnoCDcVnAkSdlerrPJ2jleCHPyqoI04oyHLoW1u2VaYKnuqvqX2VAaIx
bA4kGHy18j6y3n9WBjrZ1hinxaLHEl2OLjp5qYmO/EDVcash8Me2jDK+bRUW+zzDmvSFUH6Nlg1A
/4ZBep/zwZiA/FHtkLDe0MCdi51ydzzfZaWwfcvUX+We85NKR1oqb8E/P2yd6a1WhcMAhCGFvkQc
cm9Fq7KnX6/wSkCxNoBf7d6aMoEfYrXl91SisMqNFAqf3yWUrmchngDv/1PfIcEXgJn8i3wZvRw8
jfxZmHtOaFYT+RBTIQln/pNSKFzM3xtKWt12GTfQEBe+Iqenc/1L7OAWybMWUQov4RkI7ZOPr1TW
5Zra+MhWqymIo4eNI2DVd+k9cEOm/WAPnZi6CUkQwVyIy4gzxEKQg0o8UBVlCMXPgrt4ZPJ+n29I
rQidQhBTxwEBZEtpvz72/59ywdgAFRQlkaPTEqhhayfdaXkP56GcYGVfikOZDl8MXt53AZ0dlb3z
qeJltgDL+2EOsAkV5mbKLsJ8LabBHHdujEQWgeLOTHGxtea51K6MggJdp3M1U2egn1ciO0FAJyFf
007fpT/u7LyZGoIXzB15Ckz3V8uxjEkFflJQ1q3t29RjXkPTqU/dw73CCshRgWYvrXYzOBT6ruQR
IrNGIcOdhzdSFKDjxfUcyt07JH9uVh5wX3wpb0Dj/DdYURTtIOaBM2cRvfxiegVOw/ly6PM7d8BE
w+eO4BMU2oLjiO/f+JG0u7IU8cL2S544oCMof5kkBGkY8cMPcQMj30nZTD0xlpSQjK5nkjqZ3csO
feS2l/mWL+vElHLjbDcjnJwSNGppE9YRoaB+g5IOGSPm+QpO+VCXLqOM9eBjUfgFE7bAhRSc/WWn
3E6rtzUm08a9gsOO5FpBnQHG4l+mujRZTXbE8wjsdCIQyvLX6h28CfZ9aTfr++uhI9qNSxkNPwdA
Tv0MJ3/kJpR7IDsu7yDaqZDNb+LSXzcS5CWldHuHtDdfLWuRyRio+WPXtMenyTHZ8fy0fmctXvvK
M3gbflVV5j+6AtKO/0+LrKO6Dnm5qCWXkuGR7GFkcAyjFb5QhDa2So81UzJ2aZuw9AyyjS42LBeF
YPx37yTxtLkRKffEw57hyg4EuLebgjIkBIazJSCicHYFhvb3h/zCcGVgRZgi128uKh+RJUx5loe/
w+KEMagNwEgVzUTbK56pwGL/5funtfsvE5Yua0jX4cvzQv8Z9Q1J6qQ3wNlqIRRavrgXdV41qEp0
WLU7XRs2XhtuKCJE5bMBTv2mGyOnCyWS71j9IXK6cQlKBhhDcGUIYQSlq6Wbye0pCB6o56ny9NaE
uWdNk7zxcI0VL6rXRsWTHzWGpVQxC3q4IdJS+5Uj0bhaUjIolfrKEY7cv2jafkHLbSLlGwdSeDCp
9drucEfvQt6l+BPnSKjJymiRKFJUzBc8AYVRT/RsoOYPPDkT57tbhHXH7vaEw8ocOPJn8mla7Zy+
S+XRm1FhKyB/Dhm6P1HJSCTNjCLMbPivCRRHergkRsZgwME74grQvopqHk573Mw3e0NDrcmSgPZ3
E71gsVvt2SUlVmNub2+BFqfxUFiLiYwC3wO/tB0GLMJPstITf3XVKcX67xu+6lhp5EeM39gkOSu/
jJ8oU5Wi6cPRiPj2+JlGkqx+gB7aTHfWK/HGGpx+OFmx48jjqXCmQaWnwVvdvF5M459gaYRXl0U3
QcyBzgf3Q+Yfbz+ex1co2WK1M3bkTlVG24Vs6aWhlIeBlNwcq9v6Jm1y3hOxVbArOp2/AZf8YPoO
aQxENComRkgPR1Frl/+vkJ++f2V9jL14PyDD9Bhbqi9JsEgePZqdSC930/Wzx1g03k7/mheZ+nUg
UxkaYFoLFTeac0GRGNNEMSHm5RZQlFL+AzrBHrMCGQxD7QLj+VEbx8YptN9n52wWUf6OhjUStUbi
DKly4O5ItG8ASDpzPmOK23P1vBgYFtNvdQhFjKwbR/Y/nZy4Y13UtoNEXh6JsFIfnmPrb7bE6SS0
vJgSmMLGQsg3DTy+b3t5iizk7T2B5w1NTDP29BwX+Dld7GG4hsC4K/le1tbayymyg1YmmtP+lMaS
86MvCo8Xb3p8JqxWqB39hHK+FyD+SHVhxs+nlagp3TKEug2msZTU9ByEnVguoaPU5TjjOayg8VQp
FZPUz/rlGlTMjizR1S8NIG3H8lf5cMi/HXELaYiwIv86AteCMOcVfgAuWyMCXOOSqbio7BzgDTod
jM81H4oX7fxIPi+NwT3aUE9ev7euiSaCpmccx6FbZsoQzqL0Wv7t8mO0Z8ZoAPnbdOdPdzeA+HNA
uZBMmzM+1QM7v9Xj8ETOcvtDhbTwS2OiOuwWGBYwrH/30ISC86UwQSZcrZRw15z7hr2e3LEECnTY
MkFBs4Pw2FJ336YkKPPqExUNEd0TSI8NHBE+DeisEK0sNXP8hVtXhaGYXyISX6rxl2rhdS7WZlFO
tJRD1WLUYizm1GnY7nGX7us7dSRBPNOD6689DoS1aOo+lDUE1JGAJEC76LD9414HdivC5/GF9ZRl
OMdrI8JSfXPdgwiSPGdYM7RLLuKoH8HhM/rQLBXu9RtqCMd5TgQEUMg8jhsKw37vo1n9XHT+9P0w
6FHsPLxpw2z8BSupuYGbtCLKQIJ2O9WWhs92b0pcp0RdCzaYEuh3YapRwGWq2aCxsB5AF79Htq8h
gB2JkINY7x7TuI1WfCPzOFvPJj+9LojiEz6DzJwQpbwXZuo9emXTMcHKObqi0asNPj2Xw3AunEwe
ZuAZj3SaS6Ud8vvikPzqpEfK9DW+gmh8pECeDxr0SnVK8sK/eyelFEXQcfCe2U9Yfy+lpdVURuBI
It4/O6GbFdvNLBdwLnlVcQjw/SEpjF3Fn3whf2ubi2CyoDYug2E5u0AiNgOgNs8Xymw79Ho2VPrv
wpEiejWvKQcNdzWCAanGpx2GfNA1BgMT4cbwDTgTzSWBaDIuc6hLV8ylAj78gNM8Th7nZ0/sOgwO
T3IbYH32rMAgvTJkEMe+whLSAwHanLDjRpa5p1fc5Dzui7XPfX4YCOLytoJnUS1IDf7isbwC0Efx
Py26Gc1WQ38CZDELiq9xTKHBs6YaptHWMa9ZdCJfb2Ese4ou//UGveK4TiiDRSBopQFM4wg/k3cU
xqNHk77cocRmCr9bp9J/1ZlUANGR53S+bPyQ/lND1ZxCRLOH8W4yY+Y0EWNUlnZUmH3ciJSjFZO6
D2QqgfNxYlUcQ9CBXCl+DhHx5GHk3oIBey4hO2xufb0mDRPUR+cKDR8qdCsv0B91763TyIWzgrl/
h2Djhhy0JlgCj5TVUyuGgwhSUcaGTv2dVI9pgYB+4Kf/ZPLV4zzQE2NIEuLEAMjtmMpCMtpCzluD
CKX+KjtPzpOEYT4R2Zm2Qt51alcuEqnJ9OiBreJBm7uq+agS5aCjttn4tdNVoY/NpyIuNE0Tb6D5
+omnt8g1xhwnT2t1UfKhjJ4j+WcrLJP8nxyW0FtLxUGxEQEq15xOrZVKdiJvtixW9nG1vtG9jvhM
amdJGobDgnoN9PdfkPNys7eVyrOJmgM0gxyF02oSSyHylTx0EtDF/N3pxChiNPJyU3lmgIjWpNKU
QdM9grlm3EPaxCRBgsa8YeSxhkBiId/+KYBAAJ06DUTcEbTG+VD0ww0p3PI7DVG56HOwa933jDRO
Wh9d7ZIdL3bvGeXU4VV5h3hAv4xlDwOCbcoI9RWhAn4jiMsq5ZX7N1nFIYKL4DjHqkCMxQ/qJXBb
2ijVif8kIiJO5IzCd26NrD5zGrwcghgUHqTxZL07aOofemaLpjgeCCekVbrJ1KZ0Ya0KRqYw+29d
NFPJx9DC9CB3K6mMx9i3cxVMQ7xcB+iOKhL5KJ4FZ/pc6Zyc7G9ArWaPvfj4RxbagVKgKmAmjNBF
716TamR+sG9a4RDeAzUpQ8L6L14BCsaw5QMizL40rZecQ/cS+kLF0NqcLV3/WRosejdUDnwm+7i5
WI8+cSBbXO0F9SC7w/K95po2lJnuvy9Z/BZrJuLlEGQ1CH3u0jcWshheTPt2SYUZ94vGyY/0BFEw
F6PL2mDuNDOE3dJEyEjYsX7MjQBoR3MESZCbohhEcBvyJVlcJB9cZTzenfh82o2f0hxBfJEO4Ink
f7GaJT8XtCU9mJ1ABvPJLo5TewXWhORy8dEx5zsTTTJ2nnYDKPWzj0qE0jAPeG701GIVq5S4qMPb
+7wKKlqqIiDO0+nOyHtiS230aVPQa8Nj3T2e8rqErBiZsVFJbLh8PP2YLQKLvYr/grOZIwIm4QYc
BJSoqjme7KNNsYfFFBuOmjgBzqCawllu7RIKVDWHZ9oUraqTU2piZmbgwYYsFI6Xt/dcj4PboL/r
fbiId3APk/YlFlKUvwkO2Y+sW7Yk+iU5ICZHIzCZrtPtseFufqDPo4y5duJPHtYopPjVl8Ny7jBF
yZ3Pv1M35ZYWn/LUENyYm37+98Xiuz3m6+FzX0Wbd/e0ahG7AQB/Fx5ri8sH6PqmEgZuaHj8TTVu
49mVKWZv6bZYv5z12sMaO4/rO9Ie8c08i61a+2AUb+OBEhr1H8KkUBih1ya8FLAm025jCOmqY4Vy
fXXLlSVgBj20zu4MUcjtFHRuQGtu2IIpVL4qNoE+ogHHcZql4DAPCIUPE9hoHWds2DU5LwYjaDwQ
7PA5SKbI3GZ7s+qjihm3lpbZIURRsdxNfhsoImoh58ZHMGrcdKdcw8NTXsQPYNG23TUItMb39tee
PYAmpvHRWGqjALdAbANrJvfCzDCBGJxObwlKNkAyKeVIZAV6OUAqH+m6dA9dprv4O8BiZgUa5OJh
s56JB6Jd7TfaSDiFOdoIRaF0LcqYmPXm38en+Aa2HenNOHmoUJWEyVgbnpGIJQYjM9FYkmy/P1dk
5hVSzEjb0CxNW9hL/kNq9FmbMi7DadFTDcsDeqfBYI2lHn39F+ch6DZ5bg5Qm/vaSiPJpi9lScWs
8RXN4Wr2JbOF96908XlcfrhgLYTr8H05alaRYI2neBuyd3z13bSAHfSkZaW9FfqNaoXkQmnQG10x
MZVS+84XVVqwtJ5Xgyy8AdddtRKVT8GqvOQmjB/fLHxMzVnZ/AKHLMPGMYptRGTAUHyqZU3xrVHt
a2c9SSD49aOqa44nz4avyzJfGyHK57KBGBdbjJNcKFv3/PLQW05IBFzr/mVBDzzD25EFeFqMyeBH
DrykB6ZL9J/hXTAYQ2K2WkL1Dzxf7G7/J8vLHMC+lYkuQ0KkOav7MPFOft+xG8jODLxIyelmKvEa
zerF6hY7xzfKxdG1c7l9vy7Q2E7taJor1qt6V+Mzq89YIJRUqFV5ZfALZtxa1qWSQAfebovIavrk
cERfXP1BKQAvfE4e3IGH7kOBYQiUme9Xwp/XYGs/Msl+FjMpFUgK+rfx/FQBacTu3pzbESG5SHOq
XOJqRqIIFtytt1EgCwTsrROhUjzKsjUZCyT6OwuukQxK7sOpM05zqulOaKa1gh7l/tnPvyHwA9XN
gFqHVeRVzkh78uNLkDt/so0uTWOruAUgWfl7fWA2s6YLyFK4vmnB4j0NxMINcWeKpIpqCBdJY5RG
0YqmZo7eZU7ihGx9y+Pvvet3I+rZDvT/K8NJ6V11ep9pHe1rxSKsII9JBteM/d8O86Gw++L4ID1p
bNP0y5ilJAQ1xpYXJ5NOSFKwZp3d3JTm0hYjU8YAJiuX3Jyxhw4TP8/nD4KwzG9jDyS4HndDQXsK
t7kG6w5csECUvtSijU+8dEhXdCHPa97qc0PBAVea5CmZK/+MfT3F/xyoUJdXHedT6+qzjP85qo8g
Y0gf21IISfqu6DUIuwCXhHECZbNBVg/n27NI4hYImISqa32gPUH7tHI5XTpUiiuIF3+Qg1Hp/tyz
i8ZTMK+IHNUBLyDX8+S9meki5/tGmuP/GXuurBBCHO93+oQYj0GIbCHW10t3miFa7+YwtDklJFNF
+dh/Ghzyyk54YETx9oRHYxaE8Ntu2sWYGIvuR/HvNs1T0+gZs0x8DTtb045YtaIj/cWzxUEyf5Au
7Nlxp9wrKh3Cg1UXziayNCrEShyOFotSOxX2ykl2GKpHQyj/vJGgWrahSLfuhgZDZJGwvirQumph
SEZvt/42RLPXLgbq2jtWtEmX+NweSLywnwvax/8YNT44i2nhCNIUgjFiUhVChbRk3U3gLCXfGMs/
9iVGH0lz6AZ8bOrYEcnyunUSQjv60DYjqeZivEEhbwNflqm+SKPcLyuzkh70Ls9ZIf0LOTYr3Kl8
Y+Y1dyYKrTg/R+MRDd2hvVBMEX7LtBB3PADuOh1R7j9tqQgd8DVJ+mpR/ooYBcE1+s8Wql0Sb+/M
iAp12BQe28YCh1xji6eCEFbhYjs/P9skvnBf4kKPDeqoXsgFGh32y19u4JuyUU5WmgbQaCH3qpYr
Jq15sCFoNHaleqHjnBGhxMC7O57m/MYNVPW8ALel/jn1vUF2BvOrk0td+HVWqFIHh0kHUyDyplL9
ZpSQf2uoqoeTbqkgdO8A6FAv1EaiNLS2pj8Nx609flIJU7RuLEbD8wqY3nNS0sBH3h+WWzdKUszc
WRL1GEruTwwl0hyaWmpK20ZqyWwOG3SkqNaUiUdskIqn0k1URLQYG07+FIZeZSeTzlELKE+9z4mh
DTgu5HsKXbXRzAHJxBz0r2Re2XlFrZxMpZHUZdr1IUobb+KcSWShQKeNQWwNVe0w3wVyO43H2moH
Khbmo6PMq5zLJ7+1v48GU0o/cIayUVK/lFsK/YghUUXg1vo7wC84+WbxAFvN5wjMhEZinCxjjOQG
Raze132vnvyUGl8UOFxknIkQpIOPRoBMeihMcydGWd1nnqfp2rrqtBcOqwjAs5jRMRkpNXLcyDQy
FnNJCXnfEgRvm4Ip4UxT2AZwVjBNEMCbO8g6PR/AzroFWbkT70lG/cD06+VGtcX23sIOzxFqd6Gk
RHds3LKgUVw3+JAgPHHjZd5/4hBYCkZlJ/AWsUmbxBPdT7HOvSN6M/LW0QW3+MG2VUf84ASjdxNj
YhV/nhZO91/CbTqcTWBOu8EbB5HQ9qel13bGkJtfi33HIKTcLQkHh5WoZ/P3brl2xdgpbMWeWAxn
szxJxnKAY3/GNPTPwwo6ZJAMmwMm825Oe8fSJZTeJSgoF5fUx9f47EBomuRiAaBsswVcA5mURHrp
tNxYxSXfTgo8a6nzd42zZNupxTNoMKcYHvbm/6b/hFmpqmz9gc4BYF8JwrJVWvpBaG45u2nn6YGV
kh/4yX/ZeiRRL3a7d5/T2XwmMPMGzo3kKNqjLeoWr0J+U6EuxxkOtVB9owlI+nhh4tnOPQUYP0p4
FbOE0JMYo7VRdUr0q9H+wy2K48v6aWwMKJHzPCXHTiYLaHVSul2uXamD2E/KaGvvXs20n7InWcuz
mi7e+Gx+Z7OY38nXibHdTfDFLoy67X0p0CxGZ08+Cid4sZNV/PsSnC6X2XGmcERpqzZ6EqdCPN2m
oTIleKaHHg8B9wuu3W7Ayxzw3m+sYJq0htKVjqEiORz/TskpIba8BwOyI8asTx7PCzzVVftkLTqG
gKK3NpgN+9Zq9RQ6gnrh1pw+3yhFsXCVhpgFwweYHLSUkrhtNIaxqv/G115UNgBQWcdZf4tkuCQ0
8wDxwZ1Ue89vuxoSAz/whZF7UnD1rJRYOJHqfagm5uYVbyvNxFl1UWeIpqj8cHxV0/FM2OC/KQWK
yNBK2+HfQt0bUb59uVXhT3s6/rdoxZSeqT2whINMK7BaOnGgWJJCbi0rRj0ke/oyXN9BFijO0Gxq
dRjv4pvNGE78GSyO0jW7/2ukcFy+W4mOXzk2/dTugmLkXgRikRuQFswLmhr2HW5k0/puyiiglqlg
AKLGTQgV+cj4kEeoVzLNhsRikhTskiauiGEMntn7SPKZW51oN2Q36kSULe95r2Zd4Lc8V7H2Am1k
14Yuhq9b728PDewSyiXQyEvwCfn3WESgOyZoDXWJuNLkwt0XVF/dtyXvV+y9MJtENivwmFaO3uut
NjVnlvKH8ZyUlBmfibhceSMID8IqNhdByNB1exrXM97mZfUoSSAbvV84t3V96yy7ZaVcNEOz+jO/
Lq/qusxtlHC1l7pmoYfLaujjHUhOcAhf6B0GiyNa6G7Q8+WdDWsSpEztejnoh7oPoGskANPRmRhU
pK/5C3lbeV6EjYfjo6m7Dxr+ybWZSJXFmGXaTIOtr/Ux0Fs9t+qlmovyQT9hnUImb2ASgqpucODT
YnyEo87NdyOv9I5jkU2qyHgzxcdS+bhdsgRVbhBiv4RIhK0KyyHfGtW4iGcGOCVu/IH/fvj+U9tw
b0huOKMQn0hqWanPupjcI0/RLIiafOiMhQ4REV3jrcUMs9h81AC7CwrIZAR4Jjm6tcIEEzaGNOqI
RvMqaM8N+W34RSk1A+zPRexZAlAFpguAAdldcyJCl75YO7tRqt0iGOuMEwWCyHYNMchP4ZPAMoSx
7xiiOK46K35lOcmAt3TztiIq+Ws+OXh0qNCjcUiaQ5Hil4ttscJcZVxwWAHuFPTpb7gycVq2uMUC
qSQyo40+NekJUtsXStuDpq92j5ln6hZiq/IEOVn+9Rn6JPmSnANJT+6Qfht3yjaACVS6sSqoBdC6
tESCOopR5SB0PS4nlm8ko/dCif3l/eVo1W+cgg+QNMMQvYraILSV4xljqCmE0rMcZCXDp6pYiNvn
MColP82A/s+JaLBjGJMLm/RmetpxE4JnTGXUGXu+y9mvV1bAaSri/MRP+gzKkTZ2wivF/2pzjgg7
kzN7z11aIa/k0xqoyvWcNoBRsvJf/QqNszrv85CB9AuZJKbTJThhR9aasPVUQct+XOYKp3lSSG22
SvyKLqvCLI5am1iEpvj6c/Xsf0Rq+Jf/77daOgo9EWp1fQ0st4cL9T6sHSeHBn3UR2KskHCkRIfa
heC7/bnszPPTx0TIjvetOhr/finQOlJKh8qoK88SeiyxKd9h9HmrCUe/tDwjaGL16jRVyfvIhpzz
uS2iB+1JoXp38yHpkvguoG64ZWFZdmU+7TB+hcR6DRs9nZwAihBelRLzPsT4mdGRJ22xI3OUonAj
7NqJfN2eyjVPkbwY5k0sTXrMeCN/xEQrlVEhBCYBjZ+qj0kVYU3xZgYit5wE5m5mqyc8UQSML9vz
1Sk/ktWg4R8dCKBwm1I10/dj72rvpqyAUqMksrMhJ9wRiEwr54aZmVE6CAnKWuJE7Uw578YtOzZa
rmBFfvrgahq6ljzGkTC8LVuAH130S74Cba34e4xzY8bYM5Re5d2/tYQTmgeqiIHlxyWdTT/smaRK
atr+IOh8NXRXyAlXlPAtiimb9gUM34ijMeBINC0vWcfehalkKXutFcfLJhcH4NsKjx5HZ/wvyWQ5
v8ypBq78ql8OzKQT8Mux1hjCKrHZzXBZzrqm11bmLTqe4pv1/nPw91AibGfjUhrPaPflCucFBlzj
sVjJfFYnW6ca2KXzGNO7yXQPBFTCCAetGXpnLmWWhT3ly5LL1BzfVrTs2FSFtKDuY5s64K3pO0Y8
oJCA/t7icDMAOsaXCnilHID2I13t42VIz4xeGMwwve+5Pf6gZw7OqbPfxaw/2QavopvjVNmBxPcY
7YMkQmMetSKklHRth5S4bhDl2Xm+1yOKrokqkiBPEWxqEzNEqIvOaUORT2V7wzii5GhfSsj0SCc0
R6qc/9QQpxBfOP6h8dv0LldrkHsDPsto1y0KOUty8WsrjTmFs8YddWf+jezWzMtrcJQoDQc68inx
7IZQgu5qyVZ9ZDps8gs4uQqIXYmykRd3R41CFwZnrgfywN9MKO/YApxFCpd6Z+3vNScx2sVhQuHG
5WQX9vTxfKws3zfnhTDI1KirEWa9UiLqTdupfyrFqZfE4ZS4qoAvzhPXKUDQQHGBxcsrJizneMgn
bNpQv+HmcwFCgOj9SNwjrvIEvoAihliYmRN8DfpmtUI5wzESeqH6CYxojBxtO8hZCzYdsj13N8g6
/stTiW1M6JmAlSmiRWAwHGriP9jGHyeyVUT3qa1hIEA1ghJQqkIGr21Q5XdA2NUXEOybXpHQ73E2
L+sBYLe47DM70BC2nwcSbPmm5MsDVMbTVZ+yKLhz4MKIEaDJ1VY86ezxc/W5YZof2UAtkl2pWbBy
DU6RB1Fgd9XEvanrcaVKBdvSXhGWkFgWCcxlYJ2o8O+W4x/TRlnUvBL547vcAY22PCOfZPH89Ogg
rKq6wx+cixp4pZ+AsexpU9tDf6PgfQTxzZE4C7yxTqd/2i1W41UTU6EJbbEY/BTG/3zAfVlMf9ym
Gr1NK28lDtblBX2mIHzwXd5IBDvPg1QcC9vylAQ/e7NER5aJ2Yl/Ouv5OKaKa9mdAIk9y1zAXaFK
p2UQVgdcbnPDereMAtLx23RTZrU+edsHwDk5L3rTc/qIiDaQKPmi9Za3wz/bNvsEcZa2Tmzfhzim
WA4v+2ozMQHozM841HsQAbnMKyeYgK347aV+qi0f5GhB0vmm94kbPeIZ2FOO6C/foVHgV1/K2Eag
1kpSlwV+OdryHQSptvqiHkKEgB8g5NcRWxopHNdyEYdu+fuSWTLT6JKc1nlZ1MzVv54OuJ4XwI+i
OjAy8iuUV19MCDKkimcFg/+PslJlhfdCgkQmzPYq7MsCOXatjY4bXsvGhYnamEqq3RM5mTorBPmR
jZ0TJVgE1yFqyI2+pRnBrxVCOG5wKuoF8/wQXvjxCGUbyv50M1uIMvOZuX3zsL9IpUoLNkN1oYKW
1zEPhSJzfSSblIBlODeSb9mrB6s/fVUrogGELXAVWoARGn+qRU5mjFnaA4gYsjyMh0OwhWpNeXEa
NgFa/yN+NR45wW0W5iqVpev4YBE9G6L5QlqWvxBb5thLv7AJkNuMKZVUC8f7kJ97/E+Vgj5gva9r
QUmjQjoEOPNfxGKmE3zTR5Vvs5tvPA1Uo6cAAjNAMHitwckMb63xWOUcqW+w4sX0PhYIT3lyZNw6
Wz35wUrcMDBPcMJy+zvE9t1p9g4UoOxjRGJBxRBlOB5KtRXTD74hFk960iaeGptAkHeiAUcE7IPi
u9fFpwaREx3j3B5wu8Cy9BC5lP6wvImdXxjMYELyCyzjB3T35IAjbVzInpWlP6XBog+Hqa5KlvHk
er5F2mPmAgCyXuESbhiEyCWEPDTZz0kcRzJeoIvmv6ZKNZiuZ77ZNAW9PcNAaEQpC/NxMtiUG2uf
gkDAf5pe+7DSedqAuI1O0ABKwufSr05hLScJY8FNZQYtj25xxn/We4xvY/dvg7ytm2TIa35tSSV+
3yM43eGQ0iFqTcOtV7N+4fI7ukAXcrV9hCdf3M8z564Lr19ps7SPPXF+dcJlAHuucP8qeQli8hHc
cfKYytvBzU3FRHjmthLvabVRdzNNvfxJlLvXlrnsbyF9uHkGInX5InBp5wgJ28UH5ZPGSLXSroHE
dqWTNcygNkp+phnArVSIbGIJ1YmA7ACY1ajuxZyhtbgdcd7KIqbOwr3Vsgu0sr7cK+2LiiGV6zQy
jJdB2xr3FKlTbfDYvZxP3dDq6Fcu3DX6x4/AZ95FSHO2/ktIh53WmmYeHgAVyUrY/EhxuMxTWTMV
1Uoz2ftttv0jYPxJuNop2L+a3zhs4bMF0QgAh6J+dkWTVEQnHd/9OBB7lmEdMeJss72rxUIYyGt/
kPfO+oT3DQKo8Miea5GEAvQpokoc31iFkLbwjqKd7gp1WngnZrkyefMQzOwyxndUX3eDO0N+Vmjt
A3/iuaBBokmEnyONeVtQx6C7mw6ohcmVFu4rtziZ6xwkFee4kYCXK8ge96rptvWuiQqO2O0uJwGd
kDUmvWKCH3XSBf5grl3Aw7Tzoel6m4D7t2Yb+9tMAeiT3xgAhkKp9B/4dX0fnic5MVkhkmHdEoLO
/HOH/+jQEvNqgII0CkVovNA0TsGScilEQrJmc82rig4k7kOxynRB/qgoxiURuZjHP20WuX3sysdZ
nXIIuTrw+mvuhKwzpWT6gQ8uhBSTSaxITF8JCIQX9HW7X2d+QmU99att5h3/Stgk8PrxAIxU/V1d
Z2ZCa6TfU8z1Z9PUYoviHHTPDN1VRMHjFNGfbcz3isB9p6u2WSckEWh2RIeREERxQK05tDp0qoCN
8JfRp6iEiFa+FIN3+K8OVGBJrs6cKPWB5HDH7t65Mrg8e2XoUMXNhXtLpYSkye+yBFDVqyPA8CP/
FXWSuWerQgXpYus5BLUdw94VzYMLgdqpsIAqAGieHkGndt3YmenARtjF8hjw+gsMO+IU1H/GPh1S
HzMQxS1aFEH4s/cEn2p38CD99NKhX+IM3p5QhqPCa6m4G1n7nTILwLiYnJfJBLA3OBNPLXPQ6uEj
WBqR8kbIei9En35Y1qhvDMDmwXca3d5dEVAOTfMJGy3HMf4O9MEW04PcH1lqnfdwRqsDveCYqque
QCqIon++LM9j7MoXsznXMG/WqcHFgA4WEkXjCDFmwRnp6kF7JW7hIMCQkxMtI8mAIYGplFvv/oKE
z9CG/x1sBvKAAslm4P44qzJKfK8OBDTUQ4b4yeEn4dHLTzknoqw0fRnAIHSs36HZ1VHvEfyE85Mx
oiYq3PuiEjSbzACGR1Vp/iwUcO2js5K9QZBOPsmOyi5pXl2VLwpFyPtyuxxBHVR51VM4pC1eaGwt
cK0Yge/mUV7BQc79ReDAxIF8LYwAiMCKVeHHT8kGHavPXwrPpfWmInesfp+72ISEz+GvbOMfW0VL
lBKH/8YUOAG6a1t+LGAClPIXnLMSFMhOBT6ut3L2SPbgjsGwic3Gs9dDj/9r050LSEnxgPzuttqt
8fZfJamS+nzHy6AOjgMf6pFlTa3vmTl+9Xo4IRHnXfTDv0BIjaomBmUhAsKK2Z8d4fVdDrCgVMqb
X32AG4JvExTljVXnrqtX1Cof2aV7M/HUK3FZny9qWsit62GrT58J9ssY6xQYOzOUojy7mUfK/zqw
xclgmBI96qHndfhNi+q+U/0aaxdtg7tQpoaVVIatYVDvAdOTTHj1lSImBkZg/J6yYbigrXSowxJW
yWQz1yi1UjaWVJbYGb3DcdDdiH/79qaLmxeLQEYF4sS13+Sohlb0Ty/8WAQBQJCpxcQRjtWM9yp3
5PrRfq/bt+wy7CFlS2W0Qxv6QAFRToca49dSvGLSTiLv1WLMNmpcj0SQs8Nrs2zr4KO6/acTwJJb
zD87ydmnTryYc0GT3reesYcZnxq84epuRbkeuWBWsSXx3AZGQqnMLPA57qJ/xLO7jxAAjxIBbG9W
HUn/MScKonCJEVRPfgCvk7H0mfs2knDTPjDyZAprrub24v2JSQ9AaepBwxjM5M69T8Y9J5SvTGNb
pytolt3wlQcNnqBmbAHu7+5kZ6dDDclqcBSHLV2wEQybr0JCCe3kScAC56znba0Z8Fxjy14D8hCq
jABAbxHPWq5vzIfVtU42tVw4wf+t43yirr+oIjlfFAWjX0ExUYZExLTeHA3EgemBSbbNbCO2bxmM
XHMt3BUVxWxhAbgVsenUnsPCTTfa/fLG2GBWUKjuOOoZG8+z2f9jm+/Sq0bh1+rZMiq9f7yUuaqI
yOMyxU+zDb3T7fDRpZgAGAOcazWB/KyUfbk2V+UpJjVRo/TR8+XusXIkj6Qy4wOtcE30di55YXQu
uY1Qw6NXdmGdJKiYA3jkaABuU7lhnzFzwxEbbfhza+lWoPCNjPaK7cidJOFuBeeyRzEW7rPT8w8j
LL57/sJR42FtrjR8EYrp7oS3vUtI+XM2wwXCL8KYf4yBeCkAtIPR4bwzh6MfeU7+odiJ8UvxfWiY
x6owkTW9sfLeKkSA4MldKGMvLfVPh2Xo7msGUFgBw+vVzN4Pswb94XFAwoNsmr1Eh3vNfjjDOVyw
loEPaJd4oCPNNOMTI4xR6RaHLu/THsqcZsGod2FNQg8wzJUC82eAlwwp1ePAeuJ32/d3uhjRwNlp
CiwNlqBoJaINY2zIfiVroKFbAqHdsmd6uWXi8tIHCpdJ42w6Bfvrjw3Qq5fYMxTh06DIWFZpGMjH
rnyiZo7I9F+zCpfA1eL5sZX7O/SNQPsFjOfeDxw6Mkt9lNoOkw3VBWZFmOXU8hZbcRXn7u/RjN7V
SFxpDBAwcOK9wai20+rJ6kW2TiPvO8/FqPeEHiK+0AhNWMst0/WcVSO71BH6EzshnQzyogjPdhYj
vP+x0r0MuaFmtGefCuPyCy8oYPR9B+03VUwUYx5FoJmlax8WTlPfkFrroik42c7Mm1R5VYlY4Ekq
ucIOPy5e+YKazl11wk54sHfzPNgA0MSd6d5MOOj/SFChsFiDk2SAfvbJosCJSsUTeLsF/Q5nqQ2M
eaPqf5wUqEgMSg23ELRhKqVS699X9EoVa0U8fSJbNSDUw92GDQcwmoPdKxzGdI2CB4kJ4QbaOAjb
LlaGgmUZ+CRcjQGhTQYrBROCW2+hf9d8m1NDQUN67t7/NitL+JvzVTfjioOPiSQB8H5z6hlmsT2a
hv7LS2exPcLrZjA97lsdNV8Bl1rPpH394Rz7ixPD4aFITM5H4dSg61EbIca/lVJiU2SW5AzDZ99c
+oamDv+8OItzauLbkMqR/UkhrUXectW5ZxcBpbFTLk4oqj0UBuFO89crginILaGgkq/bFkMllNhm
XlpVPouAJHHKOn466mrpVPwYG5R6zvhPEdVVl6LEdvYNKjXcKNwALb1NQUOVsHOy4XXO13N8y8mg
LmGYKPnTsVyMhsza+ZKsKWKUNcIyZl5Zj5dGHt1feJ/AlyRzf6lFKrscwD1eTXf3A848JNvxKJHv
BL3FaVdE41HlcTQ4vhpPo3d3uD29F8pYPksyZ4Tc+l5XqortlJdOugpyOIgIw7yFiCRBUj2++znc
thfFPp3JU7V2RZt89l0FaEjkzLHAMLKVxrzHsp1hrRWYtstocqD8cfFxJFImmJsQOkdLTI8Tmqud
/ylVSAD+NIsUVoGvt/SheNnnc15R6sjhbw0opcbic5VKOJdkfczgY9wIWuEuUFYlxgj2cTP41Yq9
7btNBcViklIrh1sA/Ze1Jjzb2Z4OYwM/AR7+x/GsuscXGKjxUbMSCgPElU/LTQ5uCf++Ce8i5CkX
YobKMUkhVAmWUNiZKudyy0YFvvlwvrxm40IdLsDve/AsX98ZsvnWeP2ygZNP6Lr2xTNDyZ0p5kfb
SdYbtwceTfsUwYws8NGGWRgvUvZ05lUWCYN6kbq0/dtts3XsnKvl1OZgo4efYvWXogA/9zclBSKK
FsjjRb5lCzKY6P//9LLSfxFfTpxzJ+4rzcVl0VRchPn3VwGW2mHOHzrV8sBsDJ7yUsYiRKOkjdSI
0FwEq+uz6nKXppL2q5dp+xCai37usWpjB/fkh2CNbKLqf8QuLbTc1AwQYhVwhUUVZUPgR+Bi//hd
1ypkJEjc+NOrgSq1mVla6JNFyJb/HM5S+3gf7n7mlxqNXllMDpYda9h8qBJkPeesOpWpOXOhxzQ8
r5ej9ICzcDdgHC81aoOyA+74izVWDqZRRQNaalTU8qvKGPTrIyCHuL/COFoPPTDXcPPUTNVFK1gi
de1gsBfit9Q6mgSeLZkZIgWPStyQOCKYVRs6EOWJ421jBukX9ufpOAFonbUQLmVHrwwh4wBD2/1B
zMtgxv/z8XuH17nv97nwRiccLpGNux5he+GxiPgTT+LGN0o4p2xRxdN7UI9KC/DtWfoyEFAbfZYy
27FijzVWH5QXe//SY9Ram7SHBhg0iPm2hI/e22ojn1XeJk5pwc2bTZLq2nZO8J/tJqfzn9RKHdf6
2TYkT0OfHWW9iDlin163wRMCbVmNrkwwEF9mtQc7s/Le5iUJInHEViQc6gFhBojZFgEps5m1CfOu
eT+Y2ejGn4ezaOL1krP5B1I3PS1fp761AuUCgxRRlQoUym7zbVKSIv/2VIxSOCLjyTOlNvYhy3l1
BsJ9wXR0MVT2Egz7m6wQSfoLHn5C1vkq3x05+rI1cwncOy753wN16ZjqGkiAJy7E8/h+Q8g7Chh8
3SBqtkMpj27bdeq9XOezLfWMZR+3LAMdu/IzPfSCPy1vOx4z9gvqA+lNy8ps61Ftq9tCYHqOdDWQ
57Cskbk0QWqQ18hndBkd5mzU+jAHLR4Ua5u/hpWv9yUFWV31HmdXp54nINyuperbFuvqtTETszkL
JWspdnlrE6RLsye3Zrf0XjiwW/wDUJrlfiX6RJgwYhzlKWWQpDBh49l+iJ1YZVkh8GrD6D+sFWel
Xhsh5BgzAxWliTvTFFOvrxUqCyJHxBHScvHezSet4Flenm3ezGqYyNnL9+npJM0If+7F4iYsUtk+
bkxauKPPNkusfGwyTZtewKzIeh6ptmXsP2FmFbRj8sr0NOecJXCKXW9Gf/4y0atH65mwxuCfbGez
btO+kfG+yb9ASF+96R9bUd6IOyaWZwuTRN4nN9LzoIOOwo4NyUty2boBs0gLt8TzDeWa4dunOy+p
lqXEt9BT5JYT0ZF8N/zVOIVbfS1+IyYH0wNt+A3eeLqIo7xRLscYiQ5UOvJ946RaCVKFwd+yluo/
B+b2CbrV5xlz/Yy+k55eByyRusk2feBVoHe3jEPguP1rq6x/SfagpFekAuAA5VBzOOYhpuvODOqp
1zgpGkXYNqSUt8F2xxzHDB5Nv4E36ffXTrY102bN/ZpItORYuFeOhPFp5jRir3YdlrzC9i2FEqaL
QLlWflOGRL+HBkfrfc0B/wVchQVVFKrr5WZAUngrv0zoRzzt+wBHck1w3kpxji1oh1Xdq9IDkX0C
DkEH2P+wd6rGDDhyBiN0iNhgdf9pnxkUVYiR3NjJhYu4ChWu9y9mM2t8VKKdLYVQY8+8xpXU600C
n+dIafOtrfird7hN/j4SlbXtyH4tLWEYA9+PbXuQgMyG6Xvhn5/q2I6c7MlAsGdTKyefUCQ5l/MS
PjbK198PArGqI/6CEUIvPeBUBkUhm2GdXnCbiBWyhJ14jHhpf93nSnUCwJNx95V70yxsOh1CEqRP
vlpG2ojAGq+ynP+eIo2106tY9PRtmgbQQ8lgIqDa2Kw9tvLtq7kAkBnH2i/dlKA+zS6MwPfV407k
crBodxkcXps243NkSHgh2rjlPZAG2JD9TXW+bQoIHzcF4NeFsS6sAd5ArTburs82nUAFRpMR/7F6
qIw3qpszRCtBgjGBTCz7NaD1SR73zy14WEmtfzpyXELjXH38C5lT7iCgyPrvbn1S0R0KN/84cLhD
5JBrExB0OBs3Zon6QDJc9yzlXPowNI1u49UFGp7C5EMYxGQ+i86lwI4z6wEwk+S0mibOgU7IvUmX
qBgBxEGBczhuQ6XGauLpHHgk3wEt25CDYpWKinrkzGa8TH2n7+oahmNTVMO/4SqfAvCqhUklLawn
RqWLOKEiyiJtNb+dQY/cDie0X20P52H3CoQigCE16Ssfd9pJWW50hrLa0FFZb3KVufqD+mYoO1/h
405RwaH8kTVur6XX5Un5SSJjYxUFJ0qjznlxTG5MXM2O0CNAtSXbTB3lBP26L26Lo2Os53fgApjv
J/U65GUs1aRVrbaRO+mTPjW4MD4QxSaVF1q9iT9uOjI8raC84XrI6JSHtF/vSGY09Onx1HRb5L2K
5ysOlGPahnnyJQwArawusuCKJ+f2vyJvJJd5DaKs2Rou6SQD5M6POwrIgk4ePLi84QqVQqiMYoXi
+Szt4XsNaWDQPYa2/mABnpMEdP+j8OOomZznXhLYM9SESzq9MXYfU7QusjZ13P5zsZMmogOT68zK
FO3cfHDlV8v5nxl0XWYzFl6EPFp0QXL/jSKyUqHiO/1vJKijztItfRPTl0UZB9eDt+lLVvQQioh4
S9N3qB1AVc92epDFdUOObfgVnNj7s0iKSS9Iwf38ejnm9JjhK1R1YuezLNvpWM5z3Rvvp+NP/Yo2
w92Y2Yywa31ilj43I4dTY5bvhV38zZ367GtePwp3ZkzzOa3Ntatg4vYu7y42U2dgTprNwLHlVBYa
Q12JSxzhzVd0XTxd72z6rPfjwMrdjA79ODP6BigLzOHIelTM5jc/s7VyWKdVdudShRYF8zOCgvbB
2thEbkxAouO7VwsIhimXrMnrB6JcmLBYccfOSZHZIjzb51sXjYv/UaxW+tFp9wX5sXuRsxQ9tG8c
QdG4otMIn0i+Nu6MN3y5HOzJVvLIDo4FoUNy2u5V0RUuhC7sl67NhAIUMZkR8ZkXjHGc8yKrWw4V
vzPCVDHmQU1AD62Ky6CaYufBipy2BkhGOFHWZSD7JmNDY1lbaRLIDX5WSQpyVxY4PB5YfcC2px5p
UYYya/4frn+FRaAVdkfVeHZAXInrqS/l4nlKyDr/qnXGhFab4dQhmClOAg+90a5zQejW2eq04ABd
BAkQS5QvJE/vFZAsQgMs9RoNHzpdamj3dxVId+ESjms3XaP9L+NHdCxieGAcym57wR14Oxlyw4bu
jWv3/FGoCvj6adTmOdXSwBGJeeeXZ6qRwHbkpINON4RZ5QHYsYOMOuJVzCvyoPjCLFxtnm7mowZM
739NuzNyIzIaBTQ9FNEMR+v51qT0sun7YqsU1fYr5YO34OmbA5nblRrAJ15GiVr4aF8+JaxA2x4j
8tNq/nXh/niXzLAfk2/RzKYVDdLeXis4g0ICtpHKBF4VjdtvapxbBv25hfh6386PyUqkLY4/+Wt0
oHg4KIA39BI4Uqe4eXNLR4VByx7ts7ovgZZWaWhIwABJm1sh1GFinVKxlhJMc2/8lO+B/RP2Zi7M
K4ITuUs1eKKsv8ZyXlpm/bFq5aar4b817S3UlCOA4sIQ6ZNjrXBTYBRRIw0HDp4XI43t8AGnIkhV
DBOIG/0E9yLRK25nQ7Zl/ZLdTaopBocG0UbaJsu/UtiltuPfQnfIFp2LWXlAHWDRVHmySXjI1dZt
TWZYkg4xJDP+W1G/Q1IZqo1SJltky8n+sZ8GYzt7e3l3aD5K8SUECQjFgj9cr/dcafKn1GSo4uWj
Sw90GMh+4B8dRjvpMbExop+J7Gab/Z97KuYaGQzn+xGz1Wxtdsh15CXFMITwznysPfXtL9NfW8z5
gfwKolToggSk7usxsK/Ca7mFnd1nDgvypXP6DiONVcD701oVToeoIXpLBIuSmAG/7cNV5oC89J9x
yseHuC9V8dBck6MD0FHpdjfnhCY9C0CUO/mfUu9iVNeQDy3ANRzKsBSzcZRetbxy4vlzRgPFPsyf
ZDR4kVko+lQLiR0f9Exf6v0OfYd/mZHSn55ueapZ79/uLQZS7K6dcAFgEWivadoZ4M0tozK5mZ6t
VDJ8YkOVtFII2JPHDRhxXmN1P6SX3+Kse0LoQ13zdtjSAnDKMChzK97GaNZdd5NANp1USHVYyJ9e
fcEzysTzUvqVc3Up+Zqq3Lpd1hu42mH4H+XchI8003EIYFQ6FfENWV8uSwMh4Xmx8xVQpGt7D+Sq
avl7SqS2b8m56FuBkxAkLxUJMU+lCxNTEIJma1u+9m3/IH4AsWrUaWS5FtZorKsQjphefsVOn1X9
1WpB4ujKeq/02jsW9ocGWRckNnmODpfs7+Rl12iQnorH6kuBqENVjkV15VZUF0G26pyHxyYl6ZZI
SD/yj9qrLET1OUyOsomqXD2d/x9r+z0vQbFcK4qT2Zifnxn+qJ9/5vw1KH+7X12OfTfsKqjbnLiS
exyaOjVP/+Sv/gM9pcLLb8fgMGAnoiDPM27l+SEoaDg4xx2p7goYHQ8Qp/k4ovnqyEsgg+RQv/yc
eNrd0d+KksTUyYBfbuMmMRYkZ3YK2nJaN1obeo0/Rb2gO9aoRlNmYdcoqGcBxxcraQ+g4k7Jzlfm
M/qCwz+vINqnRec7d3i2E5c2t2Tybg9vgUT1LHLSUWZClYOpr6Ue/Aza7YXjLhjn5TG/3wSeVO1f
Jc33IMapBmSjDh/DbM9ojhrRKQ7xLG5jU0b9/a752ZwsJ6Ri25CF8IJAXxtTHP+QPw2ymF+C1H7U
cRUK6s1yhhpha0KpdAOL53d0uoLmSx5nU8gIKMw+cBl8Yzgmo8ypPUiIx5TDBIrkaEfvLbQmkiat
bSSDgxRi4P5LOEURxHs6D5d6dOenfvP5OAw+r8IY60v/jdJX95IBMuUkS7OfVwSXK9q6GA/kCI2J
mQMtWIXb1Pg6FqeP18BCzV2OU7WFFuBRa9Ly07yNhod+sh8x6LjnNZ/NoY6pqxZxUJPj8L0HJomF
L7O8yqWpzQl792Qiqt6/wat6kc++boUjUyMoItskfg7kNDVp7NCVaUdSkpQRFauq8Ky+E83B8rso
jc8jHvxZRZ3hRHlCZ8IJtQSQiH/Cpl0I+6+MP25yiXm/tqzRz7U9fL6w/tJ50628ec3u3w0/BzX9
CPiwgW97GSPH/OqoI5GmE4ENlhX+wa5x+BQmSqqn76wXBIw/oJ37nd6JtnsEgam7+VlMcVSEqAiQ
NqfYkNUG03hlvOvdWkzSMM/WjSYtq9yysXqKXSXak8hqOqmmTGMknCIxe4CRsuhlijQ/Iet/oHrP
eGDEINk/UuhCQEnI/LjJk67tHBt4PYwIKGUnj+eJ+1d+0MZQHRBlA3USrtNPs0WBlGlUCSr4INCu
UwJiiD2i0eHdi7OJhPUjYgNEGTSub9t0O9twLh1Z3uLU8qy+FoLkFyHSheOBswE0HcZ4EkK86xud
/1FBwuzxR5TlSFhHlMs/Ng+zX03ehrdhrMNm0TQGo71yBCMxuOAqXfFVlIezN91j9Uttbf03KRjz
lme76uRKG7zHFAnWeWJA1h0CrNUJwm2dRoZ00wKDxuAjZLPiCUn/ghgjySCSZiLqyzpJBOMGNy3r
UcmOWwb9BIgAlASw1xhZGkNbjcILUVeWKs4NynEMVsggivEWuJHB3D1ueD6PHIprv9XTC+/tCvK4
h0d7gAGafKUY17VTEJDg7uWr7eJnzv9Iz2OF92wzKlTRnQ/yP9Ifsoe8IQIr/QVBEpm/Hy+Yf/Q4
cDTLxjLvpbuqiwKd4bTwPlQYbHlg5mP90sVYo4cTPZsFZ443OAJPdmVGKVKMbPHYeDL3m3/R5/xD
SA3a3X/qSai5NMQr0/R/Vib5m734tWe8CDQyVr8uZVOR1GkcW18W2Mgr13Nt1yHQvjFoisX32dS9
FGFN1d2R0PnFuMdV9TvEkQr57qX+srwXXNe8XUsM9WP6rJhttX5Npx8BjwLy+CxwzpfFd4EseEyS
hb5SvhzHYxJr8RZxvABlQexaeknwZYZZu9M2jTcWoqUKQRPhRC8wmmdBVONnY6fFf6TWJWxOc5HZ
SgFR1QYbPAQfnp6jEpLCFKpgy0U2huhUdqeueRxJN0yLEuudtmKN3g7YNuLIrCDT5Uiu1mJ2KEQx
BN9K4g0YCaOg6fUoD/mQ3kIMHbY3qVtxAOt6kI9H/xDEPQ8sHhAJ9oGr/WFcfzlwTC41BDSfMvBl
MBx9oG7yksRsW5r72Ny6GWULnpeYC1yEny4KY+WiIbnHam5wS/Vzcxp97SjaD9oZc+8cIJe0O4u0
XwuZOzo0jXh4C+jnHYWs3METS2dMOtGbQkczOQbZK3QEyHEef73jvMQn6Ygl+99PipfnKfjVujvW
DAzDcbvPv49d43OqlI4IUt/b4E++CsL4idghfDGcwzDMbBeBFxQycz7GzqHnFGCskdtNGJP3GM7U
x17Fd97A/PMXSEClE7qNodFlT40B3RdfIOSBIHUrs0Z9IDgUCG/8GvLwr3Qr8GjC6rs9cm2vKhDd
Kg0yrI3FPVqNsO+sVsz25jzbYMul0BIRGJiaH4t8Lcfrjm+GXot3ahzPn3hQl6fG2xpogCZYByvT
M94lvS5hBUt5JBkYxJ6YItwrQuS+LD9mhmJHexBTm43tT2oAhBzvc8uJ8wNApkeKM+c7o6XqdISO
e0tf/mbqaBU5bLodPz8rH8XQiyU/w7D16MxN5o80xlrS2ofguJqezvVgYShqFnCfDo63z2FG19qx
1DkHYQnpH4ZNTgufSPAWoclHsB5FTG7So2uoRFbToC6B9Gpqidr1+p/STDBAjw6rRwa62OmyFYB6
VATt97yX+kbP6noO+1tTklRQfQKaLCehXeX2ZzjTzCLNHnQWCPFcfK5u+B2ScnxPzmWeNs7I0mBS
KimYqLIGUTECI2dtc0Snt/ASzXVey39bKoAQ5QtbO4x3Y5VjJbjg6hRxyB8S1Vpu3FnaACyPiNwB
o25wzt6KXvkmwGpp4nu0fH8LVCWs+8EN+E1JPRTmukuX5V5NFljVAc4oWsihRAQ8Ej6TiPIJIzaR
MWTpX5Rx0iVME36pBh4BgEYReIdCVoVZft2iME8QS0R8jBWB4CersFGshTI/tbKcc/2hBtlQYvk/
LGeSmVUU9k0nZSaqohJ/VWKojpCMo3pzjDB6Oz1WfgVWkFHta9MrSLZ4b4nPYdcyUPlVmP4WWyDp
VSiPh15aN9XZyc05CT4V8T3y7/D2hfiVpNq6oG0ADM506bhz0QQqd7nHLU2iMTNN4AnTt4w0U4Jr
4A/Z5Cjidttu7k+EjnPhHLZMSPbTMQA8D8vF38R7BuJbdjUufLqJvclLVg9XvtjgIzu15Rb9+6M2
rTwwIe12XU3861rykCbOoRm5iP0fPLjVr+bGEZ4FCQ3OQbgmW81FmQMC3G8Ahs5hVsgbGoqhxiYh
DwyhpyVhqCzLKRZSm3mwimkZELxqr8a4ydNHD8wd9DzdvX3gIke3vibK9NnVFVasM5mNvXcSpHqu
mf/ONXuMNrFRtioyILQu+l48W+eRO55hXahN/Se+gPzZgabeMg8N7qR/X1Akf95rJjvYGpu4klX+
ZLhMqzeCxMjp5JDcu2H+FiriLCqTaSg86+EYVPJHow4sidod76IZjXimjV6SOYU2km/OBfAVpjLQ
UUuu9bg3SbWVwK51zqr87AqTMTZMujYtJ5KwDNgMP6mMaXdCUq9+PKqerydE/ccTZ7i+jE9NeyDc
Cjw2ADvEZec3xRneWcLwanFWIxhoJjkmgU3MWmVwJ28hsYHmqPVtZJ7ej4dqEw647tD6SKAiHvV2
vP1k+zvmA2KzGusnxFdY2ydoQDcWT6dYOkmN38LfqYJNwdf5Eocm/lmBzHehIbtKWNdexGqzTwMd
NN+ZmcH4DpMqGXVzYtflUARXCMB/2vNjTCjhuKpyymgZrxXaYxyjh8+OyIJYbxTPS05FUehGHcXZ
ZfogqRjAyOpoxVyGAhASgVa+tzt7Hdm69kR1VIMT72E7/M0Nlqf5mtjbX1YX9hlDuTVmGsdy3ENv
MYkdaa0+xanFvkhBcr6qJcWqqqZiadkrPW9epnyNpwZI69gw5d1VRQuXOTvpSx7FGFCytO9FlPFd
xjJMfibpGNOYPjgQSzBHexb6dmH8rZHwiBqexGkY6y4TEuhXfPT4sXKyKJfS4iZXHalX92UG4TfK
kP87guDN1BdRfJXqhkOaGf+TO14VqO4BBJXdPCcMBdKegYYe0f6lJrWhEJGSDmt0Oa/cuAivpTE0
ShrfAQNa/Q/yam9mDPrLo82gkIhkN4SlV7YMJvbna8hZG5hcHhWBn3D6rqRWFfrBwRfTG7gUrk5l
rtk0ZBFPeHFZk4wm96FsKzFr9fcQtldWUZEahz1T+qhP2UgRk7EAwN/pshrqL0Ru/y0DE5GJ/g3x
ztg3pIA9xwgQiy/8qHEameQa3Ywguec2TlxxYaCNSw9bSWyRc4WuNQxUF12wRVv08yBcbGjgy5WA
nWzCii95Z8Vdk4yBYBWjd28HINJ7yb4tVIpIgFyINjPS++LglNGzKIK3X5Sakk+yOt/W+HDFHkvk
x5vUvp4exzO8WgfuIdBRYT0cGDWd2FOOaeTjfV8YBHBladUPvznWpr6E0IfmP8/nd/ta3qHFmZUP
34SgI9jbLMNGQH/5CgsXmANZiUgbA5OhtxBRGivXNnnSY9suIyq8MM3olQA4KaZQQSj4oV7yYd3p
Vh0jPJ/1CVE57/VP5+znBRfAbL32L35fL6VhwNE0na+bIIwm6R2JS50AdcCunvT2BE7XKv7sOqev
gMlrSbE/3JEJ5jixurM8BpbgIvcGynYdkgy6pAHCGEZv5BVgv3M+RyRxJAOnTDHnRsR8IwaMBcA8
wV7bOkj0KlO3Q4Mk6kg+9l0uKjJSkhvDg+Wop40qk4xFIVhegAVnddt8fLas1ru6Fq+99gX0t1Cy
nZOrTWXArwxDzQrTd1TjBeOfyiH5FPsxpqyROefgS3h6cq/UVXSpRPJp2Y/NlVDYj9BHCzrVP7cS
7tFZz95sjINZceceqf3BholMyzyz1ASxJu15pQkDK66XUD2oLwN3mW0EP9pG4NTLESJZkwNZHBmr
yd+nVB+xIcmxhptxRvLSPjtiq+ERg8MdplG+UlUuIDj+5ifL4yL5cS7QaxV6qOo0zT8TJr58kEdG
w4VXncVk5DtLFm0ySrDU2rqVBmdqhjumtWFkh272QLINvDq6XeCQGOcFlrXemWvTRaEG2Pt80XC5
BtOumFExcRKBrHjztr0d4b+Qj4pzMUQL8N7xyJzbKZ2SuHIYdj/F6++5UEroX5/gO3muTYSUHo+C
jShs6TdfX6QdEeA3R57cLuFQTB06P4jns1YAM+vqRuncwXRthfYeE16E8XIFkNytRK0ZTY+P/ULU
BL+aRWvkhfq1Nw7BqZcjnEtNl/EYYjizC46iXIZLKyIS3mf/nH33YGqntFYPdr7cQi4/umuIXhU4
YovnF1OddNmMZ9WK8kLb2wzf9XwYBJHDsw0lLr7Ptuu5CkBKkYsi/cJKmdnQgkVDh8J/dsk+Q7n6
hwLUD/puKQpc4z5/5qEqOioOmVDWohlLqEHpXWMUR985rQSm8CRZb++K/HCNePCsCbsFz6Z5c1BK
r6OAtQrZUwYh2OfntmqwJgGgihR/NYZ4sKeYZnaC98TFTGsAbn2P0vHQxkMx2/Ub4Y26521w4tD1
uBuwQmqdmWs5ipFhWJx+O/uZOyvDYumE14qd3Hgjug8IYSUD4ZHDljg0y8M4ljilfa+58AiFvN+G
ydgTakubAIBeMfUKU72Z3+LAjMdzwMyUfehNMJ5kXxU+QjpheqP3ruG5rjqg5nx6Mmsu1UDiIpjJ
mZEnG3TgU7ehE2Pf7HvuShBQ8bnhwP/iZyLp+I2pJgTw0FbJgh3uF4s0jHvOm8J9uJCJ6H8+loZb
fXwSU4I6vECojJJvz3neomsjzQNb4GldP5aZUSk9JoEQ/jtuPvstoLAwoZ4LbvBi9XsmPWsG4aiR
LNri/qZ9+oEiRcm1KONBH/0sALa74C7oxOlVy97bpxPqO2KDwPmtyNOfmBh39NmNx/nn5ehvPBjv
EVsjueAnUBbtf02k/MlWj4jmOapUbQXjduwf3eRKS3bt/Lel+3XpNIGe7oNOb7+rWT5psqibagFq
alJh44MzU3KX/JCCyauOgaJqDOVLTgk0dzeywHekgB3WDi//RKrgoGCElWXYvb0vv5F4n9o5lK/C
H1Yr2rRtHZbq7F4Hv8u/CrsGXcCHuiwRjNdZAAiVK1TL957Zyi2I1PFvPa3RunBo3kFX28q19shN
r0aNReQu9gYwrzE0XrMrMbbkmrB7uNSTugx+CTmuUn6qiOiv8G1L45uF84bRtnI53NH6vx34atrV
S7E8u6jN6uHWY0fTJcbpIi6vMOR7Gh5GoyuD6Ni6QF72Onwg7uUZgTKctSnNYQHuw5WaA8wgXKP7
BYNQmw2iWdLGz+33vr1RcTdZyywGPO5/laIXbzTcUWWC634q2QbErr9i5TjqtW978Qw2QDxTWyCT
VJ+2J5254sPnf3ncIPdtapJskQ3f4fNigTyA4YIZ96odzDTl9zh4kr+fZJRoslvE4NXucq3nBB5l
2YgRawXjj7PSSbG7qKMuNdnIuqMAk4sXcObIrEG8dzB1qlXkBLgLj83Bf/Cdnmdc1ASmsIq12AlT
TAMrwGUfFhCStMSB03A+awLJtPrUCnxjO9SRrt9fQAi+CW4K3sb/fIsGx6HF6uCec5IbapRPVGEE
x9p8KselhKfI3osP15MUYoJdw51H4+YXaAgwhFQTr9qPlItAmwZEJj68WF/BIsKvf3LL45qWicKr
sECgGbH8eCe0uJYwCHJqvdWt71Cc2P4pNeIX6E0hwRCLWh0KmPllY1czSP9gMnInwaZXRXQ4iIxr
iqG3p/8NGEoVUBfLmTK7WWNpIAPgKtu8GWSDpceYlKwhucfyTszBLEA5crju83ICjSksIiqS9Z4I
nXCAhnYR+6yDxuSSvMa3tc+j6/9GxJGl0IDl/gipKR0puDjCTFo2SRmM+njIp/AgltDy2OuAXncB
1Wi/95+LZU2JSnFxYPEbETsTzyOF5ZSjWLiUuVP3DPZ27pNbbMbcWoShHMQwZqkke4ftC1cXRb5V
hqCUb/27Hj14DXL7gIp3pUfbQts32qeZUKlNOW8PnI424VLDHAxGPDsulAgb6Cx7Rucn3SaTc47E
J9k5uMweTAX9TAYkfiUrpYVjzQ/1Cz5X/tFoG0tf6bpVwgoeK/ZrHc7f0b1DcR6I/s/Vxf0Xstx/
WD+ym/odZulx8f42E6gu814iqhTCZPs+HUPz4SFyUzkRRiWdQE47GWQnHKatvtNkVt6rXJRwTDg9
Ltyd9AIsmihoKVwP+Bz0Hd4GKyia4WvvsjaFl1B5RDouh8IpAFF+1qy0xPnXi1LUG1942EdYaVl4
y/66CKdzfRLSHHCQDTZSBVQ8o2+I/HxcpWndAxwQuREexguxZSnz58km+0MLbazX1SEgzDwvHT4m
Xf09RhhotoO0bTSsdQyuGkD/3fBPE8GYPiNg6ObZxd3S+B0aGlVVFQv03iG/2evXIIXFF5U8sroP
On4i1tcE0TMEfWFxQ0vDNYx5BBFpHwcfHiJUO5HRjQczLn0IgczkOhVy5irxD9uYhNtA1f4YHtsr
ZP0LslIV6v7NkmRyKu56UVoA/oRav924wllINmJN6r23OtT1jyRvdCptiSrD2aFyIV39qn0w9alW
hYpSMGDnNMzR0gbtkio7DP56xzDA+NuTMDDlo/fOsq6cSr7zqTS/rEzkCUJEKfBFiNOm19nxHyxW
AU5xvfue3/LazqoRSD8lobs6637oOCusTB64YJiCTS10VlPsUDQOMny3YqpB2JXd/BDVYs19npwQ
h9iQ47DLRkb925DwDMmDBl3PiM/ztYItWDzo+PpEGpfTfMtVfNSQkOpnUnjeZS+fqniWB9C515yD
6FaIdPSEr5ydWhnkIhstB650tzY144jVxAzPmKji9jK1jiq+aSunt+LZY9w90UlZDwAN0cavJjoJ
nUX5eldTRua+NX+QOHafdLVq2UEHBVuzWqZLpBVXeYwRcA4mHgPo/ScmOKVkreyuNqwrJux1xFrT
YTXyeLFP4Zl7y86g1zbiVeqJTYctG1MlfnlnXxBmZqt1M17uJXYkvaRx+ooavihbsrEaQFhzaMuE
aH6mDTUXicYtlhaXmuuhCGJ8Sf8FIWmJC2mCb7RCnVEV63f2ckJfTbgwDa+0BIB/gOe6egaoVz3J
KkaIUAiDM5OvQgZDt0I9Pz+dcEfqtL5qVIogX4h0gDWCInknC8rX4iCvLhPpQAVqqA4O2fzoReYY
xFLOREC1KunHfnbmMFU3pMxdiCCCpoN25g5Qr89DggMoTC+VmrlzU7f25opyDcP6CzjCSRnMEBRx
7oc9b/ir1QuiCCNB09+I4yzpD5GhWH2SWJeIAvAVi/BG/sg5W2PbeFnYGl7DAOTTfqtBZIUs3dqV
Hc32tC2ekGn3FnSBLzmRRE8+y2olkyA7P0gi7RE+Nro7qZPuVOvKVoMRuzLlKcQ+k/EDa6vDCKH2
JV8yZS9u7r52yK/DfmuoQkEj6tMf8jGAUgyj4acJ0osFacVda3fMcA4AyxIRMMpNCKavpo2vhSqg
xOpFQ5O6QgtudSoH6ufOM1rhPmCKx2ovnA/0qaKfSx4oTOOxaJlfW52zxVGcv/t3/VoNzkmpTuAu
tfcKfWvgaL5ht23kWJwrKsALWYTBLZqZpEFv2OEZXDD7zDyGdhKl0SQmJ57YjFpVHJEGKQLGi0I1
v5SU1a+9Uv517cOm8U4K/LcqVdNUGDivQjxufyMuz8m0JQ2IN62k8xWRViqknv1uZ3R6+5sHqPgZ
cxms9sKOHWGOYxZdXQOD9ieCnr5TOwoEbStfAOWo/oB8IilbaJGNtlO7s+k7StzOPUAEYonGg2am
4K+lxxYXgeAs7MHv/QrHsAh/1c5dDXvYZ92IvPd6lSp/zPiTY8dG1lxWxYAkqB7eZHiemECOvaED
XBBsLr1v0DmqzvJSD0XJW9HfPwCf6/ONTJlqkT/qAhiCxrPJysCgFVP8UE8uUDivSKuc5+7y33E7
heWl/ziJW7XRpG6dx+UvJVrxPg9NNxhwuZSzSjwuTmSJSzQl5eejpYpxpIIFYdmgcZvqjumnp7VJ
3iuAeX9gkxMR0HI45t2DhO2iwpPeA5x6m8hUuWyi4+7QEjAfifhaooBzq43lKAVCj2QmGkfmecyF
IfR0SdOzkmU8Wd4M1ntEYoNuiYmSOqziFo15+f8yOlfXkotbR4Kf7oheH6C0AX36Z5o++NgSCaD1
7aLmB59bERQnH7jc/I9SHANbFpkvMi/asJV0RuKfqcL7+M8afjIhyvsqisrPiS4qbUmzj7OSBEVP
YV45wDCTNxFjgmb3dVt103LgXG/CTXsnNB7dv0gpxIxBfcFkzV0QSBgYNK2rrsXwpATGPnCWbsE1
PHMjwG/mGFALF2/teN0rhQ+5WiqE8yjyBWJ+A/uX5VCodDbbmhdEIK56lDGQv+X1HqVcNXx1yVNd
QFnM2iadk6pyO7z8PaKsHJG3gpL2ntBUAtO+RxKsYSutNAYe7t7jd98LLxU7W3S9wOwDGY9SK4hs
giybQ0p42dWk4XSZBppHMeRv3jscxivubK4zQ7dx7Akr17uA0xfQI1qwuWUAEVf4YeaweBytdZKr
+igIFOHpiHkEkJC4rnw7+oeg1iK9MQIr9AJa3DIMzfNFVNuc4/Axeb4BkA76fjzLzz1COcQcybhx
53CBcNJ+CatADJxsEwRE4NK7pG5ogdKoSrfaVWMtsO3JcMDXmM1JEdZWvHYL09Jze5UYhSEiCKBy
GudZyRGOYZvnRovDAHhIx+hQdNiXvjEvI9P9/sMcMikJXlFAhSz/Ebm4JL+QoySZXiDsWi6s0+kX
WFHLcKJB6xBIonjjbVBQQ2JSbetr+bhcOJhxoIkc9LAd3v5n2lxxxMCXv+BskJ4WPab+07j0P+v4
4VakNIB4EmvjLXVXoAInFknlahkWhY96qW2v0/Y6mAis9sIaoL/HcBWse+xPLlCwb8TolJmQ4I+f
JAp4K3hhtekRgZdVTgrn/p/n/WyZMQ005PqdnQyKKsKtmbysoJcOSok7iSXzO9suYZ9cuEF34WpD
igt8nb5sNgKbrNmz4Bv4Qsb/Z9HluKcN5pYmRQBIRJ25/wAqi+JWCi25RPYKIF08W4eC0NCQQdEn
NQD/6pUnqL29HocPSXAIKWA+a71G4ybh6VhGUWo4Kq5isAhmiO1vuG1cn94/6InGekionpP48WFJ
wka4kV9mxG1qk071ZZLosbrlY4G9w0jZGE6dpqpKaWnr8v/UHPPZIJVEHngQ0nXM+m9ZDCUIf8XF
43SqHsM6r5yiNkk98VsTOVElmg3sUY7y6Ujp3pCdnCr/Wqvga+V853l8Ty5b2HVPizG2OvErMSdl
bSj5WAmgpmhXXOzAeO2P+fuUDcy8CJ4e3GeVd2UWMGJYXR1+2iW8TKbvHMwF7bUdmwcrBfVnFuZU
0wDMy/IAOsTtc7/i9bcUURqLwAgS2SQIHu9iev/vGnt/iDpRY9i8DUWaZ8pfvPsa3/E6q2DQ1W4O
M8ZFcFZfKlpsEiAoYJKMf1stD2XpKxB0rEQOdzO1nF7vDOtCnAass+Odwa0rHPjAU8zX7zRHXihI
Hps8tZY48rOfhIgKp/V5/XvgW5Wa7SeP7pbVOzh1UCRp59BjUi9Oa7zRG3kPlQv2Wh4LyRsDovTt
768v29VT/IAu7/+Bx0fr7g/oPfx2xFN7essmsdHs9Uls90oePXXa0y91cApn4jKoI8G/QX/A/rGP
thBrD21MGtWWUqxknmnUihX4ebCbcUIChxeRXEe4s6ea8eOWS6EFut24zlbmdcbcxpsLFYjQeq1M
crGfLJsSNxyKyv4VfBYo5XyORMmq2uSYHQQudyAjD7R8pXQGyxFbQlTThaG9eUYdbOo9p7gRKFxt
hRZbRfEt7Nlb6jTUjz3AcGb9O9ru9aXfRi85jiUfkbBBDMU//7sSCsUSiQkCshWt7sn8SXnyLUCe
6nqcTK0dK+gUSi5V2lVct3HaMAQolfWnbHw26ppaTro/GWFTQXueIiZYdiypgLddVDokOE4mFOOY
4mY3m2yOJQKZGaEy87ICOHk+yDdxqKYiioH0aeHJ5OItYpys3LwfOy5owfS+1VAsZxMaO5+WoQrR
KySrAay5oobY1/N4tkuwKaiNg7OzI5S73bpt7tlscAIzSVZGlaovxt3+7lm0VC72R/hAA67LZ8um
ho1L1yITRYKKUc8S28SrcQuWPdIzrUegsyKa7IcywF3FH/nGXxjGexS1TQVKKlm9K5qkzYMOccY5
kgelG2CEKTQen/tX9qVIzEFVlTOOfxWu+UAuMqxe6DuBswDI1QcgXUxkv4qwZz3h9caCen+lufnN
/JdHJrgpIjrl3eJal7RwTiQjdqUT7pBtTIo76bY5nVVboHTX608W8WHijWSKeonSvCx4PC4FyOcL
Q2Hwk0A5Fv98j7TPvFMCkcjc/GxBbpjC77NjIsZ/DyIpMG5cmcoqlsi4UC/FrBwEfTSmTl11H4TB
aKahi6rZBk+UyQrf5OUb2iHRUi8z525qnX+ldfhmIQ29DLMQFgoKjGHjtDedZK31EDcnivgZdR9j
FYTyrl8WwPdO8z/Nn+T1jKQypH19+mWd223/bw0Ml9KBrDRHUPsmMyTbe8rR4qKOhX47s0v7mim7
1nJo/XVY0RAgAYMqtYj+nKHlmpk3vOkDEEg3LTP87bs8WGduoveYo44ho8xZeq7Tq5fTboZ5ivr+
ID9UQVWfd4CHzydcz0pnrze2EeYuvBfZSOkyQz/peHvivCAPpjOV5+ArWgDSH9+8QLvVaf3UVq2+
H0Rl22MfEx+bIwUZlDNOA+FnHCnCGcVpeFaiyu/p6ieWX6RNt45b5Aw8AADetTrWtNcWpkxwMZde
tOsNI03l6Cjo+hhzbS23XEX121+JV5dw051KQ08PCS/FHAnON/hD8ihN4ggXLW8/442E/oIqaX5S
lVX3x8QasHpuNbtWrxFIPjcS8zEJPfTyOVK2orEr6J51MhO4N82Y84+v1yqFYGCPtrn2jqZEoPZW
gDy0eJpy26y+RkcCVmid1kZu9q8pAV8MdIxchYXmy469xGsK5pFU7G13E+vfnA0eCJezq+6QqODz
+xIVXkOaZ1aqRxs4OOQqeBWNEAzrLos7gzVzaNCyWyaymEnZ4JpWCeVoWcnZusCYQpF34i3brc7J
0AnC5FQKQFqBHedB4k8CrpjZpdIIciwbVZRxVUDgDawY/KQPO32YMK7M+9ZvY4jmNzRiu8iVgM69
cvUVcDMWvEOkGHR4JnKQhhlDS4fjim5+d25Vp7GCk3g8bQ385H6UwbCLdIQox2SaRYzusSP6dqdu
/EqNtS7VfzqtyCnHasxcj8y4Sl92qSc6nzY0PSUq5eI3V6dS566PzK/j2aIPSp+LyyS50txty7/H
F9amTncuqUaPDrj0JA0uCchdp9cVFGP0lCkBuz2S2HPKZO89UwLUbp4I2htW3SpzfyMda+BIyA8p
l0GdMFbrQAe6UAvYoDMr0221QQd19+yTJVkWDZFOdn99xHPAfKh25SULsDaVuZHTa1JWZ16izC80
AQRsUnxQyWrNz6lKFovdfmB/yNjz54liKEZgQ6a/wFaqXddvN5VWjmyREil3hMsx4BTnlseeCRJ8
vKNPh5snXN3wmtt+94PdTdbzJ2OhdYxWZPOjWqYw+en9h33vpeShZNv9rZYHXpgXnST24RUqTpoQ
IwsglQmJ7sbQUd63sdY4W3Q1v7ZGoGgyKzuywd6nX+bUi6somLFvCim3MjqGwzHcQcVhRHi8Kyaf
4IlVMv1zJoHEPAfiuFvGleUkX7cikc0/FjGVl8M5erHnKC6pz7VwpbdCmis2UWaaD6wcQOnLQ7JS
xBzGCfh+RwqqiREC7ynQpUYxf/QuF6on44iAsk0B3VpetDzm3MRHLbOtYNYTeekwTTlWzGAEelnG
gP/0GmvcvHaRrMyo+6LAM+JyqqdIHXyNDFAKvkVD6dtOe5/v+kQUaDu9Kc/5hDNGj3ZeVi8nEsha
uO2QyRlKyx3rHUBqR7pJI6guzfq6j9qfSjFdvrGv75NDhhKCCcnnhd1p10XLcWhLIQt9grZSb+yK
C+A53rOD/Ju3pS2i99JO1WW8AOagGpTF5FkJWK77JHZIyLnR5e/4e3Oiu/K50q0nzhHNjj05NJhM
dCq5OSDCOxE8oLIBkL7wltPIR/asUJg4osZo5Cp60F7D8HM4wdU962QtC97revV6A3CM/9gHQMST
+C5pkI45UY9+7or1/dnvk4Ldtn7SpjEg/73WozgvMpQZTplne1BSZaglibrjIUgz+ltYM2mh+uqv
0mF1j7T9N0d5ffBidiFYQ2y2H3ift2QBvtQXUPxYohXkYabTSTwJoY1/ldSEW6nbl+wzybW1XFsM
HngSdEM417QSrXfuFAO0VeIDlrVUr/zED2VMQyXr33dLYszLAnZae9peczb03uesuv8pJFzNcAK5
o6ibBd2iwc+5s8Tc5mitwFGvnnArw7tPDdtIOb5ESpe3SjxB7BSgysixD8mEEu2/CX2OlWFSnCcS
DIP4j1kAAJGdcEnwQZufrGKoh0y8h4CVW81t8/4sThTEgxzC6wEHaZzU4u8eZHZxORfHxbcPMczv
8uuOf7OAmn2h84enjb64KExqmm0kQYe3UBP5gvJpkt/MzD4EQQ1PB0xy+ujAb8+40MMzGwjISa/j
rvxliBzw5qLSPlHZe+Pfk4TnntAu3pJYUUQbIj6wYsi9ZLTuWSLbEjVfnp4WurI7XZSn15UPwpm5
5w4zI5khYg5uoI0xyp5Ci7rNOIBbdFqPXk8n9UlPupn2C7zPw+pdg1Qjf/aO1mIXJth6jay53a5k
f4XTMjd5Zfv160+VZw5fqFhx8J53WKnJRL2IrHQjeG4ZYhl0E30YhubzkwvO/AydWmrytdaxhwOy
Iy0vmL9KtLprLStUt12PU3NmLT9azqEfvL+WNAdLMBuAgPQdHp+GqJjdi97sW2ch8EYOJX7B0UuQ
Mdh5GjGJtt3FMxwIScPaw1TaDyJnMcBzwXCvmX21c6YZEly70ohu7mMy/yKegxImM2DsBaf4Ushk
pKU+3csvvGCT7I/fVXAmHNSQzUi4luyEd0y93nxs7ga6IBVfsEVkPtHuVbYUArYUtiZAXw5CJboj
0qBeO21TBDbb7EdJ5veDecVQOcDAOAwyjK4lWvmOCWq+CYH3juZPKhkVM224cW+QM5h5rjO/B6Pz
SF/UvxylJgSq4VI6CMHBI+thMBJvKK0i16XSvgIy5TDX6o7cDW+2HN5tMa52nTbcqfVTTvsB6ISD
cpdQ7FBRxe1Dz4MfYs9tlk+j8WIG1nXsMoFCTgdLVuV1QG4J+h6NY/HhLFSCQbvipLNikBcvocJF
w4T5uHh+Y7mIxj3sxo0L0yJHU/twRIXtAcUI575DQEdmaAX11OeM+dwvCqGp8CQQQfGnor907poD
f3odFDA5Nu0NNgn470gWxJaB4JnPTOmOkvVYlN2sLloRt22j8dB9MrQTz0Uc24MVikRg5gUq8BcS
GkEwSPJHDpaxDZEHZNeKsx3ime7njL+kOX3sOnrhweJXKf9x7/8x0YK6CqCh216LY8pkAn1VxLH6
i8gGysqGfUfqOmmQYKQWGgKvs7cHHLbzpkUVMRuN83HXy90hD3vjzsp2cQsllOZ4LqUgwqOyjnSu
ybFvFFBykkjS8x02VuJdzxwNv/pJsVc4byK7b+MEM8UjuG3H2kheLvrYFZ4an6Q8K8Iz6NV3QIAu
nlEtXXcNSnOhKnVQEt22cCuLgUjWjaP7VCWS6Vg3w86FAkTh5EVucj4in04kheqyFZ1y6AQdAI+d
zwGzNSwJ5qsjYZQcmXhPLR4YOLAfwj6Q6QKNST217Nl0odrkXwB5aDmY5WQxDamQBwvd1+4R34SH
6rOKuVfSphVaQaKDML1B/d8IRiIlebJD4M6DtCRz1WK9McfGhEGAU6Jx8FgE/MDvRp072cI+uprI
g+VUwNZy9+JEw7uGVSoN1UaAwqfasA/H1X8YKierhY0GK1fj5EF3xrwdksLjGoW34I8OowUMYyvk
A84LrGcW5ugYWgEHrY7AAg8jHm5q6q/fGiBixqp6IN1FkRCtMmjLq9m7BpKORT9d4AmBL97LqvBo
aMQcaaY9Zwa8wfDAb24d8TEQ/mR6QE3ZXOUDvjLwzmeuqEe/0yGh4h5KBJATISX3Ua3JRPRbklET
u3mlx1VGl4RXUeBye0g4AbXzm+xp+Y/Sh4smN3Kier1gvRU1FTp1kt1hdPPYnl5XdJmxGKiIlR9A
daiI4+D25dfeSEJO4h5W1SZ27ho0YV+wtvVwT1WMzRthRcnQ2uPsxQD8rgXnD1RgOUrUTUUy1J4s
4+Ms5YC7ixXVyIjobMSzBzZuZXnOP0HX2LjtkFsl9BnqeVoX0DDtVZsniVI3E3ZiVfqFYmNPV2Yc
BIHZbtOfPd4l5yGKCyn5es5mq8bnJGTyA5XZgnvt7uemH2eKCKjZnoZFRQME+QHN9P9PnEBtzieM
39bHBXUFuET+Xx4mTc6he3lQVsOsiAsIu7AfJHcditIc13ea1IYIvd8Ezah0sdVOh/SnXk2kosQY
3MdDsuZ8vNKSEP8KsLrYOvoCCs/YvnNujU+n8u4Yn+HgOfc3C83clRipUErEgMEBbfYkgwre0dXu
BNn3My2qiX+ABX9T/N6CWBKm6MXdfcikde0BVkRsGIV5o49j6fpHajXxRUvaF2/pRde6EBin/r5t
GmclyXt+m+4uuChplWqPApC1pwwf8jm2ljidhfdGibX6X5KTt2jNJ7criqnRsn1T/lFS634GUJMi
b6Cv8XI2P/WORrJkXIOJEDfoHatF1s6RjpQJ1sl0M96dI7Wk2E7E+kyzpLQ2OnLDjETw8gVl6KHH
/r04/ogrQh2BFZkTIEA+xMEIEm6rWB1ng2NHfbwLUEyeKD6057ESH0FK0o0mCr1yJubUuOT7ybG8
5p8LPOPynvvOXPQ6SW4SrSj4U/hYqBL37eG1LrHj7nl9EGC30Yphu+lmddVwTz1IIldSl+TEWgoI
SqbLjwoAxiOHsPHWpqYEM/Eq4nIf+kfPKeCdbVV7YYS6Pv4SJgGGviU+3iF4Z3uhgZ55J55UJJbm
5/1ug6Hu6VOZ70PYIaJdi/cQ6NA0/nLzmgcaNwrpES+UqYYnSRNY9+ydK+OZbyF0ARAG7Qoqmhkg
ic+ByutAm3EmWp1dT6GhVAuj6m/XV1PUqQnET4yd8VNzX/1cMaBx8vxYYJQclFSSXt686ICrXk6x
wATQyYZLRpU1tVAx5LxkkgrL69OQdtBNIx07oOy2wAjiBvCsxBFvE4qa0Gh/3jTL3MhUlsm1SBI9
t3/483cg2puKQIqK2iDTpqV7OsoR0cpKZcGe1tIjdvxE15fdor3TdAHwtpyKK3Fl3A/UgSzw8JVA
4nQLajKxFWamYyoTXY4CqBYsUNEt7gR3QTE4tfCluoLgt1CUmmO4Gd9Zcca42af+p3GkfhOUG+71
k9GW9I6jE7GLAFekFcsbVhlnv5245Nym6hoMaM9HCqp6XIAXv8VFumB5YBvRiEVvPrOvjA1CiOY5
f5zIM6GpyyjD31/gU7+g29r7539TnK+i3HtX5WpXm3Da8E6+chwQkhU+Ca+VWiwDnJh7rnpYGo1W
yY52p6AzyyZ3Vo/VWXV4r4eTwXMdxzyHaLpnRyDkU1p1gcZ/HmlFcN1dNyGjNxew2ptj6UcO/76B
bvyNoAAAOWDv5Ls17m0BTVGTv5yWCsJsm8zeV3sYAwayzJvfItAKC0hauVdMn/E3lGr+SDjxtDC8
9Vi/1+Olk5X0NZU460E9vJt2Iz8uJNqa5cggrCBHjq92sdCn77cHvPGGwXaou/p3RpTOiB6Ohd7t
3CmPUILZ6lPhwoNfEUkQRT5+sb7vFbIK05kt0bBzyqHBk6mhxGM/8DVfnUOoIQw3VOeUirz2nu1v
LN4LFMXuK1VYG5yYw2ZEPs4cFQ43H0O8dBeL33s+dcEkSlwGJf1TKTo8oFMuaGqBmgxvXnLR3y6/
3LGT2vzokO9ZGAPSf6qFVpDvCMv6Sqr2ZOyiksAsX1coX+EJ8ZmrGothzgoyaMlqTmwebgefSMqU
mbwyy13PypVwzDUEqaWpSQsA16CIQdPP/ltOJiyNzJq7BTdARvoZpdeitf7W45T0A/gPqbmOvfSe
16Rbi22GJpExc1e4uNVVfnl9BAMoX3psq7D9P6yUmCfwGTJgx27KSQ6i5JY8GElrNhlTxEGbrQ8N
nawObckvUOZWlQ9J7iTqZnqj37TmAqBEGWzB6FBlheVs5GGBbXK/SrLgQPj+aogvvYtCPfxODFey
VQrHYwDb4PRIb0m3u5EVZKBQhV/WTchaFhaW25TsRvAPHmtUa3BWHMeJH0IQMRQxoPxOoqsLh7Jv
wflTHdUGnQvaWsWasisERm+HKARPd4j1oM+xwIoII+3wNOtc1h7aZsOVHKLoouPh64mE1Lam7dn3
2PKEa+P/V5F8a/hr9RlGu/2Ljmo/fWzOcI52GGFftEhn8Fq6FNdaco5ERHvgSZRHmlfu0ghzKn28
ztvIvI8dfbwrs3EiuQsgZkR90YqPwNmRQJXJU+fDopQPniwdroEzFSG/nww9e9kbzF93FF5qSbO5
NrYF/qE89ItM98+67PBLy9aNpOT+HvNt8kbGgZbXj0hv18ENPEz4bsWFBFEFgM2jVvN7RGRsuxIG
FY2rilsQMKGw3PA1lmXzghnDCuQAmbUglYHUzWEbIAROoycz4d27ShmKNvlYIV/oYph3h4nJCOlj
YTi8o/9ftCr/gtnLgBWbpJfDR0s33Dvt6aP/WCWQnXzgy8MTMLEaDcGbInFUryb4EVaUvweve52D
zsLvf8eCJL+o5z+PhSehWkGiML9+KAo8URzGGwQn93AJpVOLEaTlJX2277byhafvr9MEByBLJ8ks
Jrus4ZTjB0/uHrWNNagYewqFf4cuVu/X63F37GZZC5RHTQAtFA4Jbb4HXLHL4ompQJ02PPB68js3
5tBpS3a8RP1fahvy8Frw6Zy0bks8Galwtc+lN3UEuD3fE4fISlHS0W0dq7EcQxJjqb8vHrylk65O
RcL9KQMXUQxMYrf8IogjFd+wU04Rsbqqd7midMw109WDaMouhYKiqMCB8N8u4a1px6sWp4b18RAY
kissGEPkWQr0V3nMnVO/7wyeGL8W7zqd/lCg4zmVGnlImCY+Ks6y9NhqHjmVZ6E5mm8d21KA+HH9
pT5LJ1nQ4lhPBeUlWcEYtrUWFTuM8v5MzL1MVZhqD6rjzzyoGh9lymtSP/rlsURwrcAuu9YAJ7Bb
Jx63wKGSR3oZa9XrTf243I1vFE28gCSR7GRq3Vns3Gb+cUUTs47XInQb92CqBiIRiKS53zeOGD8c
M0iiWVjoePWeKGItawvVa0K2zHn92XYdD78iys2wwV5G1oIh8PJJPeHwuvUbPUrTvEfc4x9mt+W1
7inC5dwqh9/T1z1WE30JMscP6B64FMJSlDrV5sPe3VW9lC2YqDcYpCXs18rxLl278+I+M9dLHA4Y
eO9IxcsnUqGZ771T1CLdQPAL3m8mconxbaEfVD6k+VpKegJn4g/SIqIiRJy3keew2crRVanRFJna
Nx0IFwa/hz2E7ep2cHKdHjsrdUqI/vFfW7/AA0baa9pkPlZTPiUzEYwgMUZ73bFIwxa7gel6d0K8
qmcYJJRUE825os2qsxZIPmgHOqgRs7m8ADyZwy1TcpczmoECfr7j9IuSbbPFV200hDtWy53+OvpT
3Ze+MLKb5R7esgFqoTJCzbGK6syOB1tzDS779DEXlbaVK/xIIZyQdZOX/0pcijFUczvmBSU8ko1S
kNd9nPQ3rHgUaOaGZsud4oPk1aI1O3HrpUgx3hnrRUgX8dB/IPMKfKed7thZ43ezemWCQrRFYKZB
ea4UoPc6Nfe1KIzkUlJfdqT4CZFi2Hb7UsO3k84hx+RVP4+7zbbb4mJDY70MDTuFsNqKDn2MQsA/
JMwZXJuWFKyAOYcC15kj2HvIcFIo/nh285mbWAllNS0bcM5bNar5Ldc2SurziiL03dywYRWcPqzw
BHmkXuQXzsHuHLOvmMa/eMK5sv6y0azAfzerwbGZOWK/Z9PVvIacdqHZJbFoTKocpHLDwAoAUGOC
t9+YVg7Aj4Lr318DnGegukCym1odwdhGWWrc2dojMoILCBtLEOUQk2sT4CSbsZd9dZpkIvIRNBDJ
rZ6nfEvuorbMsuICx7RoeKdtaRh6HQLWhmPB+yLxc6WnITjV2xxkKCcE8WRO3a7CEaPD3VEeL85z
GC2eY5Ta/MXRLoBWFnZ0rHjS6FpC6u4jDXsAz+KGLxRVXLBYqJnl5tDC/lVk5cX8XlrddTrSzfly
8pv4K4RHf1bpfadsXzqJOw9gII3ggJ/bMITjOVKGKp6WQIjSgwUqpo7eeTNDTEQTFoJqyw9h3GQS
xsIR6WzsLRMVp/dXjd+sGZ8DQ0lVVl+sZM1WIHqIksI+EEd1yjZqmA/PUPSo2GYHOnDAM69bexXB
PZMmw8VRU/Y91WLoglAehEXZY202fmcR4jLUtQ+M1Qf1DZUU6u8fXGSmmCIHJrbFwYyGjqfN6Gso
T/Lk4xRWkIpEwlhLdy6BhOmiSX/8E0UlLbDeL0aNq5m9v4/+9+/FKA/ziYLH78/d3eTlPYuIgqO7
Wcr6a6+OKmgQh+QjOYDyq8F2aJdcsBGlKfbOAeafD6z3cYhIDFMi/yanT746Q7Fpg9sy5dYXusnI
bmx+ilIhurWIiTJbsapcd8ypUu6np4uEj5IcC8ebhf6NPstd5PnNv6q1b0CeHl+IVYZZQ1OOKCMD
cL1OufmYVXEb4XHwl9zQCzu/Mm8epKEEdiH81LMHHEwvzkWp1Lg10xCMpMmpGwO6X9dkYjZVrRVP
xYMMT2D0sr1CiItbtJjfAucv9TsI7IVvy8FOfVPIfSbJDopfAIZoUeFaa7EJn3jjYS0muCBL1INU
V6mTsHd/atxymveNflD9Qlb6ufzEc1aYyn3ngww1bfna4ObMokgXDGk6ATWnKLASRmzaWPhc9Qx1
U9G2R/Rr2CbC73ss7yFlCEC5k/AyPTw4Zy/SA74mUVdh/UTK/EWEsm3DWvrDUIly5jl8l6bber68
QCNK8aTSPyfJLL2byWopOdYWbbHofgIysw/QzUilk7wH6uaF40GtQcSfZQnQLeTSwSdA83zsddfu
7pdQrkTJnHqapEM8fTfsQB2bWEGPQok8jqFOF1BAlVIleoft/ie55+hWPCt6ywhFPNrPwvepF4CA
aoEnBk5ydOa2mKqCBxZMg23eaOtf6d+NwgJmr3lj64b0oO/1JfOYy6/hqe6lK2BV71j2gVtWaFin
/z623U9817EL4o/2K8GTHg4pRxL67RvksnuHeJ8jf3sAi5jldAdnylba671Rt3NLeQxPfKCjyFr/
3Wh0vngCDskBZ5cvXPlgcT+Utb7AKG3Y86mU/w/0KZ5jWqppCrNgMgiexHyDhWP0SkTgH+IEpQX1
h6K6MCazk6CgQn7QgZFPNZWjZRr/vlk0VAzt1TLEzq0B3ciXPxTgcU9NS8v8wREpulABhuFw6eNv
E5sJsI3ldf7LhcTjPmHoKEVRl755pVZw78qF+apJ4Hyy3HKTUGImgnXcyVUWA1THtmqezAq0+YMh
Q142hXy3Sx1I8GZsod40nJUPgg/lzwoDl459fo0gzZkK9Tu/DC33PvKt7oPN55dWO25CYEJdhXI+
f/598/MNthbHt4Syo8gRre3mv2FtXZ9E/I9c2xPDVdxx4EDzLEm7BPO1ugfPlSALlyeutsaC5hMs
6dAULZYBiEsIPCJFb2g8W1dDddAVa1BDdc0UllLMdcNxoqQpn7bnRzT5p/h7jbrEg5sLdK5vrXm1
raXcZurh7yhfQTXaGF/ilYGOy0hNZuw2n7hNQrxoAArIaG+Yn1JEGM1lM7H1w4n7/gBYklD2D2N+
U23XQLgdbgo9kxlKIlUoS67GANfNcQPSej8snR4pgvFqT2PYSqPYj4Rz9Tk0+x5wY7wrjVJO3Coq
zW+iTnSktb9XlSrgqkL3OPPAJryBdDvPXHLeBzUIv0aZMdwTO06/Agl0w/eDaWIcY9joel9AbhIt
aLsaNyeJF4a0c4v/M5QO0YWn8d2h4N7Caaz/YKlW4iyxyIQyxeYv2mA/ka2EE5MWqpF4msklB8sT
IbsS5As7ZoaoK973aoPvsed4MPyAiki70zBkUEy0rWL3Nt/XrbvGKkmQb58AbXsKDI6f5HlQ5nSq
8lWkpfZt1/jg2S9/P2bICn2xRt7v2vXITfYHTtHWyrgWd7CNHQPof3e9yZCdh0LGS2Gq6MVlCWu+
jT96BBXwgLq8w1oKQbL+kmcS80rsSDUxBC23lePdsSIEhLK2JaBqVI8VhBnuJ3fns9rO3k2Agqyg
ktp1W1oS5gksg2PZx4r9ealNtgCCICpsK0sftHXqAi5D9FLQKEutqdU0Ox+jL+JRYZcQDTrNbFUU
fQVfr5wITeyHYH/dRp9T/f2ReMLf8INmifwCvYMsWBUpbiMWneOzCD9o+9Hap9uImwTWpKx4nqxA
k6cCeVKai2YWwO+DKtX20axcB9khEEDtBsM33X8qePmrNHvPKHxRUOY0maO3JIZSkj7613fsM5Zo
ID6Imhn6rY7xSJHlrNDukrqgVYne8DqiA0Nhjoba4KW9VcAlX6Ack1lD5m8n0/71QhtvLhkUN6Js
kQ8D13YEznR+xCI8vS3YMYnbcVHEsgYs4AM4O8t5dirGPaJLJbmYpMXZ+IszMnwXdU86m4O098Ik
7Mv/00r9lb0IW/xernnah+9+mWn/Mk//kcmVt4ddAC66X0//V7HVEgN5nJLJj6pillkmtJIxzDNZ
OGKNuZ13zkzYR4cu7d4MscOYHfiX3hLbfXUNxXvkc92CjZ8zzDaYx+D54VZidVkhEvC2Y+34HgSt
zY0IR9tVdNAcsWD/hjKFhuDD2wreCpkerWlKBIPctxrhX6zd1d2/E2ltLkVwNavO2ApnJbymdvqw
R7ESs8Q47Pi2EkWRY/MMgsVajzjkyFPRPwV+9R7gfPTSg+lIHZCDm0OV/N+DFupqIREoOnC8bfmf
LJc8gOZ6ADrRidDsgiGgMRVcNBfUMwOgoJBnQgMIykKp0ZQYz+QwSEW4JSw9s0siB3/pxg+wykOK
RUdnTs/pSgMNq/Wv+g2LNd0F1IOaLWfcf5Y7mKaHmeaZoEeHi/EAkrmKGiXSVrgauPNgaubtT96+
EzhuAlDuJz3B8mbbipEysLFJf9YGpqYuOSNuLJnZSIhFE4ooMQkGW0rA02Eq4REHGjylpGufcAo4
te0qayEk8PqSU1zbQ1I2zyQ0v3iCKtdslaFfHRwO5jQm+93K+xI2oyI7U4hV5I1ZRSGvQgk66Hmc
r4QXtH36NOdxct7vK9jLz1DlrzVzDcr1bulYx/37Zn+Zh72wR7jVvjKRtCIDDjWHDxTXN/cy1GFp
/UPgz9Hk8cHQJmLUEPqj4t+8/F5V5lWQCvdhiJBVw05prnE9ziyEMylSTZKNMnpCKUwE9DdyiU9G
ffu0Wf6feMLlwXHbukeoo01Yn0miqWfNeF78AXw1UMcJeICBnXRGLvC2aWHVp4rWyHmB4oFf8f0K
3P1BQDncsvGQRO1+4oc7m8oKDDuG/DxiOzQIPplDc2oEo3FzindfaASSKqoB0mNS/AzFJgiPV9Oy
BW0uTgdgM3G9mS4CowNJHxwu9gbty+9AwK1hVkjqcHm8Ogm4Vw2sDeqV2JAygJP3tkdL1S9meJJI
7GgfYL1UhBgJAAV95H9K2w68vzVmAkLiqtSRy/z0Ll5DdVDFww7BywyymwizAUDW1kfAputirT2T
j5cLPp9C0hyclJ/kiAr1glQx8ntyZ2fWWijhp2E9nQ3ebMh7tx2rYriyJVgMAppLRWaxJqbCvCXc
YrKYUTxzOJ1u9+jZu6AEO5PP6NQBElJ1d67Rb3Yl4vhfBn2fXZ4OF2BLGdSjIDzTvC8Dvs1JZ87K
qPf1nqc9AKY1zcONFaeqFsjP5AxpD5rVh4UjIE3KB40s3EhfdP2OPnkiVhqFxvolq2gWIg4BjAS0
f7F7MgMpub2WUWdoIKJAhO7oDfMWfdLt83sVtlUfb+PkVJYSXM/KaQjWIuHkbVqfVU+2koyzwHYf
1mFTiJVp7ysry6y9op/5rFhh24HQ3RY2t1w9AI9kzLTmCN9Z8Gk2HhwVpMZaFEcUoytZXcU3B1jw
/dqXD/XnC2IlfUODV8uplxtnaT5J/v9XbulBImBPJgsYSTFQvNjFbbsiN2hZXnJX+rtdY1K/+B3R
wSqPKS6FZVZdlwPXBLBcFXQb5Sekq3E0VmcCV34P7eN4B+R5HH+p1m06sD/5vBydGBMW1QPhYItu
57JR6DlXtp4wz9lrshFcP6MiWtLNT6HDVPYn+q6lZsv5qVd8w7Hy8doZYtUDnIlYm7iv6TFuEeW5
xMM3rLlREzMzMkO2q5iNlJNrgpW5Do07o1k/IY+yQ0+5bnn8KYFKlhwB4I79hlIfEB+EgO8L7R01
O8rcgFV4sf8HkWA5MIkt4XlWpYgBkjgPXRAGqpga3bhk10VDoGOxA79LK2sOHMukbX3NJ6iSfapK
6+vAeR2HMw0jmm2z7lSrguFohxi0kDG7USJF0RHatJ+8xuIZbbolo8zZTD8xDmKqK/1KqOAmdxoF
f4F+BPf6Bla1evRe79MJYA95uEmFwduqTEy5ygo38s4RCLBgggbrwW7jvNvrB5v3/ie11a1XfIGM
zMCODLfUQk/whY2gSJTJOGbUqe0nW4sld7XYXlbqanykBOMLPN5JjJ7BuefQ1rfztGbWZn2+G9DT
8vL1hygUlJ+F1xuP794wXrYtOIYrY9Qqrx4VGXvxdqE572h3TXpu+lhEZmtU2ZxG8xATLFCGEXI9
1VUY5yEq4FZBemfijrRvxSxLGXQlxKuTXuEbt2xtbTDIpsOnQdGRJFfXgl/pvqRHUB+RauyKd9G+
+zL0nkcy82NgddbdMvyA5RCcgJJSqsRoloqwdVxQ0DrW68bSTpDHKNw6PfBNqP7WclUNHl66oRCq
lRHB/PgK0XRh3ea3wkP2xHnf9qGQFGKsdt0xNSIvcT928t64dpGMiffO2J5LuM6i3cAJD9K5IcYr
HHCzRnhfsR0L6CGQtfc1MOPtv7iV4ASO6X+m5reksvh0DxH7iiubtBjom1SnXOcm4kFRAbGOz6zc
VG8R/bTPadiCBqstoX/XmEVJwI1Zoy1azmqsO2sWRklHWMwvz26uqHmOb90fozmIsbGCjomRZzJd
tEhRI2zeG1iyL0za2G9qb56tHTW3ztu7bKtc2ONupQRK8t6zAlgatngZVZGgw0G9w187Hn6QlPU0
shi2pZX0mKTEraXYC6BVzqlmRSOeJCh5SCtDBU6Wp+mZ9PLF73pOi2/3PKN9rgdwYC+U8gRviMtL
IDJasCUku/lE5xwTMIYpXtpNmvHznGwNicZj3YHT+UVtto4NoXuJa241vQKIzCosXu1qjR+GSgTe
IbCPp3OXddiIDWDmUm6hiJ0LvRpVKI1KZq4lO+9SgN+OeFDaGUKrj0KDjhLwFmDhuGlcHJbSnIZr
LTuUFqf+Klw1kjW871/1D0RDloy83Wl7kOd0sKn+YG3v9ErQGrgnOj1W6cyZXekvcLP+I5r9+vsr
0g/J5QPG9kfnP0YDSb+SLMevnLIDIzu/60HkDwOU3xOqLEMJPVTSHa8QP98TKbLLknd2cGmFjuve
V71vUrp4ueT1YJlTOcGk1C1pIRDaezAkpzrqoGGObQY/EpD/hqci+j4byMsZ6GUO9x0zt4GiG6GC
3PHfPitiBBpuMRvqk0VK4EkpWfJztX4XB7cSnw7BUvIBpYFPU8JC6oMMi9Q0QyUO5aEp6nWklfL2
eJ7XcBPzs2EVn/PaojCxwLVDVMaSneQo5QcbhnT6hWXPojzpNLaa8tBdLty88toQAG8oaoR+12R9
eo6yfvfTPNkWmj6dW53nniWIIUZYRuEsEeRljNfWy3jUQ83f6W/QSF6lwuDUk+kzgRstcpVafkOX
rvmQUeejMOtNpRSogIMUoFZM1ez3HgDEBkls/gEL9Ve4P/hz9ksIm1Kzp8LQLxakUYH3eOewY/NH
XXl7ZsYSkNw7nu4YM2smqDgBemhTHVSoagGDOQdarrinyMjYyzszYSK50g9u8nrSriyaoRhorEIt
R+IhsDypVMGHc24YKsT7iFdnaxQwmTuInGQjtSrhlwnBlVVsFH99R+xQmUvvcwFyDZUQr6SxMEN2
VS5yiYa3eudTeygEcIbDW2E8jBcJTeOpFJv+X94HCLy1x318M6dXD0lq0r7XdRrlvJA3yG+NyTwz
bwxruyoQiCh1L2xZw4TZaImmIqBlXxHE6f5MKLrsNeG9Y0pJ+YGzwnE1Nj7LK0rn+uMTi/TmUofk
bpQpCqZGJirVMs8MNFBYbnqwP1xKOhqyZI59YNNrgMM3+Ge1LirKkOJPZkgLKxehSVqNsGrlioKc
HNq9hzqhiUzNm8vL79N7srqSy+24LKbWMYMlsirRmPrWeOD68/mRDYfzVOLNOnbZkFoc5nRfWBAj
ZlV1WvD99fJ1N/JAxkRZLP3EV1QJgpuZ1dAaxXxfXr2FAJ0l0EfXPXDAQLGYXYOFVzPGfX2VPlbU
qNnqqPkMvgL22M0VaaXDjoZVq8BxUmPJoA2UfpFORwMPxpFWHRQjTOigKD/46Ae6lmTdz9ayRCzH
BHjwJEao8BdXnr3hWX5T/dV4aJhiH+THb3jOoYaKx4A0rF5+sO4mNwD3RdkAwLqT/E7Z6jC6N0xL
xjDJT58fdvgDy0KVedknzZdps4JnI6TkF8pz33LR1PGQggCKXtPDGFLoPKEm+cvLEGmfAUxhQT/q
50ukOJ7/MTBkYv0ozRe/cpKoa8FLnXN8AKmvfNWu11WPcYQnDm6SwliCHpu85nMNtgbspJIeRFUx
fabx9/FIQXx7aNKfCv85/0AKNyfUHlUic54xq/yMIvs1Sj669Y4YDVs702N/EsR0Q/yatCR+Gfc6
MG2Nb1a0j3/Ru19/Z2Uj4QssX1CjyR01IbKuqv79oFb+qi/HSJgcih70YRsxB2WkaftDhYTuyz9k
d9SVgAgZ7d7sLffQIzKb5eanyQVeWl6VndOh6Pm8HBYrzTI/6e9jKCfihp/UBEqAEmAODnvpH1Zc
+R9Xlyz4yvWCwlRi8aJN3WXA/7mROxWUlfmZwHPKFQA83JCg6n7gkDFMQ2dPnAZ9alBu90pMZyzS
I2S0JczatZEI1lKVe7vziWgmKzbrFiVJumNfyTsMW4cDNG2i2lmJNQYZhgrg9TqehQ4lHq9n+Be3
plFSjqY7po3+10u53ueWlSyaCltwadfccs+g00TcaRkr7aFZz+pZ+5DlMeZJVbzRetUl9QpZlu9Q
aj2OqYhpG2NoZ7BTHofiFL0j77RsmHnFfyDjc4ay61P2/11Q97UuOXOy0TucxvbeIFJlRpsKwnXh
4wqFck/gfVFZwQMbXQYo7P2r++oxScpHSGBfsh/J6AVmcnB7oRf1vre+XrzEfoHKPnTdegJHkfJZ
cWwzpP3YtN+VTbyb3fIBs47r2nMlu3lkM1Se1JrXhb/FqZCMJegaLi+qsnm2pqRBbm/CDSEeJQ1q
mDOVWnxcLAiY1ctqZbit6JgYCX5xNLvKpsrxtsbUx0vY/e+e5RKT741Cld8TXZ92ekstMTNezlEb
uG1MS3V5Ydbn2CliXL0Ty1T2OII4PFPBJqpcuJt/BeUG+6ecM+I1ZOYY8JVynfqrThNu5WUdA4Nr
W7zHGzynPy1UYdCi1vf4R1hLLBrOTVlZxfLuBV8UI87fwG/yUabLeqilzbwUtsL/i1iytmC2Mcl2
ugS+kviXM2m2wdVhorgG5rmlzTkq9HXflywdobVhdBU2V4fx3GH5eJRvXufkSUikvoNjrSmOAM5x
A+DO9+zhziR+PTt6/NBIGb5xlrUn03po1X6ld3BxrcGtTtP71xHYPNe0OMef8Ne7kJyRQD0LN39i
pjp7R0Kh50Pa/W8D2e2JCQr+zl/VVT5LsFvEJZ6IM88/BuftmD0uRmMqUz59mjDH8utq9iRh77Mc
NBIgqg7yZBb5smN5lgaNhINCF6oXoWicfGuAAfwmM7JdLpGpWsN2d1oOIcWIju3iy1Xw9huUAZAb
qZmadYPfXV5pGnGr9903tL4CFQkdNh/WVIxiMbRDZrw6BWfHARY9Fe5sKio+lV0tHCq5ahLO7ZoL
W9xiZczH3bor4bdCmwf2JwXaNLjWZtWZA4q5o3xoA5ARS9BfKTRbzkB1vk3+4joNQGUotfsr+1DV
OT2QP05zwTjl3ZjoWrs9re61Kw0lSaBeVHsjD5W5LLXv4VCNUeHT4SQGoSoQ7fWMxn/ZTb4Bae+Q
vCjYVmP5qhoXxCieHLhgRufnCG8ZTDj3Tb4OYU38j1MH1Tveu4W82FJyI07kSvOFuqQqUH9dL28/
YMwcDS0uMFiC4gqqMWmxNmMAijsQ+e0m52smvQ+La3FMMx5yHwTFF1Ngq6FkbNAx8IIZW03Qq1Nh
II13altlj2Pq7djEBDhwrwup6FAk3AtktKCUMG7eZub3ngdPyNeV00cAz9TFdvh1VdzRtv3Nwasx
XyfgB23Y7Bk2sr/305rzdBpMbnJS5BhGTeSRHKLA8HaoUNRKuV/l4CV3/87N+5lxvrBzIEJzpihy
EvVGP2dXO7NXSu5Z7ZtKIMbmvkS9ED0XLvMVAx1aTRddaMJDz8lhjzkdFLrBMSgY8Trtkd4yVBgi
hlKEU3dyGedAtUei9j/Cx04Uu2rkHaAJyVdU858nIfy+4rrW6zXVRXbEg6PfC90vDl+OBk1+6ANS
bXDuCm66HBPc+x9qWnX2rSIXNGYlpTykk9OZtsIPfT5h7Aq93tdrfaZboAJxi7XOfi2NY5bHVG7R
eSTyr8KfXEixIutWPybj0waze5gMQpLsODWw3SB6CzwPI/j9oX5Bg+W764mbBGOh5Icxjo4s5vO7
dBy7VxoSUhNMcSiMcRhStaeQDFmzLVbVp9XsWyNxndSjJlDFbYzSHNtTasysR3EYV4AFqF1FREj6
+Y3QxYgO0hnXih0qrDZEJDelXds7djpu+hqDZd+l9Ky3n2Az0QQ1JBULsXaVkCjgUVqGgYgvnjg4
EtvyiQV+sxaVRmjC4DnpGiAAv+Q92aqE15U0IpvhupnbLNvj7pG/Ikl5Y2NWsKlwdFboBRtNeDWh
ODqyOfp/zcVJNCStn6ajzhuPmGkMRuwMcAVxKczaQrYbtE5A1h4/Vuy81sZuaQ7Qs5pwLB4TVCgh
wuB3rILkJ2kgWqzanvV89W+mtzmM/49AbdtNaBq5D+U5CU3izQKQP3SGWMg7EibgMFAfKUXSSukX
1qVunf3jjIiR+1Ybuh5XzepbQe/SeiSzFxbQts09lPSJg/EZmuyxWn0DwPbe+xMKBpWekHQHhZD0
yXfglT4GHLTWfAH+I6M7MaNP2GMFFys6OUJhwK6/UXdbNiOYEhMEjW5nF/LvBKynb7uHn0FP0e9Z
bLtGaX9UAK5XV7R4mI3yuKnWkNHi5PYjdVR24rzkdRBFwbpBI/vJxw09964z6wrKM+DplB2niX8e
WP87r02qK+5cpX1H9m1OgJG0YScMsppStfgFyoMIFySiKyHXKGAuklWm1jUbUe6SF9DTs05g1CM/
0cm/VBNEl0qvVW1csezDrmroHG0livHZFLEIL9XseEYoqiy7B3ab4Czsy/Buar4rmHOcCqEhQQYE
7kCWmqwHl1lNQBsWSMXnQWadaCWPcWSX4TXc9oCFQ9P6OtwW5iZCpQ7FCeXpwVr6c3/tsagvT/XZ
r1O8GfQftpVg8/nUGkfDooJVVu2IICPq/hXTycJQdE7QmEtSghqIHa/vlbhmptBBl49tahfZZsu1
x81PGuRIhmqjtIsFHfOsggNN+4fTOtAOBvKzMI2kpBAuHzerIoN60dlM9N33aEjFGtFNmO3mkwKg
WEtonrS28owXBDvGlhzhGsMl5s/2EtrJvblDg6/1VLSQUSvT7kf7+JrGM97FMxxuiPSJ6baA8Jv/
6/K0ZVfhRiq69ZwM+xLcojwj3xL9ssYvk39GLN7MVlAPKtgXDbsEZN95uLsGrDaHeQc95XNfFQbs
uLn4D86hcxOKQWoacYhtfoqONZzFy3XYMUEGMYF5UokNI7LQG/Wnn5lKAn1yZB36Aw4rMgdRfot0
RIZWpZenQPeULDMhAMBALMo7p7ihSsmRee7HZ7BFK7Z3LUbCsvuk42KcKBXXoaR5iCIwAqxmUCWj
VgTF0dCRDNXypUf4YD0vp+il6dnrsve9fdRtnlUlwqsiDUbNONbSqafhNysrGxEHOOTLmqeHDCvJ
/DJUiH4FGxpbBale6iV888eeQqZGaynbtWYODE9YOgWs0kgxoltgxT2LJLDVmrHsJdw5cuT1Mnmo
isNU9YOWClZQSG6b9K9skid4mTZ1dHDL6EM3eChBpTT7+OSDYkQYy3KSSmj+9fuASwwl1WoPr2wa
2WKYbQCLuZJNLb/JZx1UdRUiSblvO0OuZMVvEmwsSemxqWLySxJYSiBvz72UvzaDEMP2WxQDBXjl
IKDutzpufCvonU7xL109EjiiYpXLGEMx9/HfzXMrB//LifIpIBmiRkRXfyYkvUsmUleYTetSWCNW
9nGIgjpmWYej0UQs6Du+GL7E05L3RrQZNFIrBy3rfKdCyr43beDwrcyEH97dlugNXOH8GHz4K2CA
IwSlBT6Iwue6EY2MQ4bvVE2N3T7AS+ZzH45Kg4IlvxpMo3lY/m3oxpDRyrKHjWhkyPnCiu7wPbC1
14BwerEp9elGRAHh+FtcG4jnbts8Iu9pKHjs3NuVyTqM3Rz5bg2Ee4F7HBITcwOnaCoveJRVuyHE
5UJJQY1F3yt+OMza0MmNMjzhKJM04xW12uvnzLLQkvKS1cv7n+yHIhKGBle1TXYAN+94/aKqhtRj
8IkV85Us3u45/og+gMLDsTpa8viUbG5zUfyPrTIdSiALZcxZksvDbYWG/EpBN9Kfozop6FrazQ7V
SbZ/ubSstDRu1mhpupolp1Kca6NalErezu0RV5oJS+CH05qD9rp20Dpm0kIu8r4ybgQqtRM3KAyt
iFQb4lRFVHLa+p8qtcVTOcicqpm6UeHqZIr3kZkQwQcAbKrRYzaztWoFImXApIdMR0irz0kcLogn
Sg1DaCX36WHA92QtilmvUe4sKUIXekOolnrJ1bRHT09j6a7dpdgZ+0YDA4v/fI1aq0amNpFkxpG2
NPuGZwUWqPtEJcmAcNnXxjTsSmhNxYOTO2lpiBbyqG9nmaN48z95eoUZUF0KwbEoOe+Z1uBTBqzQ
wnE/S1ldG+0ZzoQvrRnq8C1VBUh2sLjPvxCnQ4i+XAxAFE0A25EAyPWVueB0OOhBgyjqRg3zq07R
V2MZVfTQMPl4VpaS3AeM2/s9dD/rsV5ySwciXwWj5SsUxaz1zIo2cm1Jc12n2i4I6bp8MGv+UKLZ
zZVhNlTNu1ch185u+3P6yxNO1HkyGoNUKuicumgCkZTHAA4GvaW2eDs93GUVI2JQU0Md0tg+Dcy8
Zajq+pTIl3KNzrMrWJBjj5Oy68ZhAIcJ0PD+6tHIsva07rz0m2U06mwxi1dsv96/bofNVnLETrQ3
zCAsg1/FTZSbaac/OQnOfNWRsokCd3mNYPikBwEjRjK4k3mzjvIrm10t4GSl5oxgzrDwzINwm0uS
rYj6f5ZKoaczvb0O9BNL2nFenkx7Ih/do0Zl+HMnd8M2uX919vV+6NFtYswKF5xCIiVkmKEBYKBq
XtUscMVzjpPKO8kxv1NYZq+s+C2ROP5pwhCzxKrD1keaOLq3fvMkstvUZWVB4h83+SngI/VXH4Gv
W4SlplTJJ/Ne//icHvYZ+9eejuymTmd1GB7uQVNcM4iF2flWfluRMNPWnSpq2pLkskIPEDsTuynd
bRw2/8WJlkir++iGaCMFVbsfb0XuVv2XoWozg9sLQnvhG48qPSX4zZKSSMYzBbFZN8W6SJbaz+6X
F+XbREBDROHUrLYPXzdg7OOPaMnjafRdwKhBpl8W+cKLTbkOjTitYS5IXE8C+7i1RkLB4pAUzPxy
kJlpt6LVoTRFich4S/vi7SaqsUk8BzN2w74CXRuifdzWffWbz6g0uR1HGJGBrAoW7RvZ0BvVFSer
27paQQ+pujCNaxY2jbzOU9ohUbQTU4ehHHJpAQoVBjwxRbfXDG7Ono4gjty1KktitggjCTc7TgsP
fq2cL35lv01nBhz4ynEv7lrsnRJrhXF1QaQDgWmMm5EyRWJjQaDE6xfWF0gYqEVZLsPQJ4yJDyE6
b29oehv+9FoyEziKXCzisxUpxtABI67ZCiWmVocUeQMainRQjM+PjZvIQfTPeAouIo+r7CmpVH0+
BA3spKR4xP9NYmHOY43n0y2/kyMoaUofV+NeoOUAwQDV3B654MDY9TYvjvcR1umf7MHqLkN5luuQ
u+4Gg8ifG6fW/zHF5mJf0FDG8iK53ZTM3uzNsL4P1VjVeoNnk3ObuLS3W9nvB1EI0TaYN675xQXH
v38kPfq1whmht3Uwk9XwljaZUEFOcqPMdrX1AYEUXZCZbaq2tW4yxMwJTdFIhWbkIpQJIQlYOdBp
UePXvj9AKiLbVJbZuNacPt9bPmexJCIgmNOfjtiBUb3F/qeFXllHa7GbPjVzkIJIt3oVA9D+deLN
fO0CbioOdGIDxsuAxR/z89PiP36Mqeo3QrKwOBVIcYOFrce6JoW1KsquKH4O/BZtZ5uqklN9p9KT
erdD7H6J/kRyELNt4Bok4335GzgQ8aC3Y67enR762Knel5I7/pPwIrZowKKuN7vvM4XIyAtmnU9u
KkihTvAMXDEn03ArhH3CuhS1Fx11eA94keRU8m5B5g08fmWvohJR7hwjv1etmkhYTEOzd1aG2Jdu
gxiIy+EjpaQPm4DcnGQtg0Dfuh+DFeUceghIRqsb+SsD3oU9A1bfWjYk/ERUN7FKS7UT3sCF0Bpl
OaH7/zjrIe/z5zzDFU0ldcvO64kCS//EKuPXgDYHquPTl4LHJ/BleWyIbQVOE8bKs4W1a2IUK3Vi
GmIXgvbP8iTOOK53XnyTmpw5PBi6Ov0nnw/c7Lmv3cx9bojVVQApUGkOOoOhcbUTWSX+bURlpFur
xQ73Uq2aOCzuiaSA8lm6mCxoEcV4WtvsRP+dyD9JYc2Qut3V415V/xnslVZFVFQpuKa3DRanvamx
f+SDUk8Xr15uTouVs4jIrv5bfk9dBtAA3blmyHUL4YsIapFeGoJ71CvkYC1zrR3JTKyaY8FwV8Mt
3UZUc+21MNb2P0QY6DdIR96RVAqg6BpwAJkB+28pYGqcd2vNMEF+s2EKOI/J7yoIyM+zbvcO0Gax
yoAXK6HZJDXqTvWQbXGL9gKGzzYh4A9ft69805hxFoRcIfVvZZBaceZr5AnE4PEmp57JO17v8Ypk
AXesMKB0hN1bAmMul2/8pV61rr2+E0V+eIF4QEX7jp93MC7JKiZpoZ6PNupyqWBV7dzxvPm6ctso
zuLc+hzsfxyxP4GJ1aSVGob20BZKqurXskrbD2axtk1M/X1Ep+NB1/hmD5KCVoPzoij636tsY42I
vZ+nW3cHdUKKZhvQlXuI5Xl0i/mVHoSHV/UqhVs/Yn0c5I9S12U7q9eiqaX8saHNL0/8WBQxTaqj
saLDxBlXOMwTK7p9evqVmV2veiqe23+W2JoXe+yJ9sNIic7i+kX+xQYmPhkBw/vqqbQ1gtmyN2QK
CWwF0cRsbggxgfzKGZQ3T/8WVI4BIYipVxb16B7h4mTP++Ex0cXUk3/QLd1iy95BHeKKteuWv/hZ
mIX40+e1iIGbX1+cloVefIR9CNFAHqzjb95oDtlJS3DlVZI+4OYbDXZkHIBRVShnEnROOVmblCHN
dju+xyJFyLy8+WztYq9IEY3sUyQ/f66UVbIQ3YwsZxN27xg9s7Fw2re8J0ysxznN42jaSsapKOpm
7BA5KoU74CM4O8s7sCLiw7tEKzv+RF8kTkuvdvf9aXCCyZokNrJ+pCr/Owtv9ibGjxmNyh0+zfWU
siPYvSTckWx5u+kFrW43k9WICe3KK2aZrFwi/z85wWrSPLJh0PHLYYNmMB4Gs96+n3DfzGeNFeG+
OgaZ1bfI8qedREoLoCLeGzKhEw1MPSl9EgK/ofUNHCQ5YXhhKqvebELZeDLBqRAjEyLR6nPHqj2q
6K8o2tDWiZM2Nv+zH9LI0mMYCCRA7v8iTOafcHVXvmYM/cY/oLYRnzeYWqkCe6MKvudEFd8JC6C7
F5LwmzcCI1Kz7v7JhG+9sp1IY/NKhkVCea4fFamcpR5vDtjGKsUYEAGPy45kg/nIedyd5YjfTMtX
ivCOUGioWyevCVOITBLPKmcbRDWQSQWOKGfOvewuJIwcsmrAqtk6y7hiEMS47/0wCyCzioI+wbmL
5GGYtmt0PA7gdDta3w3hUMhhi3SdUd5SvDvCo31UyR961RfNALuwJ2XQGMNdwuuJqjsBIYKId03l
UwKBscgBXQrIrcPVKVPjTwcSPUzscyoUFKcKLuX4a6WSLE6vn+t392yGO3eSroEg7O0gGXI6dzVj
6K4c9zYqZUvjz6u7pcPQU0Cg8dSXbjfbS1TJP4ZpAXP0RH5QQset7fHZs9CBmHCfmHIZS64R+Uhd
qOcaIU5vxS5U5SBsjifygN1z6H5Gh5V9qTVt4HS2fNrLbyY6svBOLbvK0N5aFttkrslPUOBKvdpr
FIjr0bG/5J5Vnnm7xz0t0/+RMSdT8oxIU37ZSWhv0ka6KbUoQ+rkAV1cjZN9SagISlvHobjWbtHi
sLCX/dwjues4wkJ6vmnL+4Wzm1PbO+zNNZ6XgqZy0tmWP3x2nV9+OCuQJZNakXFkWE/Wu6kwAbSC
0aonEhzA7wbEbPWlz7oCryIsnoBnAmE5eZbaUCLeaG6hNXUtyE6hHH+YCmjvnOT0ZGCUBCYYKoRI
Bc+kh0/iKZvIrGKMC8em8NV1uHyf1+r5WPmqWVIwYIQmcYFowDODhvKsJRgmZh06qDNK2yz3Ed3q
/OcVWVnKIRInQTaWDD9iImd4tFpFpXXYBhZqajnsRxbM2XcaBUSwpId5tYXse05HPuYEdss1Cuz1
h+hcdQfB2je1pPQT8V8eaSLYnu6ihjU32vFIB9pO07ulg8s1V11FYu4pPgvZsnwq/Jc2+VSgYqm1
G+Vo9AVrI6pQm0rqwfCgdfnPMJOHmWtcmGxfU+YC2Hizyjh+2cZdV3JrSPzVEbHuhskouTdBGC3U
Vu+eSjGRYh4hW4w4Y1K2qquON3Yj3KD3yN4TiQf27X7QqmVhwIgdB/Mmm8kfypg6RbuJ5B0RIOCp
Egt2MkzDJel/2lEFSCq/b02JIZSz5fhrpzINKc4PpxLMEisAK/EUeA4kvHg6Zq9c5WmtntDgFj/x
eSdGzieSzfmk/hvmldM1LYfw1jddYP33NP9GLVVmbbn2vhi+fSHnUw1e9NcNgRvc6N8jbVVVtLZT
KMjdCy+wHexxXDJDPn46IlYWknxNuOLHgtikHEDjtTic5J8VxgZG7hYX5uGGbIfQrByARMsJ+xbp
JcuuJbShlvyUvpMbIAjwn3bQPdmhyL3v4O75Vy6FVRAZC60QNIVu538nu+U857pvTgaGZj65mZxN
+Lt9Mc12/ncOEpg6n7SK+NieiY3R++by6N4sZm2g2vauzOagHONhekaJlEh76p1eR/BqmVnM6KMl
vbtRzngThH1cAkfnQ0YmawaIflUo2bbK90a8PEzmU3Ngirkl1sAUgmNk1Oyiw8THVj4UBaEZm/K0
SpPlWjN7C/f2K2vuxBosqWFoT35B4whnciIhtRYSuKV2nxSYLAbTMvcxd/c9QgZ2weHcNRNH2p8P
dgDKDwh2RNGE0q/M9h3sXaBxUytj8KZOTrHf5JzT8Qwa8n1tsGmd/txjpLoYdMftMiELIBDlV5c4
kJv6oQYer40lYkxUWijL7knlg2XAJEkxtiQqtAPo+HWTceeGbLO4yxTLMxgYFr1to3fsMSoSDbX2
VlUvtEVFqHZHxWaRgHhMoevQfsx1hbtafy+tfvVgIJl4yQl2cL4E4GLrX3kzMdJUujHTRaEqZJER
r1dMb4O3AdQr2cpL4rRnaXWmlcRGHUG+/CRv5NHA9ZTsAgsUtyMGo8Y0Q/k/+kkp4yBM6fAWyq9T
YonEPrOB0u2Mgqu/epylLw0IOttuVDHFt0EcKo0j26W/A1lAGqsPM6rSaoXz0DzD847e9VmCUm49
TAPbrYshQKPWGEjm3lJ4XKDM+tyfTwitZl2UYryrM09Ccwzal0SaaMKuAIrn+fQJ76Ns/+3vi4lz
99xBMqbY3oNIMCNoooqekAA5tkcPID+LkjBJ8eaUYtbmma+UnLJsfyVr3oG1fFp/COsZqUkkZ4bj
/I1TruWudT0GP0UTHlOoKTT9NoZcK+6zV1f0u4Vsxa5cy9h+dxmRyrRu8mLaECuW6ZQWi5b25F0v
0pAY8qj7pb11X/Hed3naPU4mUjBn3YTkj+nROLPvAkBw21AwhTegj5dgjzVRF+f15jumLO1bnYVo
ueOFBsZaVi5Wix8OTuTdT0b2lQKlC1foHbgd1iriom/XmDdPoNrjIBnkjJDZc14+60E1yV38t+0d
knVhZm/Wae2mUVaeSoyKSCKGfzP2IoTU+IfMzl3XrUe+Lr03Xoc8rCfSlqNn7glPSXYpL1FrE1jS
QXe2ILNPDfyI9ykfiCERpQvhlxn5uKkmCR2JW4I6cUvxB/14qZWsIbpPwmFy076qZZqaHJwamN/h
Xz+QDRnSOQZvG3isyXhL25W1Zsumt7GEN4js2RqJIgTeC2/4eaby96Dp1HHd7utNbu1hsr/TJc4P
ULEB+J6ZnrSl7tqZY/ALMSRn54YLdhtD7+sKW+zbuEaNlg/eLUl85k4Rw6eBLueby0XxS1BKfx8r
OsQ+p+TpvW4N1fWfl9HE8351bN1MapMpbFSZNBZqHFO7csoR+aHvv8Bk8hkTNPzISqYaicAJaYy9
Lq5F2wuDsdlaGwoOeIk5ZmhqOwtOtOH6pEc787bJbut7X2PTbYO6eO31OJk7p7RfrTAu8ctAJHWq
a95pTuk+4OUxmhezxGVCTWNed3fCKTqL5cxCHUdM1OEOYCLniU/N5Fv0aZJA6usPHB4rjgvGKfMo
ZRt9jHgo6NmdmYQqdH4No6rfYbdMXhFIvwtEJvGwS9ajeMjCbTNE7TCLawUn7h8axKjEtL0FHURN
OJTHLQGZnpswprg9xaEts92frUSfjhtbeq0ZS3fZ/XcWOwiKK9YxroSxQYcBuW6yFHsCdgy0VeNJ
3ZqS1cxYwFyMQZkwxT39eN7bc3/5wbu2JsF98BXfAl9yqezjfDQ53V7kSbmu5PB2yhiLvm7SKsU3
i0qvUSddV3mnyjTUSJ0osHX85uJa1wjFdpFJu3L4lAfkqCwRJRkT+jGAbuYDECKMxeJYDdJ0JPAb
juqfsIURBEJKu6h7FQkcnNa5PhPkMBVMPMWoJfIm7UMv99tlSqGKEQgYHFRqMc9N2rM9RK+XYHHE
OtutTyt4VLCY3J/X3LYkZML54sXKbIjCXhpAr0oxDgQQ+6xxCqWVMjobdnK6oQlhjxaHBB0ZWIu7
Kdjw3hBT/mMmhBdceBmBPhXrnyloS3R1upCrGov32aDLNJ4Erp7uRfF1b9rA5i9k+kbBujVOyGeh
ibCPsjtTviRRS77bJ5ZoZzPjgyq1ISuZTXRab5Wzh7MuJKEnHFtIhiuzimli6P+lDNXYZLR0arJT
5bMerw5yQYh6qAC28CtxtRT7IT1VfGkmYuqRWvUSqHtqbIR5d1vHK2YkR+arxFSGBobUKdv/QkWX
L80HRKBzb44GhGUAb7GH14yE5EtQdXZqt+nWK1GFOPLf8f+2M3c0fdJ/nIeSFur79glQvAHp61yT
gs7SNdDR8mcj41PS6T+GXDDwLW/GDasnAvyMqQrPSwP9XTeKDP/M+G0JdE8htPM77Zo4LvHWGZC/
55YeOTqTfBl8XLqMx+km1sztzXXNG8d6bnscU4gJLaSJe+zCP8/L8FdZK6S/Xl2OqW1MZiETS7GU
vRVtP7dcSLGjs3t3gVLVyDMYBBpzJXBLL00QZc4DVMxhECqcpsRNPXBVCMGo15ZYdSmP0p9n+ATX
sHiV7Ax1xz4LzEGHbKiolNlK2AliO71mvbR2V7IbAH3Icy4tgNHrww15LZR71ysbAGc8D3/sa5dx
U/VEpHzvwATbxWIMPQdU6w1E4zxaq38PXKUpVxK/5wlzDeGyanCenYLwCZEcU1ziHVshHpQv1UYv
qAqy+BKpj56tkpDsyCtuqH+R9t78QS5IOgi0wIhv0Su4kj8cjJ1eo+Z3qOWn2B+kFRzSz35+NCQE
SBJPKKjqHHTJFOSKo9t/vNE0UZwqTQmNqGOFNPYl0pY5DQJZFVPBz7uXpaqInVuLcB79XYQyinYE
tHZgTCCqsbk0y4hXYn7dsMOoATP0hypAhoFQqjXVdgl24fogRGtaoOf5mkaLbTupYb3ylxq2zdkA
+IJzaA1tS5T0MPAU7Y1ZBNYEFczc3lOWJFvkpsMUUvOYHTcrBJg5nrXYnElqxzW8xqa2/a72Pryv
n4Pgrr/HX5cxha5CrJkz/utSfZVSuFks4UZ1ieUB5I4vcp7POisnpbuu+dQ/jMs6+Dka/t+C6NY2
tVRP+SvZb8QqxJGkt1cxxUAgedzXvDfORnJgG1E5k8xi6w9BnPrdQZwXcfjnaikBb71mZ5+9kHjS
LDOE+dIhvE8vQfGCJhgeaFEUz4sCZNBxIKGF5S6IGO3HQo640nycWhz9T0osiXjyV760U3q1y/b4
49T11f09NwlPXpXkgSozwOKnbT4MNTWorLvX58DY7EFvZEAmXw6OCYImGUdgY85HQK31eNstL3C8
tdOzyI8Iiyfq81Dg9IhyYzWmzuwkn/XvJZC7YD/gtRNKjsyZqLjIMcaHcs8p/uTXI1ZOs1lxO2KV
zJS2jtXozxJWzGMQYGEpiPMarrV13dKdBUNSSqtBGvlQF/QFPxW2y9FIH11TXhyl2zelnNNFo8Be
7gl9Z+3fijdwr3OqMIXuNEyxVJIG6mp0I9YcwpNTlfE+UKCVxcM2A/4Wn1HTfV6BsrcL3RiwCvRp
EswvAMPbR+4jJdlUYJvlXrqUkRXBCaPmEGBNTf5qKP+lh/jSBdW/liamxU9LwAi8n3+woh4jiZoE
RJ1FO+dB8zWhd8oqrYIW/BOBzgudk8FJfMRWOcn7Ps7OgH31GqyHqtQ52eodY9WGTt8WM0pqB0aV
5slmsi8lYbD8SRFthElP+ZthpZDwU3Mmx8ZJv9qjU7rZAsL+rDPVgbsmHNYiGAtGHB4bNrMI5kvd
veuHQVEnV9b3fhsdwNHQF9QvpQfQN7pKi3d+N9ccY4RO2AAM7mgXOtxl9j/u3xflQfb5n3PgCTV4
76ZcGn7pDq9BnC2nH9YkzibmnteCs5w/m76d5Nc59ddtU4mzRYZkF13ivlASDrOeOs5DtJp9sfCS
T2+nkoVm3WoaxgZHGLNCLWOKbPlMxSOSEBsjAqacEXZ4KExT9Wu3g1fAt8ew60TKfsymZ2CI+0pP
2xUpCiZEHtWL6WiQXpNgO4Rp8vfnx1Oy7y1Z2zo9f3tsvPU6IGw1KaFUC5G/+uvE8Cu69QxiVilW
bZ7i1Gkq0EIcprYrHMQ5CcZwcn/7vRYDosDs6kpJ6vnS7u0KQKZnfLdJ67IvdT7rhjAk43sHpKfp
s1JdPdL+NyincSAJ6H5klNa8feTRzCJvcJkn2FAaNmKSWykMDpxeXlexxjIuIlJZslX3XH0jYYx1
4kn63ATltk5/CJxo1+lBKYMpl/+N6gC2U6uBgJyy0HqLE8GUiEKPTi6a1roRqLHGqU2ScFMHAC/E
llcTlELvJRR9/fc/zk1wGxSBFSmsN82IZr3xjkDL19a1hrN7xLrVXNW8YVPYQupQRolfOFmcM2sB
vYo/8a8bWdCLbFWOhgzfNFsI4E/3A6xPipVJfur57dqpCxVzVuJOSeVF2A/zXzb97Wq/2uzs0xZZ
hOYvheD6G+fNc2Xkdi7bUhEhjx1O52ruvcsCWitgMLuWcK0a7qex3Q2g1dBCTlcVwuA8kMICABD2
7tivnO+vfzngnbiQEI2j3ieiRZndWRpwhvluhizr564JcDXRXsPG6Z4949gbkZBl7QymSYRvqRI/
ANIvnGEHqUi+Rea+FUXYbFffAj27CaCSl72vtPU3tFeJmIvqvQTRzqGiX9x9GJzfdDbZh6xPdYNR
rhEcOxV3NXCEAruDFPQcAeyOugCCZcURoj+F0mDwW1unt76VW0TfrgzwOX+kWz78GZedGQUeslnG
6lDs+GvUUqUyY/j13zuLde7fJnYhGliC0LrNgxfxnJF6MIgMLYknOmkyG5phID0SWcmuiEahn4yg
G1xE0pKotSpGhUld3XWMkA32GJFdm5kEuuwQoEWgVQSWaAYU2pxxc9SJAp5TNsDt1DRC1jm5yhpF
d9/VQDmT6JiNdJx3j8WPz40R2zVBJBngES79F122wn3KgRtuHMwnGixiALsXu5/4wJgPobYNeaeq
rbq02B3QpVyscVPRMNThVGgEc+7s+kBhaVYgZJJIa1BwZ3oU90OzWHvrxNNRy8H26wmHxnrozRef
B66XSbPsU7CzSAC5g++mjZ+KHTnKyW2xSBvMvx9R+3Io9j8pYUTnCp2TwB9enrw7O8EABlQymkpG
LcPNDkARE1tBiKKbX2Febhw8gaNC+FZG7tYB8FlsDKoWUEd1xsi70+LqYkVl8wb89ImpQnM4hKEf
DAT8PG61aoz4jrm2kfUE55HVqtWLANAlHM68n3piPaJ7ZFFetVEJmdFgd3/1cznv+1CnGPQPlE+K
clCzyr7Ne5CkmuN6nerdGqeIvVCRyYqdwQuRSSg3R7DvFHiNp8go0DgpwD6meirLRq5/SLfVv/J/
S5sMDnhluxWottn5N/5/276Bv97iVstg1KBzNdnu+/2ESigX/7m1oLf3iBfMHDnaYcQgV7QWw/1m
gccf0q/CqiY3/PAFjKOyDNFseLO52a3yeJBdSyycDfuVwt2qPfj/Ie5KqSCG/Ugeb+mVwu22weGf
/GjvEbMLb//9HGxqp28mnIehy217+Szd/DorQW0KXJO2PptmX2LYN+0tLv5dr4+//Mml7ujHjZMy
WRzjBncgXlwiICnJG2ih32YwGBCfsYhi6h/ZwjLfKJROfaS3aaTWCVV55Pk1qWd63AqWWJAv+drg
PrtYhPEu6tBj3UefmbcPetLRVvaJMWNFJB+6A5prE3cakwIoq4Bw7ewuk8cCpN+fst+UypxmuXG9
WHPeIn5A/YjhHIKue5OxQu6eQ++zPZ4p4iTG1qW8fMAczpdWp3N9ftw7/Y9J3St9IUDhFviPT7Ak
u8Wax9fflvPXLPASvlR3O3wN7VgdUZKYayzofywKCjJYb0S+nZRlaOmyWgeMRI/MgIg4FVW0rHfl
DQfTS1n1qs4ugG6wKM0SuxVd0rV7Pera/J+b0VqMQhNSHBMZCm+mDNzw0wdL3JAfVDx+wXxnRF0A
OUPdTAKzl6JMH/D85PVYpYwVeA9DY6NEk4BneoN9dy2U8K4VPUXGSvsZvwfCrUlJEoRZUhkyv4GN
vfnI7nywxQPU+TJ+RHtd7VR5BJqcOHmMXJfxTqVOfyuOjoWc2lgVb3ybUYLsEgzXLrA4qjqzm1cD
ywL9hd+LJrA3Mdy4mLO+HRAFwbmGzha9C0huQ/w2jwCa0vpFO+mne4BHuX7A+Q0FK+kuD1TVkyP6
ZaUUzBqKqBo6XrAxO0tp2T85G02KZ1td6FvDAUlZEm+y6IyEmWQrgueWoB/fJS/P4GNbW0tFfrGB
VYy5zzkY5flVaT8QAEStDXHvcikOZg5kf9QysJzySkgAklRsS2/ppX9dGjq67hhcRWp+Wy/SYkWZ
DA1sesoo4/y8Z+TmlZDVSEmf5eb5msXU0IjnEcBVm6ZOzKzQPxgJXEEp3u4sGwT5HRO9eVX9G0mz
vG5XejxGBZtgKxJHkWRr4ra8u55g/kPV1WMKuDbDBQw7/c+UYBFWrZtiLItZyJ/4MaSzRfrtNfoq
q90m6ClEsNqMNj1+eWGvFyDoXLX0i9UveKjq596NRqNiKdbihFYiZMhwHqwfsGbo+cXo9A3OzxVD
emhCiy0p813wr+9MjPz3cMzH6Al7fs1NjRL91I7c/geuTHJyQVDbihD+xYfnKZ9obE4yBwat4RSL
Sjm4Yazuavq+Fywx0GzVHOFmHLB2n/jABQ67yxRI7xRB20KKaSD0iiTWG29Qo7BaWwW4mJ5bqtE6
mzVQGtt55l+yHRPbouQxi880rou8N/cDgOFCzJ8hGYu4+yNE5TZD+lcgtHMgNuJkkaD9vQv+jwut
6jqo7uj+lXKze/+60WyPNxsZuHx8hapdK6bGRslWjns28tSdvlA2BNAt4Txn7QBBPztvRJNxskh2
9Fy+RvPrgT8hCkV+cNixvkiB5cJMKZHBmHHgOpGkzEl8Ok40Twuq3ESV9ITznUbQptDO7mQNsxi2
IpcNBCov4u+qjQacwKye+AXExewocvvnUv6KTkxHCux73kaSCZReQSXfjwRuQfG4LxREGx+sAoUd
NpfzywLLFN2ybL4KYSKdxBgL2gg1dOx3G1hAWsYrojtW4vt0b0YqTP5pUNItj5nbvdEn1SeSGyh+
TugZnoHvyrsUGWX4Xw+Dhy1REGfY7gFxh/jXsoOLvlkDOnqDPRc0VV7oTycOEDiVsZ6UruI/r+at
q01XZtlk9sSB0sVHmjMWbpf0TZq8YfLNYjLUkn1NLWLJMzR+6KUw46a2AUCMrcu3BWZ2Xp9Rhz7Q
TOWE1Jfl/MgmOERSzOiNdwzaHCDpoG0TBAjtCsg7nWmHespLmGblXDWvKfAiEivO+/vAdK7Xd6z9
mB+db2pq40J+b1ok0vUzSiTE9jM2frMJ7gM7MqfGCL+wo5EZo9nMGq/hTrrsz2mWVtjvL0pVBm8w
659xfGfGjv/NLv3UiusK1HkqBNrenpExTF5lCSBQy385g/y9XuwjXsfiCCjt18QfChuB91IxVNQu
xddwSNuHyegb5/rnsFiJS87FyrkkG1oFOpGJ8Z9GwrCR29UPAA5Li+LC30gkVx4SYcVa8k1hrO58
bCIDnJFVtLZu6bT0Rscad5gooeqR+aaVakLf+K8SsVka9Lv9AD41gIDeP1yzrdjBbQxyYgv0i7Es
p2VexfynrCQK3D6hnBKyJpnhTpoiORZGd7kEx/BEPEsemJOqwR2iQOQVddUp8qMz+4MH5oOSVN6j
KqYwXhZs1vI2SUQSX4ta9K05Qs8bHRFy2KsZhJa8mFHZoq+sWc07JBm9cbg7WJ3/6uvE7QA55qPC
sABAjJycT7qjNfqrKhRi6kmY5CN5jyFXF3lH4Lp28FIieTHX+IKLFfGHn58143uQN3TMl4ebVMXE
ygRe6VUDjt04D9Crn6ozWxtOT/OSj697Ax2s3Ah2QTrF9fW46g4zA0lJBdr/qyKK0kHRFbD3CwO4
XVwdk3NnZRdPx48pwT8cMl1cwI+xl4IcvcOf2XkQaFK7smdmxq/IQFjYZBMBA1tNtlaqQYAEUIgs
82ZkFVdBrWpbnr8xQdgPgaSFKWEcGzC1Cge/YcWWxqlmRQxxkN+4C0gsP/VN7I/cMbwduNRtuhKk
RfDM1AGhv1NV/ux/h7EpUt99DNQZo+cGWVx1x//FG8ImgkKwat4tgReYLbYv7NjkiJ0Un/OZc/kM
tWHDyrUFYlFFbaSB6WheMxm/nAocOtUJ/UmvKVoNos2egiT0bKzAcOI9VL7473qRG26ngJG10PyO
/JCr+FxjQySlhusM2DywKna1GM+Fin0cwBF36APf6VNyyYfswzJ3BaI9d5//mnh++twwcq/60oYd
ZsvCa6JJO0WJe6dQEhQBhpOJ6XfimVGuMq63ejrz02VqB4hFUz4X369X1fR89doyULvoFw0xqcqd
tH6f4Qb3YcYWJNV2BK46zSqoc9N8qfW++VQUIlchtufqUCHhtyhk8+X9f37CtpzX2DBFCtDvdvLL
c4XgiGz2m+3smkOeLHCnw6ROkeQM+2RCxOuy/SzDOg6LGIr4HDIadvAakxpHGTKDNAM3eRlQZHrA
KiVwh62qaMns5VwDqKuPoQotC6CuF0uAlbRUobIMW79MkIrCWYnYOgQj0SgD1SEfn07IeZ538tk9
opVlXMxBdmb7UqHeC+tFvbHzTab5EYOzBigSS5o1Tst2x/UfebL2fPfssz8cbUHlYULPin6JzDe5
smBgV0Mkz5vlzHfbWnjc9zcvkBTEB4W6z/nJ5gqZiiMFBf+ic63o6d1QmgYlnPWRdrb8UCRWxn9y
DvetIGP1wWQsCDJ6BcxMliFIzXkJX2uVqrMe1/FSCKtlBdt/c8GdBqV3UGsCYERvBMoN78PO46AK
P9m1HUBcxjXTMhDwCNHtCzZL4pX4E7R7qN2JBKaN0C2yZB9IdXxv1SAtO2I0pV+L2fc7WLvDPuoi
jRCuGO2sroN9tBd/0tgyA4wF/FcmH0/mvo7P2QO+3Yj293yc6OZmw84RjGdD7DnjEkUV7BzaoyIQ
tjXYHkheP6TNcYAlIFOpw+Y3BIEbK1C6AN2iEkG3g1YyeIeKA6a3RFF/MkyaxsYe9UzvQUWbSeon
brsPKkbQoHzTFULJKshJtrE/Pk9JDfrJxQZR3y0wKR5Irea/qlJUOiCQB0n+6ljdgMWcmPhQvCD4
cISM++SjxNyr5jCMWuuW7a+CWuE0/Qz6R/VRhCDq7UUvL9Quj3mydAnY2vzzIWncbc3e23eKwNDC
dL5/V99LFXlss4Ajr0pN/BBgrgfk+9XBMJbfgBxOYgvhx2RLje2zZMoXrcSf/hWTEmL/5EYJCyfL
VfwPZJUkeFQzAiv3PEs2oAcw95vu5wbP8XifeuiJyxERk+1GyBI/OBe/4ShQmQpj+cJ+Ov5fRzgT
ifT5+fUABdojf1NczJLzZGXCiewHkcp+9YYSLHDciIW5+o6AAoo6LTOvGsNc5gjWMRLhYGXA/QnC
B97zfPBm3pkWcOR1lImspN12coGkgQy54f6AbvNXS7HfCXY9fGRq8sfZBo3Ask3Bd+9xM6v7CDlN
dzt3WFx8MnmJ93bQYslpRgKbcS7ArdERQG213Mg5hPJQcp5kjN2Q5qEKJZqj129SAKW+fcmmZptl
f6pPEMP8kcpUB7pL3U0T2K3TuG/vIJRFzUayNgNHcnL37wx3U1bCBzDsf8mR66K5j3ezlUcn+7oK
7cYP4otMf8lHmPGvxGdqVkBGK04ID3ENBHCEgcC8jzpuwIlwi5kixfovWAvclxhS+5h+zsMD5IFs
O0hEuToo6r0yIisRzp+98gUzVRPakZxzuGSvjgyXr2mZZEgT8/gGS3SmX9XpBiV7SlOo1z3CvRKo
E79W4ipgiFTOV7VcebHCF6DmYQMaDgKmxUgPToikZxQFUObY3G219TjUjt68JlxAnz0akjsr/vxq
WHLObXN/4Y2XwuWIGheuCx6RBlKJx5XW9EFwizzvWJNteUdNReWWJUBudCNx8+AVtMJ4nwnb4eaC
8JeZq1sqWpTs0mWWCbtTi91dwCaCySddTli717DKoK7FPoNf+LO3o1mNTG01D5m819LTrQXw6cvu
nGmpzjyKCWCjIPRoqXCYN4/EfJXnrMWtUuBdqA5r7Yh4pkOKDYk0kHwVWspokyFss72gJLPCJBZW
2W1cwDBbcu5hDYuOF/J8F7PCx/PZDMYJ4HdKunCtz9WK5Z/LzqGsn01csn8MWzrAAID2SwCQ7JGy
WKUYzv5yT3zuEm+ukkfNrgfW2e6IyYcXBYy7lMh9yXf5uWb0xRZqFn0rbJxcnpnqXkvlUTV2XI3K
h1UQ55pdQC9MP2EbdXWdgsTX3L71ebg2hFMwKzxXPudle5BZoW6hg/rjSP6jEotRVqT35CpSrgOc
dJF7c6WC20nh6cIKEdf/3HIE7DjOoxIrlSK++6kuwo8AOtiozFBKJIoarVc2vqMLKkKf5iXi0RMi
PMw6rVJQ9Rk5CaSnHuDBEHW+HDz2gRv3pGmhoCt/QedL8PedqfH5SwFjFk6cXNrkxQ7xYFcG1EzW
LbDvVI2BXKZKPXhul8NUPOF2M5nv93Ygudhx6p+9qFvG5KujAunjIz/p8NAUU7vje6/1YKdiDXE7
IrDdCDmOoX6yOVYUcuPUzFY+8k8EvhSCbjlvU3t8b+LWNPGtSFJs8RUxg84WCPzqQoXj3UhjBaNu
IIExjtaFDi4sHLxaIvqGvqOE4fs7HOyZLHMgtYupfjCkvgcLROeFFhtgkU/d1WBB2lcLgQKo+ssa
225tVmA+in8LQywuhsK7220w4cJCVpkKDq6KvI6Vvd5OTfM26VhffRdnNcCffu5FJhvMDucwvizL
Q83ISkeFitFIjVFZwpKeExI1FP8uSrTX2/JjEOWOA9yhrNgmaoJEM6m0yeXm/+8mrTLvs0+c897U
NOaVyWukp3aXq1AIpOK+gXxCIloe/1nt6aZz7gwvLXF0wxYwdQvCNFpce0ZM5eidh5lDhbSn/hGE
39Mh9FxnEesonEtnClMwHm10oUNxztp95dSgE3qFJW1p2PCvbI8VIcI+EQgMeG3bmg9Hk6eZl6At
EdxmSk8PltggBGJ9LwQGIg8XhOmPhT93XWTNR2cbjE0+m/15Lq58s9slJ3EZ6s60U2h9C53xvr9q
BRC96bW4alhMMrx/NEkF+Lk8XqAFfkJ/aiNd6T4ZDBsSbnrUWEnAsWfzEngmgK6JvuH3DfeJKZ27
+SU9/Kd/odGOwJ0pNOd0lgTNZTTRUy2VqpwX2ZgRS6mT9ayRTDvdpOQha3tflp8djMgEthP32fum
Z5Y6rjc/duN2v53aAllXvjftJLMfDDWsMrVbvNkTOnwFYVcm4mIyXcE3fArX+9y6JNfbrZ/n3qk5
c9uGPIwswwXigRWkeK2Z0GsSFEgrQqUj8QAvcazaXxTmgwcI0kjFSbu4L7U5M9y0n9AIYVomoGMT
LLBQUkUO5VH8oAh8BkZ0oo7PS6BSd42wRVYNrZgCySevmXDKB9LbXYx5HCJHMT0liBrqx72EFbZO
7IWGyQDiYv7Tc+enQgYb+2IGzs52YrJOAZnhvbSVYJooRDoHlT3xqkolhGEHXUn/510obsEz9ukt
owCcDvyqytm7iwLpcIWrspHENQu+vY6UpPzcAm63YmYp/UCmSoYD1YsHk6DKiSvKYHVKGkszyjXA
+OvGUplCcHTqB7bltjDuZmN6Plf/ucmklNUnWtgKTzmZsFENOdk2US9e0Mu8Jq27S0mY1VZNQ0D8
DNWCsYgRDCtMhmDQslUfkt2KMSdYTyXotJ9zwhNA0nPED5BD4FxJNn1ZDVBPKWWRS6ytVHQgDnlB
8/HsqZxgdqsgYoaabuhB8733mtkSsyZtZYWJF0n/JxXR2ur5CGFxxUGCsB/jObTm92O3prMdIQ79
bLKSFnFT2npwhuvnhAJQqJArCoc0cgWBdy8GvcQNDgFcjiswK9kjKbgJhDQ/1cDVQ/P32jJ4vq0e
CbXRi7hAwshVnwJxIys4Ha8LIi0KnqSgcqwlHWNu2KFMxqp7GX8G3MjxORQun8auTYOb0B5qvvBv
SHMO18AZRcGslESrS2EsFtYt3mtt02qXqTIdqNs6M67wDyo8qu7FiNrIMMO7BXigg2u7ds2HDKk2
YmOPCp+5R+tYVcyIv8T6CsgmAyorEj47lDDJ4u4E/3xsdPieGgsnEC+54uD9jz/y7k1kJiefttO8
0f/t9DkM95RUMjJZWjszVg0wn+5O4kFuR24gzrro0vkvqOStlKonY5MLVuF//9BCodTf7Xj3EORp
cFUo5v5bpvWQ1HUenyW/bjIcbQGaaaejHnI5V0D+XMSuf5hgMkIcTkhSapKulAOMlbyRxono8ZFT
EblIZc/AUz548IvnarOvNMn9IbW5ib2pcd+uaQPwsmltUFwmjJvK0oJvJGdLIQAjJfnE34csKvoM
NwmT3ohBzDFYHh9jhQLcE3UE2fRbyE4G89lIKO5wNaJ+9cRIMx57UQ37BuzSbRKDKycoEr9afiPO
3GbmpamAad300X7CTtzOh+Ec6Mf0VBOLn8oS7r0Mc+fEMs/FUs0f+WDI7NEzrelOCfb69zkzwELh
A3Z5LkCGWWpBEnRFNg9mjKN2HfG+C/y1VYNI5jiYfAMRTYp0RqJHpZdt+3oj5TKkgp5eVXO0kpat
X4FvkynJUBKcFBs6QWfvmA1EraJ1x9Nzc2f0fjJqUTl9m92bq6dG2GOXGQsl8+CrG4FS6j+r8wVX
qI3ADvusvrb41qkSedKkNqGKT8mD7p4yEcfG3sdxk77YK42TTg/DKHcy5/tDKin5rczKEcHCKhUI
US2di7B6zQPd6LqxJ8Xen4KmT1fUbIslc4G6h3onjccXxOi25rWP/7vllvNIbIyv7RPuHe7XFie8
U95qNDmqOYxqHjEmiyPlcFNP6DrDx60G3uTgJKZU7CuNcWHBKaWUReeFmYpQAPuSy585UqFVjvT2
h2+yFEhidkXlbMk2gzjLh5qHbqG1kpbZnRY51bnUqEHSYG3cOXdoTyinS/u0NbfXGWsPW6Xzltif
k/tjda0tR63RgBkFmRI34T/IQMIXFhOFf58o3RYWdmMEPwuqjOTP0rBBN7RoofLJz4GDPuw6ChAr
RXaG3BPBCHKcoSYKPXbYkMK7m20I+GzYVv29ioVhPDlXyJrWKp6AaTNRJp573tydmhJh31hjVX8j
92Foww/QPEvo+1s5CPLo6AUk9ZD4FlKI/lSpjlt15MYeLQqvVmn5f7LbQeWIH02uJOJLyfpHPq1u
OFcith0/SjfkmYROHHd9vgur0MpJ4MC0x28rS26T2+juynOVbdyrOXJWE4Ef/yd/matcIm7Jpkx0
BismX1/cQBNmexlCgiSQj0lAZOPfQxDPbLPP4FoUKtwTzQOV01dxfm7E5d7nfQlMGushwbhs1s/i
zR5kAhcCWTikezR74RxAowoyJl+cfujTS2hp9MnaZU9syd9EyZPDZpncWW1/KwGLxNHU2eVUT3zx
VQA+bgGbLI/mqB2w6AmaNth1xgLv/4meMOLNfGOI573bn7w0A2GTs05tnbu7KjXoj+sIl96qcUaw
DnKFV7AR8jlLequ7nYGtFljXWYWORLb2r2yFP2FLM8OaR/eYGh/v9rdiMGhGNEciNDnkxn1AHHfI
ABWIVS0ozEnzBp9JLWZAI0zsJ3c7pBGKFzSNcuvXcCK2q+5cNPIr1L39fKqW5pLk04zbOkC6Q4D9
zT7jVf7MLQ16ycDCcsjVOVtaTcv0GqluOpkPnOwfr/zieSfRj8EBdbqDhQu9v8thJb0IHzSbuzvM
+ecFC4RUlLL9xq8vGz9kAkCQtR73FpJnt6+63K2E03yrT4TMSfcwBCAb52VUED/r7hbKNpyRxIvh
7VCGru7oVHDJFeGFlz08jszqL3gtF68YhEqDQke7izqlVrXK3tZQOm0FNj1/gw9zNLAZWyYo6WXc
H5XPplilM5k31J+OcDSl0f88c0K2BEo7mtN93a54ebgxmNlCpRPVA5LBXjheYvCBRblygdQdVkaA
MvYKYjSSlHXGGS1VfxMJIeaRX3gywwLmCO3u7YZxD0bp4ah8mt33iej5hbtE8fBnQKBXRKtIQhBl
ArrzixfE+dCyKwWIWiilVo/si9WLyOTN/xIHGYX/F6pRnunNgtrhepQUNSr75Qp47fUy8WZbn48P
JLGwt0UY7Ohg0Hjjx6/RHEZ5b2Z8zmRmBJFNGgYQAszhW/zaXG7FiKQay0NsaWgQzwDji/FgkbVu
RoQxY7WBhKi3ITlxsBT52P6NTWlobb264eKkCEKwOX2TO+kaUyQr/UEhpjWoTX/27OcZ5HXTq3LJ
yZYkgu7R3sjMOLW+DkqyYtAXkKR2C1aJeuXv2nDfao6Tywt4BOFn48hofVmBmvpN8QzFFnP58Swl
dNBRsyOeBUXazgcVGYMu0IUjTislf2FrdiKPy0CSVP6JUOVNVdS9xp296VXk5yrrSql86VkW2kK2
q2d/xInGTiprfw/DWk+MUprDgo2iJv/R4JLmTEBWZJNW6eAqqqhcEdb8caW7q5p2aLZ4nCce1Y9t
rO4wh9RROMp/mvEkPO5GOxLkVl/VuNxR64llqwcU6Yb6iZkMAO7aTMDigyNDBsWKotYQljszkLoU
jCF/ewRFwOi1opgyOdqp9z2KhvqwY1RAKVGGK48cSb0YDt4AZNwBE+2HIGT8rK06ePe0qZoo8LLf
ptZjuEbCPZpMbOgdYIBEoPR345HWr1hRXJzT9VUAfHdAN8HAsmqQlNkuXLFx2uxG1HKMqXxo1obJ
8P5ybqHLW0lGxWFgtzh1dnr0YtWui6rmohjis7iBz+Y9JBGrpKDEKROhHA1Jc/pQTHz3pOju96ah
omaNlFHkuBq6FebgrbfLWhWgMkuATJi5Q09S+scMlVNxNf3KJJb90CpOhgmEgflRjUSFcfIacW9a
d2lUIxKGcjyjG7CwtPYDpcYlLZ+Fvl2CK9YE+ozTGmcoYRPL/iZaf5O2TIQ5wA3KkYZ83r9CnKoA
3Y1BwkCCJ+8gsYtpLHQwo3itLN89DY6P56gxWaAlV+vP6euh3/4ZhAbFo1bb101SyKVph75jDLbH
JeQ4+qm7ABSJZja3ZNcHIP1cikNZ5mgHUJhE4XNwuHQvDoQh/pTia38WGAXd/wAFl6C8cQShkWMk
hVRaxQ7O/3VMflXLYsoRsufM4TUpmABUHkHeHHDfUSo0N620DhfUS1qlBwRalj38WnkfELT0Iycj
MBxLtQ2qWwEdyzhxlcWRPpH9rGGs50TW5WaRFk7xMVTzYT9dYEf/AlccFxq5M7OTd/T7tC5fVAn8
iehXtaQkts8FxPqlMOVgCWoWPifEqqkF5UvUiuE5L89G7Cq/DUwVmq1zoi3Fdccr+tsSQ4FghHdK
W6DK2NnQGjLQj/qAnJRxpv9ug5litMrQ4DzR11Smg42+L22rhWKpwKm0mDdQjZcLIr+Gw1xXLMGF
V5fk2zc1bRewBucFPpjC+ySnuZeN/A1xV3WOnZhLyJgS+ro9ciF2GIqUecOxtRYXO0p0yjQ5XBRw
x7vgaH6hXrCjtQ1PVOPJX27o2PgpY5CJog9kd+6dqteYxVxeZy22kQIJbYh21rNOIaVtSxLc1B5j
0oIsteuefAHLL6UXk6jE/5oMQiu+alMDVeA944ofzZnO4qMRMK1vJqF+ZZKJy1ErBfMHUUDq60gw
J44Tq6VjRAHa4tExdyxI/X47W8wQ9ndajmmRM6DxoXU3ondN/uBWJGXbyVfO3dXyaQBfVyDhp4gj
haXllquVKeoStsm5WZhg5w6ZAZDSIEX9H3jnzGc+9CsWhY0dNCqKu7fEE0BgjLGwqMOp+roCsrT8
1u9E+off6rRN/ZK87K5+cPMBGwox90vWQuvGBIEfXGLiLEzjSqX9tQxiihXQVPEwE/MBzkBaGu0z
i8B+w+BtPIxtRco8/UkbRZsrtduTuZdg767ODMSIbrnukCAilC3eXw3EMgt0iliZlVzlYbvWXib3
Edsxoh/rt7iHO8eHL1MZaRnyHPXDVnPN4NTAKLnwqnQY46alYMNdqExly6VKTMpk/f6BENYHXBUi
65abTzbPfZG6sSKJqGxuphslRtMM9YIdc9UM2jmDO2lNB0eUYc7Qc6nL2YE4AVTJGgX0SmYdmCE/
Q36/bgBw6CGJEGH6gzZbr1fgjnmXkt2FEhMxa5mzQcE+MkGRjUczq96XkSaAlLoCRuCSMQ0Zz3PM
NrHoUJxaZ7DnnneHAVO0hWvQsAGGEo5zz0iXFgjCnnhENRDWMpWa4EUeS2TNqYVcAR7LQdgLrG/9
tP2o4En69oHSLHGGvg9rpqHptYaqYvLFsrPWrlQSLDlGSMkSSS6eYZ1Snd2J0qD5oAxRmSMG/hFm
r5vPNQLXQJwNuVRjHS4P6k5njb+Phc+MXT0Bm6UIuP21cnB5DxB+64WbyfSSojfgOwBx3KPbiSd8
PTUM3hwRkNI1espOS4RN3GDpNbewZSrWh9EolP6NGeBL/Kiku8JWjiyllm14sTGnNbfpziD9z5Md
KPmkkeSWIGO5QlgwcPG/3OvS2n3z0tC/IROhyM6R7u080t6xz2LfowHcv9lISWjbmT5fvACKuktB
jOJRfuFIon0jKnyRNynF1A7StrP9P9p+tH6/HBDVOTo2lvlK76UI+OhbMAhKB1w0tMnKY0hsvWMW
cDgJLYWoAjkWpskOA5jblHa0m0P+wr8FNPnnYCP+WiTVrDuDuL5dpdsNS9grRe9D2MLjoDr8zYdd
pscetC3+2REthCy9c9PpB8F2+oa2TcD7wBeWaD8oP6pCTAGE7f3wITMJ7PraTzasDrdI5VX4ii5w
MZJCb8zdvRH8WwkmfaR/eMNnoGlKzjbQRaLA0z8DCvJ4QzYEqKfSs+pmS4TRPQ17uGf+A5StDsL+
Tiwl9cRxg6YIfsSfem3SWHkwm6AaK9XlePf11taN6z2t/XJNXeLPholRKKoFOqBBo91micPJcqya
SPW2/7oG1xwCMb7N6FB09yVQzYqF1pqok2e5A0HLdph2DMK+1YhBurv82+yGsZ+6STzDzSNEt8nQ
IdNiCHpRruBl4jRB0tm7bdGByKgsS5GzjOw+DCKCN7LprUeCBF3dHYW7wIElIhr4NaROiIIq1dmi
TyWPI058F8MScRR+C+fmiViPag1s186rOBAcTtgbNXy0oW0/xquliGW5oAonxPiqOrH5fyt0dbAJ
Z0Wt6JiphgMkQdPx/kyzOpKdFhBjymhh9pWnEwerVW8aCjMe4XUMzcvC2+6JuMaTI2sYe5dY30XB
icvuofWoLGIlFtQWNk+82a1ZpIRJO3ITd+a5G+ONRo8G9QSb8VUMsSmrzrW9jfVPMcDch6vfX922
q4M8VY0wqmZFozV8v87AnklGofaBfNGDw2zvE+u+TLxnsV6mWnycJGe+NnKislwy736pAu4IByhW
K0du4XIaV5l0GYuWg13FHUcEAfl8mvojQYn4An+Xjn3g8ahhTm6xwOjTg++OQ4cHZ5SMYygZv56g
lXRtYhoGimbBAb/34tU7SylNaAPlJvUYDy7h8SaI+ER4/789Ka/uaDSHFbgCDxAylLvzPUgCyGSH
+tYAs7fUvSqJ9cH1+UgmZPJeYB824/bNcp06P08Svw1buMSLQqsFG/OUl2mQffX3FhiWIcXZqVtg
NJCtWIBGeO+qnoskvj88sMEmToYuGVaJo420lhoIgTpiCnAT0EHEtLhNrKZONIOs7Gt7MxDlIZTS
1cDr4HwPnk0pKgGWum7o+ouK2FO15aMt/OzvmA1NWRRB59L2bvS+ohjZhfxd98fFWNygzEXGaoV7
WMj3zIxc+1WhUAYWu7k+5DFWjOg6X/6vr/RTNK20XoOusoM4waxay2npHNpXiD5RfWweWToUBfZS
cCwkVotdIbU+SZ69TtlF3zXAxTh6ZANWJ23s7Pec3zymnK5MHNnYCw0YJ+sUVYX+qfkV0IZJc6A/
VEjdKjE6vkWorECGvAwtwUgE0Qg3kEC1AERp/Ye5/ETNgmDO19XYdRbUN4AyTILwVGJZco6d5Cep
tTwU1tcWLmUVcFPayabgCpYBIVoXWsNvEr+SqeosnS3nYrDj46I/sKdF91veoYCtA3tuXenz9+U2
deybHkq8pCBOK1Lyr9ggTVGmwbW1z1CeLORcXIMQx3s9INq5oA1tn4AcbvgDiXtCNvhvur//E820
ZSJ+KL4Ie0FwK0EjTQPMlJfo3nsI6I8d8xwGvDNTDRQL6W9uBMnR5O739ucihm1KIsKyX5h5zLAm
4gBizk/7SD+mHnLKCOHW8efHTELySw7VzkKMT5pVKJ+Ggsbj4MogAafKRtiqzJVtP1zuoTnv1o8Y
UM0WMC3S2f2MX24AIpixZTngp15HtGKAtO4Yp+1cZM+O6yjjXWBy91Lm1QV4QC8+m9z31a5FXeTH
VipIIEbRUJzFwBD5gf3Cn7HoLOaTIHh4F68xWCUSHJ0nbLqmL9gWnsjsv+6kOgxJvk1CrXEI1BCp
+9sAw9md/kwKzGCBSx3m/BLJRIqW1SiG+skSH1EURRzT1Sbg7S01vBbW5Ei2rSii+wECMdA4hbPL
n1T8uUaxoQ9yYgA9mrT8ZvvoZIp/brOS4xFehWnyI7vr9IgTHd3Roqyh1ytPrXNV8kj6IkwYhRIc
3pZ6UyDgSf3XDFPkCAfxxuWIsPjtcznjTjoxfLS3AHGeLSc6B1eszuxihx+tRbGihYnshGcUUSmA
yxL75FaWPP/SrLgTbAGwf2fLzLGBR71dTnzXx2kMUBoB4iAw0bkK/wx3qNDHQ9Tqh++olcHMeMYN
Jvw22PUuwQ27lkKEsSqrBn0vLNyD0CY/H8L9d/Jj+B/Z8D1Y4EJALj/TAdV79ZqEqlo1W2wgLspO
tkOG4BNEYPCm41a+pgyegEUoY0/HOzG+dAKeQ2bb9haFj0Je6tVLtlokMfb4yz0W/6C3SF1N6NmM
VF8NSJ4LUmSAsjTR+ZzqPFILfU0uJ7/dgJJNifnL+4Uv+3Cvl9VLLsYl7oK8ot/pXNlYyt99YT5u
srTJ/HdtJC07JSzPB7imLtXnUbs3JO1wUgt3ZM3/fJdRS/KqxGc56XcpNhsrBiY8RlRzFRYIBnxo
I9w9vm5r3vrIvIEjGM845vzAbXJsVMsMq9RYl5Rbehcyg+zHI3iEj6eLdJpl7h0cFgasbKmZqL9I
KpqHrsqifmOia9Zr6IC5ld98g+eRa4/h/WUUjOSAap+J1eBPifrY2vBOkaMGJWWwEIs+aWcgi9LS
S9Q5/C7wZgfLfUAl7I8KHN3yyDO9HaaHYUsZhrV5yGwGaAOd132UvHuANJG7M3rlroy/DCGCF0M/
G77EH56rtHWWCArMTxUdT4tEMlwgYDi9VCGt1S+Ceu8D7+QFs1RxZfqgWPQVOfWHBX77mvWkIfaG
oJvsjnA+rlfAGm6pO8gvpVRm9P3UzRTODI76W36lGwvBGxspd11IC7x5opXWyPSltl9UEfFXAcDS
nACaAMni92bWDx3j8E9VvqbTXiFBCbMfV0hPTdzMbWIMBkZ226zKxczScq61xf9SxubzQgvU9ne+
JHbWD9q2T8JchWeOoX+UXCayuqTdYOeh3DFA0hPn7QRLPI1OIhbFxsZcQTVTRPSt0Sg/smwKd7e+
lCAGVKdXwSxwDFoLKK+slsT2oRIksBRgZXi1sTjp2/8kxyJtmm0yby/Zjtfjtzc3kRdW+n6Vtd4p
UrOt5oM4s6R2pnHFfjiAZ2IJZu9MsmxYMgCkmNdQTgoP70rkZFdiS3SZshUOpqXsLpghggKwQkcc
kXHm8UvXGl2J08lmC3EjQhUHnams9Kt18H38F/2En67AzJD1LJnqKh3yCb5DQAbW4gIl6qF+6KOu
SubHjFbzYq816q2gZhaX0qlatOoymqMYVUVVCjCTcG8H548KrjuBc68fIldZhSkpOvuyI//tifwR
K754zO2oGddrhiwpVsGTQ7SWWOL7edKSoEudu9bTVe+ji8+JKm7OvDo+4Xum1Fk9Ji0ZJ6Kwnjgc
OUjhuOjVMo6XY+K0y0hRpeKGkWlLDr9+S+ylNPKMF026aVXTaFIA95JdPNefV5MFQFS6ucozJcTN
RaIZq7oIj6jKmLIFEuiB7A8j5kpt4HPEyRj/hEQ6n1S5iGcXlfWcKOgpqE6ciPP6HuXgiCLCkfJt
D8eHTSWamtfiSVg6ufHHG/sIB/vo5Gu7SwGlrDtrAEU8q7uXRZZzbxpGwZ+076QQwcbYrHvtoYbQ
F/JoboIgaabHLvrX+FZkAO6HE/KTPGvikO3lfuiuE5YWXl2AzEzYTjIuPITbSblNniEsgqRQmJPo
SfXoMf8W3UuiuReLWHbH1j0NvI5gsFCof0taPmOq+1Ex8Qjqt6tFvFw0BIr61+FBw40bJsqB6MBV
ySyIiI56BxiVeoZauu8rh88jIfXS2nZdIvb7cMCgFTuqDjhjAWP9j2kklbotH9736u6LXLwq6i9d
SIfD5aSlwrAb3VSePPGibi4moZW6P3SIDb6N5mhR9hdDIhxDWPugJWOlwFGBI6RX6Mr1SVlFoAuK
SIXUeWRe17/yuI1H3B2CVG0y4dJ7hVxxeGGMciWIhTl0MMuHeTFS8Wrt+7xamIqGyMUhrq9NZauY
TQKpVOf1kKlRjVaPN6a1aoba7BhZawjWHAPj9sdiAmcUXhJMk9zl5gjru6K47y9mW8OURNcEXx43
IpwmfS6gu9x0LT5yaOmK2yuzuJ7MVCpYjWq4j8AWuB+OGStw/K9ajleqvg2yOF/6EvUANd5etKQh
EAlDxzw7uXFVGYgKVV0QdtomKwz14ZObokOMvkJthy23ATxUiLQNEqTfDgGaash+/EgXJcyViHTY
rjdGffC/McbqWDN6kCFEL+UOuV1rmrtgzlv0/KM8rry+iXg/lMyxhyU29bGeYLxCXjiD+Rp1NKNt
g8QN0UKiQP1tZ2ctdvKTY1HI4SfrdmRoG2bVGzkiJx5/rWLCePCYL8YTfP7hH0LCkGcW8KGLY/7H
5BkHMzjJOx61dmuHVhxdZJ4aDpm4abG2VbERJ4q+uw02pHT5U+6RdrslOgL6XvOhJ2lDsFr7Hd52
398Lybtz+hqwOLAt8ofRRwqVMAvNGaVrWjDs8NFom82HGf2K6LnKt5o0mMaiT+W8XqoKHCZ0S7SR
3F3Iq5OlH9Jrycadt3oYqdptAwIRB7dndsTsVsn/6GjqRmjzldB578tscREuGH9xfbyggyEa2MPi
V9p5iakIE6da8qBXcR/j8b5cG/Lhg8VLZrD+0NCRj8QzfFj0lyAi/seDhYb9d1/qtpgjNEODud94
7rCsYYqt8NbtJ754oeaaHAE15z1phdjt+NC74ptS0pPFmfz9wDuJ2da6qCtTrltoJ5MI6+TXlWdG
H45r0ofOXCrytdD/VKbk5InmFVAxm/mDpGqy64DmlkoLaUkPIsb/gjGuVN+V1NGTIF2QDgoN0TMK
x2uw0IVI8m4BIR9NdsDJ5BnUhH3J4MxrHpg8T7QXvTDzudgZufVf2+IaWZqH2yeskz9kPXJrXv3i
H3x/F+xhznu0eSgXzwHSevScvQnVb96o/oGGWC6gB12b0HsPxsL8b5JRnhHUURAJc7yqmKbEtZL2
YnWELHThYUc29t7hjlGdveNsaQBZ0b+ZxuAJUDFgGrvDwot+fb6K+sQFhKh6qQiZ7V6GIUMRsPU/
xt02MNRinfuTBCIkBlImm+KTVEvJkzi1htgTDyYJZwobIc89j1EgP99p+GhgwzwQqFOaANcibe9k
TMKxUeJecS5SRg1SQ4Lixk9T6pxk6I5B8gUoH/YCquxhADEvzB92bIdsMC7Z3iW1BQfFvC+yNaau
YbRWVq+DwgBSyB6bzPrFltrYTtjwF0CZDtmjTlRjGuvHLNad+qBULishJWD7aa6MqymEPXaJj+VK
lKTZh/VYmbcLN8Wd5uMoOymPlLwwaotrQcDMYfjszPLzXLSYIhr+y+BVMe+Rf0XTnrJ+O25pSxBl
7hUQdlAivKZWVuSUF6xxhudopZ2DXKyh3X1if+exww/dvJ+gGgimNP3bQGtXV6IKkI3fHctNq5Tu
PVqjPBfNkAqTmSgVtiieRoe45Ku+gZmk8xL93UnbSHa2JunvkMzQ0wMAkMKTPUQNqxAbXKPOyn4W
dK/cInC4lk6uhHfd862Kb57MnLRmfFxsowch6ARPXYlGcaEE82+du3VqxoyRNl/WOhRvTvFwqq8r
QqoOb7RkG7Aw2UFAcHJCPC6pezId2+9gnK9ie9E4M1cFu/Z8R+cx8XNw+Clnjjj0OzICCbNBxMxU
R5p2ft/tjjpMp67TvIMj11+J9gWf7iCAQFj6as9ohtMbj+vI5S6sf6PVJjYUFpv76u/yQGxLgtY4
DY0htQ2EJNZ/+O3uRuCmzGZww3OU1X42yzKPgW1bdi07vFtv0hq+Yd6TMaY3dVWzL0Q95jPa8qz5
UTwuMAFDfy6ndaLmgW3zIpYWaE+fdu50zalWmlbP/ACEW0jHf/H7/BrMSRbv/jV8ipDtqCDFHYyI
Tb0pGdnc/cFpEm1ewmN3n9UHRmpXBCnQSNwjBh1KI3I/FGbTHj7EeluR366yMmh2EXOXSMpXFC7r
2rMZFLMWALeJJ2sTtfW2L1jq4Trazb93AasGy47gMF/N1blPYm5rVsijVhepYbzCe94c5FCC1aYm
Fs7nSeybv4x6sRi6D/CulRBqVEM4MT0ML7QgYoKQNwmpEscF7yGXT//2UhoJFUubQjClqwNIAe1Z
GP8MJBmJkDyvl4RD4B/HmqgAsoWpzNxDoAZ+medxAoBxD+aKVb/Mlcom3DMwc9SCA3B9EWP30QPw
mzr73S9J3wJcL8z+GIQgEeLsOTJPH8ZClcdBQVoL4Va3SGgfV2AH9+HXtHVW51d+DxoNE+HTe1gi
tM0hlCAeir78DHhSEMmoPZeXOOf3zbvWia+E3qPsy3q9UUc7kxBSj/v5fxY/N4LwLbHurD7Yn3xI
CivGaO1M8Gj3s680bw3ZNIzqHriWeUXIaVSPIRDLIhn1noGdVTirh1bcFcVuS0MfUgNk5dHDdRlu
JXR7zR8wjeXSjSV7Zn46Iehb75rPpRpzjGpiSciB1lceB4Tj40EUoJ5+mA6DHNqD8FzXVNLIeveU
RdgBCnEYE6VzDB9Vy7Mxr6X78tcn1sq30EgGVZ1EwSiRALhYRHT+9WTeSCsJ6r5Buqp6DGiKoeOW
oyIgPD7j4UbJl/JscmceU9xKtProrDkyO/OAyA2lS+Kzdt1Av6Jxqt9SYhpmYo6TyiY7IS8AvTEF
KofAH/IJk/FiZ87zJlvrIO68GGMrLXHZ8VdYQXmP7L2U/Uafuj5Sm8UvM4g+Hayt6nUn6qEjY41k
7yMXoTH7mS2II05ZiYjJl6LPJHNT9a55XZjVjggAKu+sYhIh2CiGn7w348m+U35WrCDMFg//MI96
WURd3y2QsOxOFSvC2pllhYyiqNkDZgbXh/FQcqTd3L134HJipBX1VGT7Nudgo1lWY1ywhZLgE6xT
ONOZQsecYs57f15efs4PRrno1y9LzGKOTQ/8Rf0azVSvhN58Z8ArT0CEV7/bZy4edQDqoBaM+mAy
ReuhwPMEGj8O5lHE+Yqyub1oDSNFOabooJXGy361t/HXgYTRmLFlUN9bVAnGzRs2XtIdQumKQL4/
Xo7vv/qLa+9eWKUkUtf8ghY5rCPeV1d6ZfSPQnchO89az1bVayfjRwM0VZvGHwE3x7YX59nVNR0c
312jqrMmSPIBRjAFlqtNbIb907/6BoaYqEzsVM/fOIwiFv6emjclU3p0kpi7N9SpnYoCqbE22AVM
YUgw7mwGRpdGpBvBBxgTVVOlS+/g7AjP3sI4qT4Aig/2Z5JHMFH8maOl6hXhpBG2tWpMmrOPWPEo
Wf/2jch6m98j4MzKvtamwt9CRD7NPQdemY3dFu0dakVCsDOnDRgx1oM1xZt/7UjcVFCOMICGXWD2
J4WAnKo1YiwSPRE4uUIJWfHck0reRx444RwlAcIjI4q7iJbhZOYHAU5WlxcfGVhYIayhZeLVfK6U
sUawck/pxeHzEDEg6yU3W/R37vE9sHcJQw9wEHbQ5LGzBoq1ws8gSgRlWwA2p5xnZLUODR/7Lj0y
WuYiRfPkZnL3E6su3dyfMH25wLQHEW7RqUpW+i68KIaoqtPaMRc2aT1beU6fiW0n01RyRsi/Pfb/
64M8/v5UPLsorAYA6PiiLa7d2sH//n8vNuyWpTkmw2lR7rZqdeJT3pqwiAVuJd6nviB/xajP6vSA
rANhbjkTRwyMZXJXOBhXbL3qqsbN8RUzzQxM5y5wdqCLfwi/VBi+asFsuG5SFF39Ld8cxQEttdPY
uB+K4pc8uBzOdNH8YtvuVhsGHiKGK2LmowSAd/dMfMpAVqGOpPByQ141Yj9g/pPrATDnSF6vpsB9
rmF9Ig4/iZqwULc6Uwcx/t+gL8i0MPyHhGxzcZ+I4TTcGlbcrmHJQOBo/U4tT1hEQFoXwRn4ODis
fEsFG+FkLBKJyoaCi8CdoMPwBTd4nQTgtFB3j9oQ26gg+thUcQ774Q82bDn7NkaqYO/E2SR54seA
gbmrCA3n2B6GlNh7Oc86+79BrUyCjqRu6M/wrBJYqWKS5nbfZ48aQ43vRSFtBj1IZsfygSmHAld4
YHAeccHbupfov26LGYvrUsdpncNmgDFb4bNd0QTJrd2q/WX10I1MOmOieR4X6/wv9VN3xcSdqqAe
EOpK8QVtZWEtKBKzkULg/kbDOTnC1CzRiNCRmIg3siKTZGPvK0/VVmhB2RCQ4YMtKoXiYjnkrWke
9GJxLbkZsG0Quo6xarMJ9LPxajwIUkfkjb0ThvoR5qcbEgyIceErC05fabeSEzDvcBWJsAQfKb8+
jzsV23Y2UOhJ/EA/GbLCX8c1K7WmUnyghfgxrnTjX72m4dnsDCOaOc7BlK9z6Bx87vjkC/mp4rqr
2tEXI6L5zs7BKYqTwRQTYSEu/+8eCBaX9eiQgadqAOCvysdx3XCbsXLO0iXg20k+aFpG+ehzCpto
WUl8NkEZGCsLxrtFksdgg9V/+efWlGbExNCp10Gu9JjFMffqBOpzXvU4G/ktA+xeB/yDRvJyKIx6
qRPvmeasGIi7EdtUwxN8TgVzS6D6uRavZKbesqJ4V12VO4ikXV3VF9d4GWXPJB5smncxQiC3islP
qwYTdCwfMqtTxGu7TXr02lEvjtx6fnWQOkGTSkQY+JIfPqICXn+4MXktVbbM8IMjZapNKD5bGyhY
rc2xQFlzCK/1ajQD5Ipu/c0FujsU5oRypqOTAzcAfJWNXFvpRzd2ue5DZDbp5+natGRaHTNr62PL
p0Fl8QrpawSiOH4DAmGH8EjHp1t8b0ySAE7cVMirwda4lmIpDpVL6EY9gIGQ2PxxppQQycVLyt0c
wElSDVjCwxemjOqWVIxEbWmnwq9LBtKD2OwY+SfJPdXgkEK/zRZ4tZ6D1GuVgFgHxhc5ACOu5xlq
fesDbqH4Pc32cRb+piH+RqpxbxEPBLKyemuay0vdcDrZjQXl5xwQEfkvwQJieIkZHx8Li5n5XW+V
2dAtjCWLPvo8UCXigfDayYl8HT9XzpbniPtehwA6WDSR2vJwZ5+9MLAlaCBtPGWedOoAd0lB1Bj3
UU+KkUS3vDBSlNMgeVZP1e48cB/NSFDdkcRe3JrfjUwiXcOOs+rsKBo9EbgKd+kZ8Ae45UuzE9GN
8t8+p+4jZv9GnntEJhL1l0KYSyUPsgQN9ykALuHJGJVl1VU3qd28r7wfJg+pfUyo1DGOUWcSqmav
0pco8qg41+E4Av/Yy/cUsGqZEOU6TnM00bDtnoBsizK/UxB6L/I0ZvYoxNA/V2bef/oFtyBnZgfO
Z6PpZaVEEPbRb9gnliqv39JFwnYvCCbNVT+FuYlVJPrY3ckczUv662hzfBW4t9PlpC3asO2vItOV
blLjFPvk9gsT3jWQCdFF60IZyuqMMvvtWIiHHjsZhm7uTq4C0E/bhKh8FDFay8/zdw25HIXifdAf
nWd/5vErzICWpzVak8kv4uEUBXQtLu9/DW6Zc9WepsevaZjpSUjpRLWECIBCpGlg79kQHOBPe4pQ
Kb0SpXlAsG3//ZXKE+hmMT8oS5T32K6hJy1KZXWXQXSjz+1zm0b+/nEm60DBccrKeL/IbFshFqvg
bbOxbwmPY1EYVqDTbdgCariIl7TFAYEAD0wDcdy8w5zA7xpwAonDv/fV+GuesEVY6q8FYq8P9vlo
InnR0720lI4vIw52VndUVqcfGc5xZdiw+upRHRePQ6qfLqr5Zl6muPo54Rtr8ZDo5QGpCCp9+zyX
pmK74yklSIvh1vkyvUo+pyd0buk5cMEC2FbCH2ob83ac4gxp7q81j1y269+4nMkmO+9ZMkwVSnVY
DOU0xtm7CJeWLpP6Hfm1XA9Ih6nqcnAg5xLYd0fQbYnGUsu7ZxAA7ng1puHEFLJ77y/UlzTGeb7z
yttco36GBYui4zJAP+EYcXdyTE1QY7QSZAGDn82cg49Pk8nPp7nCLTAwyOEwrvyvBaIKYFsP05oL
VeszJZh20sqvqpT9uK0YCmGNtvot7AekJCCpWTbNDxcGOWtoi3XeDTTBry8+7alklOFEDoontRCr
SIrIOYD43ro6oRUFUCHC7nveZFkXNEcFNzxLETmry/8bwZsBGlNFrGBkdDTiomAQCjIw5gRm961+
kyb1Yb0vuKEECZL+hrVTwWHIbPtqXrEl1upeZG6OyNDzzcm7TSkEUWaZ5+A9CoKjmihQHNdwTFG+
arwyLy6MdYZymooGt4q2MXUbT3JaHHUc4ZbqWT4Nl2zV/Y5rTy+CU3i2HO/DtyDOKAH8UfJdwsb4
bJYD6ZHfHDuSOamo7w3MQSuHu+9e/PR0hyB6PUTviA76QlFMFYVJ1o62lY/eOrSkzoHSa0Zrr9Bo
L4Nm6b0tdTPDheDhcg+k04A0quPadefIQdzX2voGYztXYs8lLdOf6kxPx2fYX1QUZVKbLdcleneH
1teHTw0fT/vBGn7XuSsj9Jrm6MSitoZLJ8BsT+slPDpgtyizWxZRplvxolbXFt50GuN3vVoCZY2+
5BeuhOENOm1Twk7cnw/yGdnA8EQVwGKCnHjAv4eBBmV4WMHhl8/JSpnWGeeNTymz9ezIAqF2bPcl
llDgaxkhGzoqoDkSQI2phHF48ctrgThe5foUWZhtEX2xD77kl2WL8gRFaJnRFomK5FiIOgKZLHsL
6YKa8xzPCJeR9gXRxCf0oCUGoxXTPS5L0rqbdvyD05pVJwPS9YLSBnyazTix0RgQ8tOMJ4C11UxO
h+CFYkg1qMzSMdMIQmxUqqYH4clwbaphycB81CT3+lRqUagqY7Im3IKbFaX9F0IFhAQBWr6U6Hzj
c6vOWZv6ygkRKgLSAwCzGCzP1yLzcXdL3IaylOhlaSBu5bITlZtXSCHIWPCuAZSqGbMOlzBXCrMt
5aX/V9LwvUzqBpLlzfSdwNPf7Q4GpCYm8HwHwbFTLI6IfWeEYcVlLqWSTMQ0+A5RIR3KHUeECbwl
0O0BvaLI0s4ocvkOpnbwBBfy+6rV5c3AnYBRg6NmFX72otw8OQCqqlSCltPFqvfkETHDWjZO+une
/5j5JkYR50ZWJNzx2oWVG5q3Yd4rnslllTeLzvVzIkSl+4kCyvMp5XE3CHyQ7E9av9EBw+DtcIFT
leUPQgndosPWdWHfM4ej2q+2/jOmWaR8L8lXJcvuV1chr/H4l5FIiEs2DVFQhsuJP0nVa7AU6Xvk
LnYPTCWN/kBzDD4jdDQnFm2BsN6sTkslY79Y64V/xaNxr/KkCaOk2HjorE4VsZgTUYN4uFOEfq9C
X1rYx3B2sq1Fsc1aOpEgOpVJwAG6NdydjjQ01xn7rd3JgdTpqNZvdw3xY+wY96VZt6RUKutRnDvU
zop/8/FlflqAjVi4kM1PTEY8fG2m5YL4QA4HLVsRaWXEXAyVQB3Owtu1ANE0eOG12evskK9ONirb
QSac3UdVGEUrpFQNcPCCWN/9BMhYeh2ss0iM3rTTfHE+jL4cFC2Bt8PqNLm0L1+Y5IkiFFDkF9f7
dFDYBvRWqUYGOXsWHVZenj5RM+/dmur8q/j/6tywRYh7PwnTpJ8avOgy7otQMWSO/GSrBSNSaOfo
0JdG4t6FmyoB/UOhCqr0i8XkUroo9iAyZbGqTv/PyBVNhG15OlV88q03Z/Kp+XBliSq5Tuwmq1Lz
5KfUm+T4V5NNu3BxRlwIRhWO5zCG0Jdcu09Lg8dqGb2EU6kMVuOovt8ZemqxiHfZIO/e7aQ9ZtP9
g5vnepVIM4XunV0gGnTqAqN4ZU6G0n287xRVtUwofQ0TJzb6YaxMgD4rgEXmY27frVx56rl9OOvj
Pp3CNNDlw9vFZCg0tv18rGl6ubo1QdY6sT005DuAm2xnAWuHGuik39dMT8Wod9M7qwV4RZlvTHBq
PLiBlTI5MhYaQUyCsOsqVXLYcFeKRTvHC+lR3JlkqUQZrWt7G345uwyfIzcoFcysVkQwp3OvtT4F
ZZSSgrnSGC8JpZQDrmJ2uzB8rVDHnwt3aIpaaiensuLQ8o04Kwpents8y6rRCqm8hGm3DauNfp+2
b2HJjQNz4OpsyBCJRgMCrX/+zYx0PaYOxjg2vhrlAuj1dTs4GYju8cmLVBER7wwszv9+Bxe86cGg
9GqcAjT89iXukeWy2YlXyi5DXOVpDmL4tfLegUQEaTrjavlAEOqngKDeWce+12wgOP93MeHaSRt0
8nwRqY2zWfBS3GHdZ00/K0Tuc8IfVxP5jkP5GIUbYiZdqesyrZBEihuS9qz9HkUE3DBmyzLJ7nAi
j47iKTAqdsBh9cX0qdZIA20DH4+Y21aeW8Azd/dPW1y80h37w2mbZpU8r+bCh5ZHSMrIjb/79fgw
2WbWz7fmUqNvZPgXjjnDwBr5bJ7Ffyhm/pofasO90txnzuMVEQ2Xfp3EXPiQXM1MpRrtWOUw0zfc
tTElVGxbyXJFc+ZL22i8lqoy5sUTZiNqWI8FAsDhsmQs5To7VbkkSDRn7f6zVdcMmSz31bMNbnxs
D7L3JbFS6h7CKw8i4/lPOwmvz+0B460Pk2T4S6MRTIwd6lj2Ps+qibaK2H5YcbiEsxkMi7qbd+71
eWrGaKvQmOwFELt8e73cllRjuuOtWLFXc4ItKZf9xPAUUDgCK/E14qE9ceCAURUP6o4sW9l6ugLa
VOyrMZLpir7NM9Z+FqlFSch24qMwoVGK+b0PQnmFinZmRnNV+miItRAVfOrM1KEW40EZLUhiXgBP
dPFI5v6hNqjudBRc9241vH/OzRpwP2uG0B9wuJpFDQ4AIv5Ezbvafw3ESQCvWOFUUUe8v58cubp1
DQ9nAKuda1bk+mF1MI8/pihH1sSL4l29OR4FruS7cmQQqxa1IFjijF01vR6GxNc1ZRPeYnrHw7Ed
gRzWF1iJJIBOPOFYVu8mbT0vGI5IGvqUSexeyUzSRaOvuasF/HTWmdtSDKA+vbRkubVJHSII1aGu
dZFWcW/W63PcKlU1LVKM8SAjOulh+fL4LRw9G4hJrTvmqy42K6GOLVo7AWekhUya7zqWIeF3JkEB
wPriGc0iRotwQVc9kgH9jCWHsQNidwLtEYwQqI2SP2CYSpAZcs2DnpYnXsDihwRmsZBFZmOwvMnF
g0Ln8FzDqhDTN5H8c+f/2YI4F0UgOdvVuQvMpMiLp66Wl0yhkfE+GCws23c+3jxqL16PLgBopFQU
bQV9B5QJjnUt9Ats57uTb2Q+nsCUtZ8ueeWebjWBDJ8T4g7GP3+YwkvjfLB/5icu+UxVfQy5c/Mu
qRvybwltihILNm6qdt6Uyb7lFCosldF0V8b+A7gGF4cMQfcz3DkzuuQlY++pHDXMPlT96JIb2MX0
cQHC2mPO3QqYcs95COK/CxE4aO4OM0rat19O1AufcLGtl8uSVG+vgw5Lmox1/dPBKciPsYm2Db4T
1bvdB0qcxbzF6LDzgjlh1OvLzYZ2rUmx7PRQtQV+0FLTMNwlIQyPt33WmMRn0n7rLecPZclFa/wN
8q2DCJs7ZBiWm9B3nYNKTNmNYA8x66F1kPEQ0Z46OTUeW//C+aaQuDGupbQbAWUY/QNCM/6vuEyr
3dxFnmT04aqBabF2uIw9Q82QffDweRwP/c141taqK15U7M4CBMIrQhUuHJWLnWJQktc5Rx4jMoUt
VJSPslsZwkF83801NsdWvJriIG1C3/wUT+WoLnkrx/vEu1WCm27nkjW2LUaL158xoQ3TTn9+kLdh
jcVEzQ6LkNhAbTF2Lo3BENuc4+q6DlZbtx4lm4MQrTOEUQP8p+vB3qncVTKtqFxnflukoSgma52T
RDPsnTed00xwubbiixUfAQci2rr21CSsi7QXdZN1V9zb8NTNAEkEnLbUPFVt/VScDjyK5rISxNJH
3KqVxVobhFEbJ07hopWZ05gzOoZTo3cfL3MjMf3DhfeptV42hTCsHCRTvvcZiHrGx98kKPwC41t5
IXsRzObHFUXHwdBVeWdRvFSWnIDCst1uhgWm+/4/8YZ3m4qjIHUJoA7GT0Cl7JpyapTHmcIsAz6K
C3mghdBOsnhTDr6FEELScp33Hmana1PsF9wmS544Ck/cAO/6qfJbq8DLOHoJvLTxYStwTPc58FYc
lr29GDCl/g9uSS68O3+fMbB/BawUGZwBI6bwDtT6QSptuhTRwes7HWRI325K9Vp1NR/5WvKRMiAU
VdaBVVBGf5juJlgkvVX5YcFlAKjzJVd+oisFGhBUQNYNSlvvE/NI9EcfnkVZ8q6nbXl2PiG5CsJa
nuRVK8x3VIOHXfLbaxco/q1WmDGHNXpxUVu0yY7OVcFf29Ux8uxoOkBKn1+xgjq8JUmIowOBJ0gh
ZrGvBRzMJOO9r6W57ptU0WcmTNFPqtopkNdSaxIOpsz2izl6gzHLBtnHI4YNt8dO1fYJOmkPeBUT
EsB1xOOItUVsGD3ahG+TRRQDw2ppMZbo664rLbICB/M6PAR+x1GKkYq5h7koHfB1P4foGKrm0558
fzLTLuAh0uinw5+YytntblMm65ZXzQM9/0fwkKJ3327VFqhB9KHPoCogxrxKWgwGGQsSS8oU/tGM
NgqIWaLLzWFh3n09qA7qyexuToR4m1bohXFQo+v9XCWUNZtmNEghyDVQAk1DtHIpR6PX+n2tJGIo
8LPvi1cE6FluBAmzzgkWvHQIic4LzyB22XC+yLRcNwyUNmZV2ha/LvS+c7UmZLFsbE4CzLViVyJo
8LC3ghW+9JUoTub4cG3tcHVvAFeR5vJ/mST307ik8Eo7wtXmqmo1RtyE6HUwYXe0NABDG3iYrO0d
bm+CBXce0vp/QBvYsGHsf6LP1nXGX51iRq6DlpVeuK45m2VaKjljUHMCb6SUrmMo6qrxnkHh1RAe
uspi0MMQsqHaVcqzhTKnxnTQ6bE1JiUb7BUxrcdyNq5ybbqHDRhDaQLKFvTB72caeGaF+Xq4rUUB
S/demAIW2jSet+t49DRSTOLmGFjxjYzjgDYGab4AohQsPVS8fLb9N7nHh33Nqp8r3TykUt9/PXOp
VM6fLtWHVVrcXPBeKbVkD86snLhU5KSMqek6VVMSHMl3tL4iZyfXVNqWMEkDy4evYgd/D5I5aNKl
nBCv3piMtDySROLs0nRAL+b2yQ6qNPPSk4mzZa1NMDHUsBK+h7Vx971gXF5dBqFHMLhuDp0WxyKk
gT/uCPGwyyOPuWwZ/omElZGb7FAaV3wwpmlQnuy6K6CFSH80PI0tsmtZaIpPY+emad8SF5W5HIU6
MuAu9zgErB6Fy3qTKvht7HTOatpQz5cXiqmZAFpoUMTp8VYVhn4oEzf39Oty7xaxVDrl6IOo9jnD
b+MMArMIFN96v4Z8p8LGqohNl9MFed716p6ZN9svIIKfIB2SrWr19IDu2cID0/D4TfAuUnlH12tF
fB/4Q44hWzSPtfb9OL12lRGCDW2U1vxNLaWxnFnwwSqqI+m85TEBzpOHvwWqQMgJeT7jVAMW4wus
n7yvSbXEkkxsNUL7554GYivnfa9OXa9Q6dCWrnRl1bKrIZCgUTqq2zkjuW9y32wSaivMlENHVPLE
S7smtY5W3NP5e3E6+9KHNT9O1IrcPBjaOtoM0QMWXLlTu/thR430DxiZTj8CjXkhpEXLZlBTUrQf
8up64NP0HtX7VmC+3avMbIxMEkPMn7J3Hh6IVZY1YNinSoOT8Qa0Qdpp9OpQlo3t6LCUOo34DUmq
2SgMmBxZyTev2WAxCMPENbVoM4Rmwyfgfplc3/CxjztTPkBLRoJL2hhyINGtwkl6/g3Djh4L0opk
JBfeFX21M/4LDHVq08/EUhWOs9HBciuFX2DUzbBPxtmgv53dqgbnbAbDJgpY0XUJ4yjP0b0BuBUB
6ME8fLniDt+bFOkVbqgNiJGX30OTNnfIvzeYqAsP9CZBI9IMjhBSDXAqtKgd8Ro5Xgw5j1lTFmVj
xIwCQwDlANv4sXokUjkUvDTnh/bw1cNgQsS5Wc/yRnVFMU24uXbCgXUVQWCW0ltd3C/lCO30RwTP
b3/d9J9RhIYAYVNUZFZeGqR4ToAePlBdkj5fFoSLR53w50oqpcc3RMyRfLMLxi4q1RLZDZMro1uF
sEbyBOTPlibOkTTG2fXZ5gLCol3dcpBRoPlwLYM7AdCLaz98rCIl8mRniOZzhAw+8ms3G35H+5x0
57V5FGf7b3hPasFTw3qnaauBmqMaA3QEOIbCpDUYUH2xzOt4SkfBbmREq+RVAWsaPwP04RC+0gsc
VsPGHE9n9EtwLe087S85qw9QPHN4dnZ04Bsk/bF3/U232ploCLP/CcJIXHluOPxSvODrKEQwHSbZ
UeOSjXyXiX48ZpVj4H9ETqsQrfBnNDE9WBNOjzFEH0Jd/nKh3Fc3xMuhCuBUB6gXdjABkmNgNoz4
RtdPIvTQnHi5ls5sZDXeF2BRJKui3r4HdtggIU7to4gm8p3GR/po8wYd6POD3n97xr51//KDN3Eg
MMNhWGYvbOxrN664MKqVcMvuHF4nke2JOgOfUR87UkXaqXC9tauc/A6qbbq5+s9I5RjQDMQ1Jwdi
VKWCWLGfXGt1fmqemWY3HjxCgok8zRYYDNCq+GjN3dbAFiTl/ToGBDMkVkQ57TZf7E7a3eRiYMEo
yPHgbSv4eFn14UqhghNul/aUNfIOjdkWuoGo/PAQXUJnGrKZQC2KIZ/npNHkyDqhhLzBrIfbaxOj
K+LRoWzkUq+FaMFCK/I4ndS5vxoYUqDa2UzFgNYvWscCXPOcQWpbz+nDQtop/0lxaj2q/nGp0ZkC
UY1Nh7G/XnQJt+bkRuDbgWnQoj8FnjmkeOQXNqtAiF5Ck2WgPwvF8AwACGxh38dArBPEMFmUOktb
PmhRJmcRP8MMgGMmWihPZUqrFXzD+IBLJEyrEjrJ8qmgCr5H28drR0ivBQ9lDoWytwQwmlFnaEQY
2YPi8qrssCZjJ6r5j/nE5Y9pSHivDSCx69s28d8N0Pfij03pOIkIJe4pBFktlNqC2b+j6xD2UIru
FYr4kdwhrRRv8T7AEUHm1FZ5WogKAHtWddWfGfMTGchjk3BcYqfCGMaao9s+djB8rwsH58fcdpBs
oswxq6nXh+P5e1uyc+p5J9ULI185l/DCSczOew1NPiOSFGmJgNVgCoYS81oMv1MoQXvQmHy/gSbA
JkwqVbtiUXzn3EqL/ObWGme463i7Iok75JeJwmYm8AWP7MddJK27JJnixK4467fiwUOPptBS7/rz
xKShIIHaeGCvHESo0tSwdPLlOJ2uhxkfFb53zlDnIi8EjQO/d4hbTvio0JtruJi9AnmwtJiu+jWj
fdYLS5zTSmwLiBcjHYfiUnSvjxZHRxzUj/WZEAB+zNneqyZtcKQi2ze8yl00OJ2/PaxEEfPUNTfC
wAhE6zMdjTqnynfD446pTMyVa8qavS7C1HfzlL6fojWVC93guu35KtWbjp6dX1NUDp6rEXPxw8WG
tsLn1QvVFblFI/b92aizwDHbtT6U9iyo499gqiDs1tAG6v5JK4HGXZvrYnquoeP+Pd0iXWeAUvX8
CvqO9O+jQsmd9iHrSlU2s1jS2DXAqWVMzfsTf4VmKv7eJ4lUoUD7TzbTQlzqnWON4NTm6JtHc246
qo1IjNdhWKTkRDVA5dH2frB+xJaTFghYPPStWKaJhjj4lElNnzmiAUm0PHibfsurYgn/xny1yeay
0pRqcwrQOUDAHs+9PyUGzbgwbxMtptlVfSG1r51a1Ko3PLKkGbn0Kz3niwloj2hPnb+wB60Yor1f
yRxwbHQBgF74d+m8Z3FCEu/jwg8lZi6alban0xcVyXcQe97AfPwE8hpAMeZBS3knoUQjCA9wwHoM
w9Dl+vx1fgJUlx1dwLRhF/GMM+gDE1hKsfg0V9APOhLpcw8BQh6zTnNCRq0AIWQvB12iB0nBPmFT
EcNCEePdqnk1S/Yp2bj37xxdCAKs+k366iyOZUR18KST3wNeHscxBRzjZ44tkoFE2WbMrsVXksZJ
cjxZCrU9NxPhSkJJulSDs9DBzhTn+/oJPQjhG9xxv5tpOxvgy+qRhjfmOhXfO7F7S+JJqMXyK0bJ
wBSRHIG1BTNisLjWCtAI+uFShDPqDzo5VHEd37Grf6kYOYvvUpRSjekb/yzziIafg8P2Pc1JUyx1
PVSPCRpULh70vICpHBUZggtTih09cvaHvby4B5gtoujwuYplcXIf0r2ZiGdp+bp2hlj1oWKGceHd
UKkOPnRv/XCGA4VvUNgbZdBjdlawrYdKKxNM95bWcaoXUGRrkwlZxPLj8yQxdMQK5u7we5tdY8yi
l0w3jppvbJDfjAAzB0bqPA10sLIB1KwvnW+ISe9a6+HIh1UqwsYnIGIcsKZDACGz8kCS/YM+/ljw
2IY0lHi+BEG+XBKwrW9uN6tvKo5wl9uiJ1WPsN4J0OVIintVk2IHk8ZR4OFLBTODrQoTW9QsYZlx
zV6YqRwcSYIuUAhBpDX/SPxslhvlwtf4lEOCXdO6Nmm/GxJ5Peej1shq8+MhSiS63sqQOgfdQDY0
SH3upKGHa4Fhi+3/hboBgzRHIZstKG+SNgmEWdalb2IHGrHMdB/qNNv8NRDu1HTPnCHIKiksx7P1
W98oB4bvwGpftmtS3N+B7STwp8t5IDA4s+9ANtUnm0XuML30zHlg/UdoTt+coTjVF5Zn4YEdbYrq
suH/t44IDlFm48O9mAUTortuPczuupgdbYWvBZkzt60zlu0AMY9cEkj7CK0yG8ndgxEAJtOHO++2
eo7SVY2BydrYM3/I8Hi2rwAWbgHSmtIaGqZyF7EwsYSe8rw2/ZArTETPykNdiQuCTK+uBVRaSSSZ
di7bX5Y7yhlu9Iyf1zFqvkGVfI52VT7lr7ctwYQ73r7rb6ZVExEKV7dHqk+B45EVzPaHs1e1gQ9o
EiBsQZZw95v0P9ComGvOZq3HTwqrLTq17yXrZDxRj+Tgg7qc298ZGOhNlDDGcHWYQy19T1QLCVj4
NTXLuyVVL6ilREyroLSG+bSlr7WYffHV5GOFyDN0E1PtfBHIGu0bCMt2i6Oa5bUzdRnDfQYO3p7N
oxLxUDNbbNxWZ4sJ0jWRa59tRU640o5kRJtqGmiW73Ma8eZERD0b6GLCJ4lZ4475XPndYZpIGaoM
A2VnhOnIW886B7E4jO50o3JW7KnePoZ2KslDm8wiugLSuefne9jfoUMkmqjLxEfOzrXpYTYpomiM
m2y9niPMhreLzlChHvI/I7yDcDAgQ4eP+RlhRwvmouG9uJ3HTa2/d3mg+M0fqooBXxwRlcy4q4gS
Txh7Mqp8hFTDbAF/s1/jQZ42m8gMUnqxxmtAYhL45dDfnSXUVcoBvK/AbQauPp9yxzHFAyIDEGui
sGnJeMDD+j+DbXTlz32zh/WqOtYODOBGmQJLDacoxyQTzFarOJLD+v7TgWHWWbMMcVvZ+X/O4lsB
INfexVS1tCpu/G62EsNeQhUzobLRMAuzXC+b0g3fhkKw4Rt9RXfEMwN4bzINd8u+LzVTZelG5iVx
JNdeqcHOFe8cewM9vQIi8jBKzdXtuMsg/LHR/f2uSO4+eaebMXS7eCA+Iw4TDfNx4ZsCVEEuM0rK
xcG4ufuaTlBbkbM/uBnlSz6no5Mqc7mTS1g0IENQRocbjAgWwHdIgZJnSvE90DkmJl61ZZbm9pmD
3/xdR8KKL1ol6sj8ijB2afGuUekXTKHpJQw4xJQNmAmAuZlz/wkZ0VYJR6XFnVApJ/6CTNRM8yB8
uvGDzrer2M98ZMS+ZzOcsnYqP1KZl/PoY4kaX7PnPWfyApYJu2iz5dwrFIpIN9spmQK4r0bZ7QIt
7mIbsbYy9+DilA/dB31c1GjlvisyTf1pNnqRyUrKj3Wr6rFAiNWA5EkujVnHYf7q1usfCRqfBSFQ
u/VZaWT8xyRqNfPALj0hwYeVScTyhiGFQHtNwRN0Vr9Ypj3juvZU9qfhMHF3T0V9soO88eAVyrTf
FPUFYRmLHhia2PSB4yf3Alz0qpSvXyFWUS+EPnI1Gq/iOHKlU0Wx0VKfKKJAqUjnsVGiUwfzg9y1
xKV322pNRpzg6iSMZlu9WncqrswjKvl7yCctqTqY08pKNCUk/SKV3+6TxuziAbG01+7jQFIJOneT
2qwODwfW+sOn7ANfZMTTuDAixwmDRkcVRZBIzUEfjzoJdotoODjmPVZA4cOaBn+kfEAc3Xc6n3E5
ZOm2/6uJvqmAWwfi5Hcjshgc8NYzV6788h9U0Y2CX+BtfCBoHkVf6nksrRXK3BvYVZug/JLgtyv5
iEbPISMI9cWfD99jX+VDmQ4Zv+3Ai/yXI45+b9fHmYsouwELmVSt/pkWoDCQZYjkHNOWGVJ1LkpX
fcA10Qu4C7zRG1unlOOEe/JoEUDacoS5Qj2HaH9FP+ln55DqY6uJk27I5yr0fEEPBzMYey5id7UL
EleL7QDt/7vrcGYYaAIILx/8Dvcn2BC6vyrIZFhY6MtP+Ok03xK6QQc+5Ng3xgwk10T+jQbmjRZc
gMtSgiA4fbr9yJ7hxmjaGDB/nyeDH812nLzKKV9nSdzkurXPxDV2aRsBTrqiNcV5BVOwMc3Wl+89
xpSDLXRoss4M68FJF5gv2/48ZdG49Zo9YdlxpyeYOFKnsjvSwxKBIcrdH1zO4NtBrcWfBHVBk9JY
5zx8SoPq1L+IZlRn9MJskAkdMO7tQ7mr18xue79ucc0Ffgw5KSqWedZ5GW0EZTVpV82X43z9xr36
harxn+4x7OJaGyjAcag+sDhYQotPREF1sV00vost+Ot5nnKx9tqJl7wVqglH2t0iNSlsoUud37np
yQtn089eQCSc9Y45yyjYvRuQ2n1dnfzf/4cZCGrS+CgNFLB7Q/1IlmR1cGpnFI9M3mpeTUD1+Owe
kqHLy57L5JkDRiIWukmyG7C2q7Mz0qHTBOUvAsFTYjNThRfL8cNJHsErT59Jvx+phIO4EGvjaa2m
FRliYTQIR52gqPwnl8zXpgowCmRF2WMkgz5C2yHtYqKArqGgf3mX7wBEVNh+ACFFMmzNh4dPAMJf
WVe6lVQRDSQ5M0yT6kC2lfIbEltO7y4AgqggAwP+X5xCnPH5XNK+EqP+KBsvygtSaK4/vlOzpNk7
aa43UzzqUUMFhiYR037fA2YX+YTpqCiNcY8JKxQv3WQlX/xqcrcsofJaeHbjnYeQ189yembdcbQ7
l7jPeLGMck6CC36OMp59eQp1blS/0nXLg4nWG6SVsKEw4ajzUt7N1p5nErPCQ3c56okR1HtGPytq
CgLSPFcZZ2/oErhEPky42IMUOzboPTQFQ7G087WdijvlC+e+8xn3O8BnhMxR5kVnBCw3n8G1cx1l
c6TcxVcEcClO9PywGcnvqndLkyV82Rx1g3jacx2Sz1hn6/qmB/PiC3WNJNvsY+U71x1PDXbvNit8
RHnF7k5kvNJY5+/DWUwXCaB2V95RMYrrSH7iheB1iCVsaN/J2z0fZefiW3CalDCAbQh7VNylgyip
pW80pyL/bih99TPMwTtLq6EyVFW+y1/4gytTLS1dbBWB3GYCHr3kWaZoSJuBMj96x1SgjOEehlBQ
64JgZmaloUhvDKAY2J8Dz28Xc18wXh5I1eTwMEmFe8/1vLJLRWVT4WcOe/UPWIUEGtqcuYK3tCJR
VR5jjMdnQblOUH4XrMYuE3pfCeE2IOQSgwHODrF7IsfrgoLk3OgU1zon6bm9lpZZnGkoNDhyJ1rM
cWfyJ4svUFjAodzPIi/CRQv8PPDsoNgu2bIOkVhSg+hrnErI2x1w0Js8pM9oPMBaZ6MXlEddEzmn
k/8qvkwCSj5wsKs1dJvYFp/bUIW7MOFgcz1E1L+BDePOEHgRrAFjS4FG1HXuwXuooyNUdNayfO7o
D44iAOi485f5nC2glMbNTkFhrlAn2ky+Ircb73TXDRu/VyefmV5zE9aa3RVU5vxuoDL+08WY/j3o
rOmQyvhxyPXO45/QPkIY2/Uu6VhnqmJG60xeoR/zxQrfXeEMuNX7tl5MH5Ud02HVw7QQ+uT8VviS
zXiz2QD2FdUZNAE/AwtvD7NVUNBMhikWP0LACX5a4svJz3dWT6paxx7qHaBodZb1iBuCNAoz0W54
okKANDj7xNuEfLUoc/3vruNcDjho1Sko5Y0xQq40JbL05O1MkErZtbJZLgVoSziLe+yFtdluP5Cr
dNrumHC3mSnMCRgt3Gf2OWHYYZssxpV9chh3Y337kbmfZLwQqmLqh9XbM18qAzpuQEYaIDBKOBNB
brGwHQXO7RGXSzFxK96MhMZjFtcyelJF7yyii/tczA6MueaL675Z0t+8BdCcgH8C+ecR99ByN2v+
UiIAMmsWhUDkyz17ykD7v8UunDqWyrKs9MZv1I0p7ufQjuExaYpC+B9cL+4eD1lRbTraF4M/MC8M
XjsxeXgf051rsbqCjDLGssC0KLzwpI8VgJn70AAYmTK2A48TmC0+44tXnQbhxlTJnN22s/2joJhr
IPrVA7HBbsTdBDYlCpEhICgXgr5wEuoFkXsbOsa9e7d25evEXZJ5G3LLsFXPrxdmmxPJxbToafgY
zVAkabxne1eWKF92KAJGJlQ3enpAwxWl+GI094pTXHCUhAOtzh35OernfOLT7GBQZhmuk33T0zck
XciApGG0hlYCEpNrEBm69lNDB7nF7jtg/cSn3DoWgdSiqI5Go+gteD2sgPUcRRwpOropKcC4QRKu
zpVCQDlUwYhuIR4fu7Z1Rjf0YsL/vqtfO3SbB8dILG/pTzOSlPkJxNqTt1oDg4aLmUuJ6mZGOQ7X
DOJjBW4T/+U2CbEt3gfdTDOwW8c7E9zuN2gH5AVgLWPYDZ6SvRDQji4L5cJUp37Hb1EuGx2RHgSf
463yXKTucFP9O9HDAf2m8JJYyTfei6DkQt5tANYpRgzyYBn92zOYUiOBSJdmXHypqm0HyJCTcH+A
TiELAHrYKg2RvHkEVJ/+S6zEpd7/NJoPNq/tebm84LCh4A4D8Nwjb/LYpQXUFGCR5GRHPE4kJ+Kx
TCVmadN/lu0+roj+BSbr3wWKViz/FpV6WLE6APOaJz2JAvFrMrKpEbZNWvYAZC72v95fiRCmzB/S
F2aLzHG2eAMiVoeRTJJ/WmwQm22k3gmgwGfg5zmymvVw5wdu0tljjb+/yno96IAgFjI6yzjyFYq6
L1OjJ70PhVOmBaLaJWxyiT1Ud2C5fPxaQP+ULyEGQEGN9XGwaNg/eG7eRE66t4wnnJrNnI3FtP5j
Ma+unw3TBkPhrgkitiPXamystKtEylimKVEFgGP2NCQVMW3t7WWVqPCXdyHRSMse4qP/nRRHPPVe
L+yrF2A4RCdjViv3v3wYsrQyCk8YQhXClEhseJsK/E/3RZyQIKempJB95NHSj0mq3JwOXsXGSZqD
VSemx7mr1nS5SOHeENFmV/KbDOSx3QbrjQbBC8tb/2NkZb9Vg5meG0ZZ/GV2JCESx70vqiq97Kjx
bC3tjDuMaI5XnqeQaPH1528HLZFpr3xO6DwhhK+pCq9piziPx0qNqzVD7odtG/2qX0sLa7D7a4EN
gVKuJHTfrhBE4KYmxTZB+dyCln+rzjhVJ52IhB+yUiBBleUvS8lE/i5aCmDv86ci8I5vyIakY067
ZCaRyZQ356Fkf6dKEnlvVJv9edqV3MR/q56SQqjNIjwZFcJSpNGKYrXAdBL88cy4m43hRbWwi5zF
TGUbQQdndcTy/7QYVVwpkZBaaEZOu2AVUW/Fcr+yXbpsR46SUuyPJOv1qWaBtcNzU0XYgLdCW3S+
6GG59DVrGOGyc10H3MeOurIg45ucQrcan2JKC5S4HEq0cMf54zmSJmAjG6ZHdeFGhRufpaFAKdWK
B5x+Dr2fCNxU0Tvx3US7rosPRgTJ7D+VCG2tticueP+lbxNBVMlnmOW2vMRVH8nJbi9ppF2eXTrI
dEDg7nJXCSBeTE2O7YZ4ajQf0mc12TbkZRX4ljKKJuc9rGsr8YJXcx8jPcpX5y1YfoxJW3CWzSjO
rAsR/VneatuhUhKhdbWo3406p3uBxyZWUMLvVHRpU3xqacuU7kqDdVx/X18qeXvzXu5FQEmxOUyS
IFiyRD1+JyN0OzjE1U1rvbhUrGRPmW9Xpx2FTVHtK3ZoP4TNzkTBUeaay8Fz8VSsyUaxAXIpBHv4
cBR6/N7Vt0lX74gxjc+EsiHUohBYGS2fk5u6AI53YjZtyL2Tf6ZRhYE11Kr1IWwYqtEZcVX0KU2h
CbNzqaZGHOLjDh09D+UO2mks6i7g2HJja/e/j93XJYGVIaU0a+3+ud+u8PwL44XTE6K6QTxzWEd2
URsqorvvFbvJuooHKARA4pGtexFcf0bohC25QsyMnF4jbqEORoijX95kBSpAEgbv4ZfFbSejG3Ko
jB9ABkg5QyrLsl1kshBD2TmeC5dN7w6c0y9saoG8awwtaeZkqFICCe3MdT3wtra3umA2zrJ0jFDK
DHbm1MfeB+QiJNFtgxfdiCKQmfCfkZ/ryMKKrKPAP87ZmqCitcet0urzdlblM64o0J1xPIInvAR+
rWIIwPNFUUE7ZquoSBQRkJMZhKAj8uE5TG0NxCometfnCmttf/y0/TUgXIzdnu3AZAgz7EBxE06W
NavklGSFd+u6NwnimoUTFEOZVcTE7Rh84QU+bCAZldo2ZjZ0tqmlQ7apRjtA83B5R0oCcqNgIJDe
iyyeaUJK6lfwelGJ0wVg7pdI8rd7LNZlg3EmNAWG1rI6yN8kPzCENP7BP+xKmXiOP+63ABF/e4zC
byNrNXGDbsUBotSAMuS3mfmmZwVZ07+MS0W7e5o9WLmLbh96wpzZHzS4IRsTvgRLYcxBS0JXDUC0
7sK8uBAf8u1Ke03P9D4PocGJO/Tuh3Lm5o2ljNtum+2nAt5/7ia7Op3tXf6TscgArMfUVpYONIwv
eo2IvUtGIDw2E5NS4BOhOxtLekxhGbmKlJVmlhwdyc9RhK+STrbll/yC7v+b0bTi5Nl46DR7YsnH
Eu32EoUVSvT5auiMqTVyonqwUQpYMNaE5Pu8+zIwVe6fCWvWy/+ocgXDIzlLKKr2Wwxgocz+PSf9
qXhP3ZuEkq1le4ci2Ddi6Y/3wCDbLOkD5W2P1gLo2ofiJOSP1wnWJB93lxtFLtEyTTOPcXNXx7/b
pRY7ftJagk/wg4MImb0zlE78S0iIAB/as1hX97ZWQ/JJAfuOEb5ovHsyMQsTOe4oK6YtToS061oQ
K/6b/5eXPr68+0lPA09fQRP3tKTJoyL8AHLbn31T+4nmCdyAsNqTQJymlGNDVIxX/ZjW/7f39bGU
29J1olNFgr/Rtj/h8U4nimUmc47kiFaaRmVVALBsdo5vdGiJKV9F4l0IrdvEpS3NhO2mCTOi81PA
Ki4FTteYdhnoAHyMnk0t647+T06kLFqQOwzW5jf05FL/acA++N1yfA0QYnxLS2GnwI02yNWHjzrC
7TfNLtP0vH4yga5q57WUL5za1VD5K91pA7Iju161odMQswcHEuV8iwOSqradBXa+dtPUv5NZ1JxN
Y8JM45YXcxuXCWaadsUVPfmm8HMSO5Oa6uPB5kx8lBH44AFjhIupvjMsSevPAzqagZ1vq/GGbVAj
0aj+3x2ueJ/jn6VMSl5Y2DnzW8s/xZi+iKl65/XkemSTQ6qhp0vvKYwBo3rKGHFit+aMRK2/Qj1e
vk2/Kps4rHS2TjHiMk+bET8fjChMQDB3vKXeqy4CIsQdykESo3Osw4Y/qlMeIg2OESOdZO5gs6ZP
l62wb2hPAj9dVqokP9zPWD6RL3D94ugZbf9QIoxZRd14e90L4d2Ejr43F/fssKACgQDRCGM38oLk
C34u/4kD5vukROvxPx7ZnRsj+kBtqxlbnPPCOqOtQbmu96m9LpYDW7BI0CSW0DEvNsg0Ww+dWta+
D6AFnBo/uMqAQ7YnilUJBoFrrWEHnOSoST3t6/eVsTvcLru/jgWbuO9QRQT6wSTYA3wn/9MEwTLO
NJ8BkOrYAIJR2OTNfA745Of7qCducE4aGqpMhrBCpopXayHAIvXh4kgK5XYjfVelhFPHEwXew5cK
zg2xweMVaRsj345EwjwqDrOtlNBO57lmMDefI8LC23C3jztoG2IobYmW+L5HbTGPNJ1vkOwO1W7f
DtIj459rvE2AuSN8g0n0R2wiP1/Qp2+5tAvuqKdlR56yAecmA7qQ15YG85YA6T/3P7mraowgEiUC
r4jpdTHk+VSiv+ekoInnIdcw5rU+GeUtT9EmXyNCi2QlUV24nupWAArtmOG/Q8RuEmC2w9weimMA
KzFXnjxTiY12aiW4fqbRT2gECzAUGfUegJN0iBw0jtripiPA4pvJupqplg6m4Cbra8GJZwRt0+B0
V8mzFgNUo5D8/0dMD68LWaduIAg+FnJ2X8dn7Oni8pyW3m5uIQtTGb1M2yg1gVfhYvvQOA1lmAqU
qj4pDxqA1KpLE6GD5LFktRSdDNEbQE7MOOSOAEa+iMWzG9tpk6ThguTSWgEyStY46/ksN45IrjTy
/oNg4UAbls/2c4ZzOfImrDoRiBk0/PYahPhIClFRHLcTR5pegu6Z/rROpvKqiQBENQbB5omepIwz
JdlIPy/SUcPhROagUk/1yx5JTbkivU3915VLH08k8Bk+Tz48wHgcf1F5EE47VWqX8INjsWdrxDob
+4awKHX6EjPjp9yqIrAs3CcxqT913Ex6V44NWm1Fzep58Kp894iQsSMm/RNC1+FWislYRiclvglx
2kW6TqYoEYbgXF8h1f+d7GGF/IkA5fam4FzebNB88e3gHXwXNpgNOjyONEawzuH0WJcKFWQdnDFP
Nk6o+Xz4Bl+kxsIhVjlbOXKMlVmuX9dPNgJTP+KmXiKMk4zmfknT4k6xazFIZQ5O5L7hnHO+z67f
Q3BySVg4CZODWr2nJORkIcmb8wcjuF7GBqspyxVetDBAd22NlZ1rouKi9CpT5H+/uKDSSeVCLDFe
FhpFNxUJnkRkQAoeQdKLjTTKXythXoYWqb8BsIaQJvfeAZ1+eqgb6xhmh+VwLzjx1RXTkO9OQ6MJ
6hFIlZnj2agENB/CbViDCxfxNNxBQzt7jUf0x/Wp3tzK+axvygGfhedInvMQ4EAN4fOS7TveaCpH
x1wGzZU80deMxIwdHfEEoN9p6rHOgrTPX6SwuSgoTHYf0XseZiB7/UMaeKC05Z8yucx7mZHeCcJW
vs2eEt4zv2H5gYAlqqfZ2f8WI46F5bAnEfcjoMY+kqXx0Y73rmVr3LCrhsUxCiA6bGiSDMrlviH4
Ap23+Uc88/fLAJrTUQVNsRs7piZ1PsJ3NYktljHrG4Oy5ZTy1L2A93DC2HY5LEYdELK5vGvRzWL5
ZZ98YfgXWiEfu3HL1kZ9AA1ucAE0qWfEkb8hAionDVC8DDUs0Bj/Up5yAr2PO39uB3zAJVjAonk3
q6Nlpv1CU6od9Qoj2ak6MdwHLqjcA9kBJ+jvh6vR7AoAzsuOE1h70QT5krB0KMmPB1jEh8v6pLzo
j9OKWY1mKJ9JR4nsUAOaNFaO91Pv3T6jqmNRqXZr5qlnMj6IEb3MwYL4ODknzTqFxW8g4xxlDYNS
hMWYxNjynmS30VEgBUmt5AH9i1Vwc24wXFKkVD0DnIEJu2Tk7t5vjqy5fgNQapg38Ly/7XRt16DC
V6yXgonrUQNDHsIFXp7gqPlHy2o3YWZRDpkiUYzU+DjYnxj05iky4VMK4+0WQAks9O8CAs772URa
v0AUnX0IdQY78GS2WQge/UPnoJOemQgBdZLu+KnaMIucC55POIxlh1agaiRKtVmsfBwXGXG6oxeQ
lYPaXkq2N5N9Pfr4tx8l3iI+ot8vxJH/DgrQtaM9w0Osn9Cm445F7f6AYdXjrUYsLIrWPL/gvjWT
NK/e6eVfg9ZrAxgwdhfI3ZAc+JleoxQ/u+1nY7/FGY5on6Mf9DBS6gMu1ymEOXa0OLHk1BBnTw1l
IrSklfv9LxWUN/q2nVODMdSdwerdGkk5xwSi79hhSVcNuhDNc/94tAL0QvMcWlB4+jHgNxbOEJw3
dCf/GZ2DAq0UJkuKqspOlhVu1nLXpF+sQQoLHGRnGLVnIJ97YScJvNBe8CPt56H8nlO/ekgUgC2O
SwTjHMRaj8WVXkVWUsPM2A+3ZfwlwyR9UGqoq5w0N9HkrL63VTus44pG5iFBVjEG/Q22bHGijf8T
X7zHtWdaxgZ9SFTQd/rY21G00G6vepntNe/qX36UhTV5StVGCxT2Sfd3X2iV+8DMOgha2RMrUHj7
cuweBvgQCFxMAGjij5dYIvEnJ61AY4VJim/QCtOI7zdFwZxfVsFZ5Uy+XHuuZGdfU4P3sTMokXPe
Plf4k4MBOE7ppFATZwhCsQC6Q8tf8JANAGodTt/c15SF05inJH2R6yJNVUSMoGusDnrMFpJKxoJ+
VfaMiV/98Hf6aw3wApuQtYfj4jzq5dGj3cuw2YAmbvID+cMnzpYzPUQvdqBWkNiq+2+jsSAZsncK
tkRHv0Zm2idgrlLoYdARKPhvbm4E+3ZEMXvP4Vea7MryqMGfcUuygMJMwCWkwq6jHFHxXRMa1hwO
wwLgH2QIlyRy9YS47JGWKkmrRqyeMdipuwFlE4kKrjFwQavwI6zUugNdDz49O6EcrGfH11uWPruH
dFzKd0Fjnnf/Gf9obzXFJvVvy7MHRJLc5yuj6+AhU20DIeN1i7DROacupdLAXVSueN4WROcgHAHj
gUhODaNhgtIjqExPuu4sm5YzfLAntpxXT8+ub62zUK9wWbf09CNBAbfQ6tzGqDpJK5kiz3VisWkn
yKECYrjOSXzJK6FZ0JSp5ff05z6Aj3HGtukVU/MErqXqV42Z0mgamn+M5CSmXtVyUcrV4B1mA1uZ
pC1I0n6c95Uvo/Ytve2LGgdXm6T+7ulB8IzVuEqEI1fsz82Q4dtMtPv9oADlPOC9z8GcgJiAt8O2
RYVwlh4mg21fiEO9e6jkm0dqaldw6ziNS2y+KJZDUoVOAR0mw/OSayq2GpvsAGmlg2DSa7qFPaY9
cFkIxZm4vTLmTaf4F4q0Eh4i+L8UsjYvk2ot/lIDhcYZme5lZuws5b9PFhazuWRFR6fNFLyemlv+
Ibv7wvqFP2zNhF0FEisXWl1xz7agqqQOC06TbIG0Q0JPWt7Vi32fx5LXsUVHbT3/wOJgApkiLoF6
8T9LtDBHPXN73xMt9DUQE63PflInN3Bs7IGfauiW5nnlcsefFTqIVLpNFulQAAsX0oaOYzU3XazE
VnUkGWBoCoMwkY9Kiok6dUSjFKFTq/X5GJ2QDSnkdbJsYZfQhpQJ3lSd+9JDdR0ewkwL87tEP8Bk
QkzDO9c4RJR8h6DHaDwO5aYjazFK8gUYVF5oPjtZYxX+6SkKjYcVrL5SDvEKPUUxBrR8kqECgXte
PKFDwEA8MmVTrBqpXNmaT687rMq2/EjIVgkYlswAAGw9tJdr86LUb3CmUZzYVagvPbzJZe76J8yN
uS1BDDxZfkwT3CHdr6hB2Kjfm6KBAprWbE7s7+yL7RB7qf0XoAwm0u5iLxKGAlhsO4470jaWEJtx
noHIA6HiW3yYQ13vzii06T+w5ARtjp2wcm+vVp1ggM0ZEV+NYxlu1Z7Ore3aFmSbc1TTFfrFbC66
olr5oBsQbO3yosYoK920mUgFWgXBESb33LYG2G+Vm1pk4V0YIFd8aJ1kmlkJdSFPHnkQCfHUneyX
s5yXwfnCV8ncSnTM+J5+abb4H0UGqZCF+la1z1bgHCnkt+fsGz+6deern5s3yYrcTseQgrlbHASc
awp+g3jAH9LXWIqPKwvJshe/p0IHlDO5VLFDPmDUwVOIEnzryrxRE1QCRcGxEYoVOHU+ReKcDoK1
zux+LwUdYR2P1C4fSHhAfmy15Cyoi/JOQ2VXgaoMTsX47YSoSZzkT6u1GDTcd5UIad2YfPdOujyh
I2NvPprCCNdeuhhK8rqx4O6Uvl7d8aizr5OAd4pMB6buwTn8mSephAlD+BrSSZO5XgIyq1zkgLa+
ZJgpqLHOAwcH5EFTTmZjokRC3MO3/AGxOso42EUe5butlgpLRpFSNe3QsyBQVlVWlX34fx7OUyJ/
j0Zm94/3YD393em2zJERa4+eej3HxkRp+bYi5CFc075hUS4vBrOkhz1+XQAaS/qJceVtNFPC+kcS
bjFvoQm1QtckH8Qtfp0ASg4y7La3H1SXAYDbKhkigbDCwenDmBidaXE0lghkMdiKfBmSFRWO7jTp
SunyRZbldRk9jc4DKPoK4BktNAvdaJ7eScs3lPLh+fud1f1OyvKFHCGplXU6eRSYDdIAgzopSq1W
NU8E+nf8JUp/VnTcOiS0QMBlp9g6MVNUn+XWdD0+f4vxdzAqOA8xmRiv9uGu21rsU+KDZ3OhkO73
Kh981Ivh8clcYGgJr4WDGzusLTVSW0Gdh6lPRPRW83px0rptMX0RlZC5GQFjZMjM2j8xswYn3M7r
lQZ2A6R2D0FDy83mA5G8iRqaqYrW9cNPF9LTR+tdI0qSjE9Lmu+yyGwztCOrLzrHgD/zCPBUUxJ2
EqVcMiKzSogL6OwqthZNPMqFWUchEEJXLlSmmabG2nJqkiHmr15z8H5/e5iHuI7vPwez95ghN38e
Fo5cmpLKi6pkA4pF4kFOdSebU1ptK5MTEw1srhtXoUCcaEhJ7LIe+NJ5EJxdj8tIGE4LWcp4zu5C
awXyZKOvUDAVXsc8LaOHyziNc/XM1g/pInghye/y+ZKcarZupTaBYhE/a7k3Rf3ndDXxek61ZfqI
wk3Kdj2bAsnF292tqvGByOlqOX/7l17tkXrApVnImOs4SQAMr7racktDmXKSGkhfbgkK3Ycvw5Td
8IR5LXMzLKeqSxwiTdqYMxb7tReCSF27mQRLEi/48P0xa7ptlky3tfMwOUYf4Q0P8c8PhO97WkMh
7eF/9PQi7Xmc+e7LznmrhXWUw3AuOROjsYUvZY9UChbHxYqIZq/KkrhFx+iLmdvqDYbeD6SsBUnJ
NSrToi7yMxweJSAHhwYGC2DnnsXaWJjeg4ySRi8K6hNsIV+wnVb5WhPIARsMOwYpF1lQeMO/MPDK
C9Dm9caAOTrB/GG2mbfQa+WfmVSQsogKqwGE+xB/gBQSjlv68DfcOdV8bvbev7S4RXZ3N1xM34xR
CNiQs/0+YTMsi29Py+Ht9Gb9D851COxZ136xeM9D1y/esmj5hlzkG6pNeD6VZcMUwmz2QnZ+cK0o
S9lxwJm7UJr4BdqCm8L+7e3SzhtR45DaNz7e/luDbUU9iVpy/qVomnJNsAxDS9dEbMHaL41unGaC
KZxqPP6HBnhXI95KNJuQjN0J99EV6f/edPjWB2HwmSse+T3T3TGXsy/Ub5SLPDYpup1bPhjZpYL9
QVd58L57Xopo1idxnCPjynaoUIbYLfGVVBZFKTBo8F/XY54mXbe0P3/qYXO9ifAsP/2SwurUdANs
dVkZ0/lXAL8p1DAAPIv0PDHbU4nEW8z7qYlBwSKI7LliRyCEqVFk7M/QrPxvEfqlhUyz2ynSF6Ma
xdk+C3DbU4tEx39Vwp/oEg5Tha8iZVaeFeqUryWZh1RRS+SD4wKOykKqp39eAt8GjwzUG79vBciz
lnE9Q/fjORg3TK8k+OT9ypHZhedxim79rR78ZCMmRdXDox9LLRn3g2t8gGxAETK1R5PabPxhEyOV
mVtHgs7VrWVGqdR+Bdh2QV8ONi5k8wvNIIN5tC7R06XIhr+ElhhW+3Rqnh4JE4FTxw6jvZVAX8A+
stZrgSAUs1wyexFxHcZ61/KcAddHMD1FANxw6hnLF9Xrk71SJ871SwZKDKrhMaS+7hgaKOMmrhhd
8Mj9tUI7i+seu8vgnSJ6Zm8042TcvDVydllXaGq0Jdoresec24yyVw9zhKL5vun+0j5DfiP0sBYI
LrQ8unErLFJcYs47ia1EV9qULL3DVUaENTekKv+Qr6n3fKbHcXBgs58NBFleEVjizajGD0bd+gFZ
jgqy8LGSnJmeqh6hfY3khWcGXiH8ogyxf7IN/MVw3nWF0TWCHM3k9A2nrVeE9wJM+RZRvATsC8wo
tsH8LHjLQLmi2g49Br2eqTF4yQNrHvjfgDvmAOpvXY9E31DdQNLjExVnkkathjksdQgCQY1KH8f5
beaVdzmBiWykjMSA61y3LFPx/lX007PMKYNuIUWyumnvfdCT5ahrHph+CKTfBQrMr8qXlHS/Yaaq
b22VsdKGb/k+xOz1D32vZAnUbWdKJ2PYcNVQ5zATShTuBhmt79gUZh2g6JkEqe3tpfJHv8V4/ev5
Kp6UkQc5uG5TqVG/Lsf1LtBm/HH9fqXZBBwM6WsAbRywH3VGaCPZgwLVR1MuvKcDQfhfVG2OlTUS
bKbMrO1cGAgVCq2wi/JntJWlAsETihcJodOVjXWCJ0QAxkNXvuY7lJ+3FbldPWA9CospdJgb/SBg
ILxek73ZWqqk98tFchgtcpxOmTw9v165rZgwIIG/EmiChv+pVmva0edG+rsx0sKfJjYXnrBJLQzV
mKq2GpkAgIw3X6naovyMfNgWfYzYIOGWgYzRhgZHvAD7pepw0DyceCfelTSN6nfHwr4DQ2sJqD3r
pDjuAqHDCnibqGS7gnKBvtuoOKbwFbBZXRQ+pMU8qwcHMVaE2Vbll4m7v6EvrARgPTkkhts6irg7
wdzcmfi27SS3lgo9tdeOtfuk3zzKv/T/oS6+gdt6Up4D3H7WN4Tz9+YpgGKWnHABkoxbAYsj/5YV
irLzTGVBYgp7XkZAt7IMPsMZ6TnqzYfBEmKdRC8uo0Af9JZYHXWYac0qQ/Y/9uYDfUpacJnLjZBJ
AtoKiKRFz8uQZSSstS2dSzCFRi1x6AiecJiuQP0AfS04PG+oQzXkVaoGezzufi2f7PNuH9N8vNll
PdJoBRVWCGCq4bCiEkfN+AezZp4RYNkXJTjA2lRwTIJM7iVy2Q2OcfnHRVPOKxhCDhaRpVJhiKf3
j1/okoV6qxa8KJ/fwN+DHue5xSio7ygkIXzavBt30T73LAIGjLOqrXk4UZQ6WuaTdMnf/gasvrYS
G1MXcdUBruNh5lhw+AALjJCg+oixU7N70n+fxvVRIxvJnjcTdGOoz69rHqrvV0HGiWIzHbpfqFxG
y+2RR4FsGCrTPcvYeswY69WC+VsNHHZTCq2Zhz/AiCwblGECfAovWQ5BlYaQw01ch520CrkTMWDz
oGjKSZh6AJ+J68D3CWN6D8NtstOnzCshZg5QHGrFK5DOj26xnA9CvoVgDadJgeP9GlYIoq7B9g2w
RYPfk+l50Lg0uONgh85u0qWPaivNgSmvnq+B91QrjO4g4YCbz7xmG/2NmxWbQj44c7lDMkEkjeyo
iXR3fLbYY/6rlKmGuxHNJXh+2wkK/u5h66bmD0omFn4tXc81SxP2d0gcuPkuWP5DA2UweO0RMWny
h2rjRQPdrzj4wTUwBHx+IqEnv95NoEjSGlEmRlhgSpVniE60SYGbINLFDRQvM6RLO0nr0KwAPBZm
8gLLGOCVfLNpBjzZGP0mR5kPGg8vbJhFumUansQ3JJIpY81AyRUKJkBRTwsvCnH6eRNUNF0Lc9xQ
+R2j010doEJbfa61J/+QSrIhy/CeX59uhE2paz9zQ2JThOnu+xVaGhLHc7qXUrhT3vQrx7Rdwjck
3fhTMpODffWlqpHv651tosO8honUu3j7K0MrtHoU35m4Oiw6zate7mEskNqbeGWjRSEd1GHVUYcK
JuWEE6i0dGlHVWGEfr+yEjnwvYPvOVV31hTY5Gz4UTaxldj8zm1xUYaihY8oN3CBujQnpwHJzfyJ
wfey3xfdKm4c9tLVxoaAXE/Uih1fVIpwOweIXQW0HKXapg+BTdu2a7Y3qxpcaGrRYoXbgurLNmzA
YVczmq5sMUqiahoOr8+MZjPnOcKIzrkbUBYXPXs3kPkbRbro/4iD65qtVXmzCneGsVI7I2mRP5Pe
9nfY8qH4Jbnqewm8UYCP0o7+Iiqxj6aatQMl6MopY77n9jQ40/Dxh+VROAU0miptYpy8RbfpVxm3
qPwb/xtu0Jeo3FSoKkNZRRcOcEn1F4Py8VpeI0HBpK1qjEsNmyKgPutbvCZAgrt3x4lif4QMfHi2
FxlT+RB8+9oM/UXpEVdPpwzrPdyXL7COnTENMfAYx8yA25hFaQ7IaGNVxeAaXqZogQ6cXUQznOro
2z/kg9nKuMHFN9pzMjUZuVBhhABAqpxRk1SAkRouqvdLdvbHdlBk+N9EbzLiG03lxRZ+gnRlejLr
bNwrM0ttCAdCVWV1ihWPrcYw1UyCFp7GzcKl3bc4tOu5n7g2FZrLnYJZx1FE3avN0ncb1rvB4EK8
L68h10ZXYIEiJWyqJvVQT6ZleVARZ8W/O+tzbYFokTsOqwFpTwEHyg4ttVOnnaurAGX3r5N8Wo9S
ZEWKy9o7FwtDyawmgo9a9ru/1bmfXyqR52v5ytw4h1LfOvZ4dmfibIhX78odGdakBb1KYqmI7Okd
4pRkra01C4E0kLXVFGXA/kQMrdIWlnrTFpAjTltvv5ZxT4qWnUcCKg+/xahUMfLxl0CK7uprSx+A
lMYj/Ue/rXI4vGN04U3pYP2J66GwirsDDJ/cukTdoPUIEREZ9+03vX9VoGd5ZJZ5kBrTJsDqMLMr
OtFDAR0ht4oQ4HgIbnQAi8gbq5qNJTsOhErpIT5+eIJc/Lck/iHw5faMYOVMyh4hGU/J9VRbRChF
wOwtqr9+qEhorISCrzCwlPLKnzMSsApRxofOoPPx/c7q7TzEmdl4/LBBkws0NzDWX4W/E1LXtd15
eFdAKaIbicxsxu3pKpit2htXBnN9U8YgDWaYicI2b+PAks7lK+x8qLktWqVkhQ4nOiKeW9XKijei
AJSbQ3/DXq2G6nyL2tBjbzMJTaWlplsesl0gpMoNs2xPolQ3XZ+yqWzqyX1agOhO4VkMJdl+zRFE
oNV/xQdBIDFAbTyq4FiTwecQ7ufc0PuWK0GW5PgkLC11/vVVXB0Hmj9ALG7FvZIUKn1b5QlB4mtH
YqDf2A7Nc+9fPCYzb36iDP+CF3oSZCskoYG4rjpM2mX+pT7AQEhagW/PZzzkamSnExNnphE5brmM
ATPli8mXKw6vPGYgsgZPVnICsnWS76NcvHHi8fyoF8A5op+44QJ95eSf453XNyWb6IZs/qwWaKsE
8td9tDrVMGAFotLjBwrOoV+NAWw2tCFfgTMOvm/OcsM/XlYmx00rmR4jSqcBzuiEouMxvHadSxWt
uOhak1KxGN6+6C3Y5qUvZlsUIdu+AosggEBb3Fse8ZTactQdjYkJl2+/pmp2LtEH/5n3rIhjbMxy
563a4vPwJ+5uywn4s0bOLrOpX+p5WooywXfc/A0UQNrff1SCq1qxmLUBOL2Qfd2LS9DsIEb8bln2
dmtm2spP+RfeBaXXy+Dh1cIVrdcvX3MppA0Je/1eBGr2gxez6gMYQoYQqk3CSmJcwKk12RZgfYTn
pHOaVJNQ9TwS5l6LXZHoUWIY1j4vNFLWa9HZYh8vi/rde/lXAGQcRi7yvAVbfuBfRir3LjL4LcIx
uoEPLYawEKlqaUyGAOBmum+mSWeLG1/4wI2J4gMONSWM+kpUy14VyYQ0ivbEr9w4CBlU8R2vsKYJ
84G/CP1Ra1MPQfVpjLSFr+0MB9uatj9lehbyLIqpykv2EOoW6uBQFD7qJPCV90BPogZ5jNaqF6r5
G++rTsLGG4BwLv/dZ5ehiT72pWJJaaZMx4FexdS1sxssYwHu5fzaEVwddhQ+PIGoYBAmaLoESVp+
Q4IdHiLJEk0TUXrMdGdT7Htxsjsm4svMr4XlLomNIu1s21BrSc3ArcICf2TFyN+4KP3WK7Mv2KDU
52sGhTgnatA3fGymDe9oouDXODl1QC4Jl2kG/dIVyKaNYUT6SzwN+1asglYTtUYILKDnNNC/THLF
BeQmKo3JpmwNvKJVDoA1exMg13GkNAkZEqIARqRtUQCwsERsiM+cmjo02X84Qeb8IKDOAeE6VW3R
z2EvkUCp7pIHvkeukgRFB0M308pJIrWCPeOnZmH1QlFlQmv19jBsTvovxxGLDDbWCC5RhOpHrWVs
L4Lnc87LOXrktxyBOreb9uInuozRBOEA5ToMXngdpEYuI5OkxruudPwPv/VRwBZNTHMPVCm+I0Sk
LNCNcYCRTBXu89G15oBkNNbdevLWTyFE2kVYTp12zkpXyToPjQs+IrIbF5xvUAxRFMeuXGXYsn26
qlMGDI6nQKP9RJXsXHztgYr8IszLjrqzi3GPOm1fzeI7L2ZJ/kWThuVjrKgfiIutSudB5TGrP5eq
hN+9xLx8wvfALacvnW8DZYtiKDxI5gPPtzX0mjSNF77+huBvMHTqImpRNOpNthjTR9UYtf6jgvJR
UG+1KNruPGPEVF4MQpKFsFbWuTJ0zyA4rltygcVAWxNAY3FWpYhr2+1vifNL4s2rBSsQaPxuH87A
hBoV7yKA5NrbIyq/cv1bk21i+0YDOogBs1oae62dZrVKCtLXY3rRtxUN+kbUp5LlvEcCPP5gJB7s
MoSe0idmiZYBp60zcxUTMNvs3C5LAgq+M1Xpjbh+MDNR9htowaAQox7zLE55DO4UwEyOX6FY+Y60
jqryk/enHuwl8qZ1QSrk1SLnahslkXzYkZW0CMKFqg6VqxdIcICcaQtQ5baAfOqf4EkhqRIUldmF
5fHeKpsXuUBDGpKu9ew/513CDdjZDK8RMiboDc8+aA2KLaWkDcDkiLy09CRBWVuYr1D6HYoI2y0g
nbTPaQCdNSjkihHv7p6WlpyxugjdUpIS29OkrSP+EZeArVgNtUMwPTDkmhPyqCesekXlOmcErbdi
zj21hyR7seGyCrupuZyhOX3oLrSDr/X/vduxNrZ+7LoDIM+5tXxoblu9N1dgBvGhAwb84p1ODUHp
0KN0Kwomb8IKtfwUx6tdhoZZV3OdPwswcodtjIl2xVzdl/aXFdLXImQivtRejHJscEv14L6mUbnu
PfKprZS7FqqRdbwLGAYX7N0ZWu2oo8zePmhb7i66hrri/6Bt/8bojbnxnh1Zu4Lcuq5nyV6U+DqU
6HNpsRDcxiEH/79OAxONYnv3BMMc9+Ok0GfhP78AVVRNkNK7PSUwvMNEAwJvvrjCrmR9TCOh2xiq
h54tqV80tZRYkGVPBtipTH/0DAliRHlKCeysEanY1envSqMgoO2Z7IFi1H+p6ukZFGvNCsUIuzbO
D6+LTIgnBP0sRWp7EF6iFQx6tcJTNz3bbL+bpLYelUVai+Gf+VrlHl4Wg6g5toI3snFMKGLfqaAR
XnZVq6L8mygYrTipEdRKC50nUbXTrnt382PBJN95xhIw+4c9gkApNSF7MeHD+MxbEnjJDw/ohChK
JrvOWSqSEaEZPTPoxI+7QaElZcEwB5/EA7UjgSIK48iG2+NRylk/MTBX4IDtDH6TK0Kz8W765X/d
lB0x9R8dz86oPMywnMGuqOqwBrWE8CxzuSpaFWTFVmHMyu3zFKxa5QQ5jfzy0Zw7yoQYpbAf66Pa
c1GD0fb36Q1Njk3TbTPRZdSWpTMFU1axmx2dX7aqvhb6ldzCUNoALOwVe9P9WB5qxF8FQkonw74o
NkCyRUwyukeh05gv4W1Q7gApPPhYBgitVATDnPDSf1PQJDTKCo7oZbBdnhZl/kD9XVmRnLMmtXp3
aNIJvE2wYDmRW2zccHDBY4kMGjqPzUgJuD9BIXmVpUgSSmdaeWUEnYS8YgEcAQIIWO+uvjgKLyHH
G5GiU1HbPZjHLu73T0G22cwtxxxrA4FF45XK1zWy7io/vqQJ2V++hcdRR+qw5nMOAMBbhBggMRAh
oZwfZtZ53voeMB9MHn9XSG1ledjW8zOdq/Yzlbx8++MnOn8xDHJ3zF5eaFO9e8znAavjqIl5BQzq
9BCtdNhbgEuq8ivkxS7VIpNFmjVowIOz5uQO2Rmtt6HjPstitdVhID7cOazJjeGPrB1McPxrN6Zt
WDYpThMe0GCqmzOIyTPubrs0Gv1iuDVvCtZeY7Fyq657WU339nHIBm9K/KNeKNk9eIZEwnDMVd0Z
6MTzUyZO+gTmVTO6vKDw8URql045ESWRD9uIFNy1WKPJyOgkDcLQKetcYakGYOodloRpZhPn90Ct
TIivHjmeBW1rYF220HDx2JfLraAtjlrX24g3En95aMyYCJdWFGAO54TDGI4s5e8X1r0+HNsGvCgx
YIuJumWMhcW6MqBzMJtcQWzACID83vGBnM39+3XrhPdFyNHh40xp1bp9wSDjqBB3yyD2h21DjZ6X
vhDQc7Cb4CVEtLnFJJsvpTtW+N9jCC2qO80wxaDNfccWPiLsIvy6ZgmbRh9Ey+5DApbtqY7xklPg
VzOATk/07Snr/7A+wAo0K3Ek8110bWdKQ2fvdhxCfB927bSLRGvbMF1cIinikNnO0pT+RM3745x/
aDKHn6GXlbAaugGLvoHWZvTALpXLg+JMm58BQtidao6PelYQyS/Bji5HUW68phUsDLt1lWFkm8py
J+6Yv5IB/x6tqw+ZmUov0tgq7qWLAnNRVJys881Iy8AMYZ7cFQtvgAvL5NlXEUkCL7HH+DX0U7i3
eOAzAK6mxyWvwo3s2a1CHJOKQn4pgWLj0m6ZjOF/xVWsTo3CQ1hB65YN0rLX3aI1sC+n4S22z4YI
8FH5vg0B83LXODqfF6c3felpVmGB8H53VXOecEUltBH48FqlWuHqOH2um1bJscDb88fpdiJ17KAA
VgfK6bAVSxpZ4S363I8X7vD+umhIafqbQW0kzHRfLn1PtUAFGPSn0agevTmQ8J2PZwryfo1G5Vmh
K6HZFPLUAlrVustBoLu5cbm1W/FZbaOCKNLcngO6U+GgkXmBQZvnoxanmq5tWrvdFuCxzx+KEplk
w92aYmABUm9Vy30C/btTDLNRTM10XVF1VOffEB89yNNv6idDq9bed0rhyGOz6wVbe4VD8QGnrF0i
fOqta/K+fgydHggTnN1K2J3rt6OfsNakn3W8T1EXL9XdcbrNzmaTlSQD8zGbvMF+hTdzSPDAa7e7
DhZoCOpS3OpAtV8krCCIlQk1O2Y/WQea0AKaDmlJiwZ44ZEuO7LWXT1vDkMHdoFaqx2HVWk1cq5H
FGqRsvY0HL80XgX3N5Vg9SKhaHT6LrxJc0qfNy+6JpQ4ZEGWVyMG3RJtnpiuPE2qsyORlZth5jfo
uXtbSyD1QCiAOZPyFIlvDLOeT1FINEMoWU2eCcEN1Tb5jIALYERbrA9VJKwfh5yb0su2A53hQ6cy
f7tygtjoD2YRQ+aBvwnTg+0K26ZaiABPDQnlXnGLjiupfFsZXMWz+/NWuaM7wOPvxyB8U9WtMb9N
yJdafVrigpsNeRel2mD0b9XUQEg7jr7Kh6iE3Oju2e4fH1nZKJVOLBN1wPvw7RbEhvU4ZTeJYxwe
m9xIJTQiYfICLXiykmNJbmvHj7dqEbmQ5iOr4H6UpOHFQRdxStKwcrKw4mxChN3Za8Uhp69UlaAt
UCv5lyXhFxLXkG6vnHv81OqXrVEmOWowHZQ24EbD0q0k2gM2pbocEYT9PcakMFTj/lUJGsRLoA5f
GtLaUQMM+uCKKEiIaOJXFtUTaoO1UFBj5/BW5miMTzxKIOMv01/uE40fgiV+P0iwny8vdxc7SDyK
lYnFv6nc3xHWUGtQ4Q6Wgudhcfphjr/vvH7oj7VPFLuYEda9aUq+Y1hZNn8Q6+s0XLe050BnNrYp
ngd53hFXXg3p4JAOYglqDQl0Y84jrebqOS9BE4rAwukKTRmMAYIkJh1pZi1Zek4RtMqNaghFaRBU
I442N/G1A00pBDXRv0SQouHNzJ8szVcwPoJ2ZfuNMAMclq2t+L3uhEo3ZxUiU32AgD3r+3UUsyEs
LfQj3O3XhV64AqsWi5kmLYnrRFYuoSJ5h+myHqrnwFLF6K+aQG4HZ4oAjFnGWJjd1zCPfP8IjgXk
u6ODlSFiseHDXkVm8Zr/QBXO600Q7FUarJrT4fqAvSfsmulrxfpsP/EmVnMom0wkmqgPeb95QTFo
hFrWw5sVaNPY9kTwgDSemtRoutgOOWd+gSuGfAj9N0SH7EgIv71x8sHkAO4qoSgppbfH9+wpvpI3
PHXmWDAv84lkuYlRL2m+/NeVhWPzFcBusVeX38Bq+ZbWvUUyoTXSFtzUpMgz0yF2m+w9PbxMKZbE
wdT1fhcud7luP9XsSnewC4YU61NkVNSusz/KQm6KJWWbSsS6JLtuvbil4YFAwC+iiep0lWKYfxZg
bz6+CtXNKLfYH+5m3lFYOXcuhqgBxEQ28EdHtP4FogGZn0LLL/plrRoOdpbrkjCiqJeWfRVf4S9k
AKfnzT1g8f5vZzeX8dXcdGcsKVxXPtiAHqrTGLxr2FSwVrxWbIRNKsnyi12b6o45EXwxjt4jp5M8
aTXxqvYi6c1FuQwN10IP9it0v9iEQQC7TQz5ZPnmEbGfTpQQDQlqPPkuyok/LIhej7hW2rFKjbc4
SfGjY/S/6KO7gsI/FEIPBFTi5TT9fBeKo31JQLlffIOkIVvrzkb1qk4O/zRRl6RqhChDZtXBz9yN
0iq6sA+qtljixgCzQcGAI4TotcuBUgX5ZrnvKAQdE8wKXt+4vhe+oAkkE+6gQKym9rQiscKiwnOG
eTrDjM1hsXN5W5tSA4+8gwDh0R/309FfqqOaXTQ83C5Zhfap7cbT3Bp3sWSVpkG9FvLsYfVU3Qd0
2EkGEThStqB/tWkeKNbeHU1bKcuBkcFQ3qAdXjQi32+ujL6+B3Y/oCz0RrYgcEB8Ey1Ne2ZwQj69
4u2f82O+13KfB0TPlVDfDDtWbHZRbVhPCNItgQ9Udj4sfdfOX34VzDQW3ZgVuTnR/hn+pbew3VOW
4JwRy4o3GAXQUfAmJLJ1L+IlIaaCkgWTuGhgzNsyeldNwMBIu8wYWrbhZ4xbSjOkdsSsQzOWAzNG
/zKsOWfF0ft5LVdNFbiR971fc7jB+PoPPSoTxldTRq7x9Ag3zJUTVBa046qlvrF7p8ADq6L0V5r5
EyV/t+HupstUILokxyuNh1HiEC0i0+6CzUEyJkvtR6YMxedcEc1zwnEoQ6658qa0zzeoe3Aa7h2h
Ab3fuiTT0B/eTv5xJjMiqFT7IBVggK0Ckec8g1vF+QR5idc/cpuQ75aPumt/gqHpdFg/bqcH0DBl
f8szqjeTomJbg8VzoFF3TsUYiwxKqnY+ojIi1ROuXa14l5gRjzilcF9Tw1T35AL4JQCU74/MTMfe
9e6U9DIsl+cJEd1qe4/mR3XR0oxuUtKrAwZGO84VuoFxOK8eXXuJN77cPR+0ALmtJZT3MlN/SLe2
wOr9Vc8AX34/jumzemU/Of8GxzslVR2SkEq2NSJT+KbALkjNtVBNE3hIiZt2InyZWugL43YYE1ji
QShl7Mqa8IcgyaEREFVQPvRFFxVnYMOUajmO5QTpNeGBtPEluPGg3VjxdoXR7KkLCbVHcP9M5fDt
l1HwZe/lwpTc2zS4O4wFv54OWqmlwZiygLMehGLJoHnKFo4zW3yo/IMj92ZEMLRp44hgLvVKNze5
UDgLFIF8CurJGzE989SDUyTnYkmFPPcLN+kUws8VSYF/c4pACxj1wy2W3YjQgHko5xhv7I83D8e+
cfcFyb5ZvfJ4IeLQmVlLgohCRaUPnh2N/XIpoUlpaVarFvI+0GhW3gOlBbhHEaK9S8/ZvLJTaHjV
zBF4lYlN3kHNDN9YjUVOV9e5HRbv5zDoMatVXnAkw333P3JyQoLfBdB0RwalAe1faJaKJQfY5M4Z
s//o4P2+iOdUqF0cnlGjGtildPadRqPaG4a+eBPJSVl2zJYoMf+MtQIdXUQXpY//zDQDNHFXIghL
+wYBfCYYh2lE6/kZKbBQlbxO4NHZOJFej/ZimYgeKlOZJiPs26UDevuknCWXfIczW08dhHbLizci
BfT0UgSLuurekpMgW+6kR72wIS+E/9+lD/s+cjRYONcjEmu1/vBYQbVoB+glT06A5g33PhsBbXy7
kA16HmzMayYaJTiWaOizw9QnFuCqaier0Wyn2CChA2W9MUpPg3Vx4YR3uaP5VyvyDij6ZXJGi0+b
xkOpekN37U9t+zp7rE3DF/pfdjT3AHgw1hjPvLXcSD2n3I7UnCKAh2ZPxLsN/1/76Y1vwebzRvaI
Rc+AWN/HjUbyAqfERZsVG1+yCTVmcje3bQ6kW7VSqi5faJTXxVhxlrjGc2159d15/axw6QkM3ZPT
Y7m3xk485cDuhrVPb9ovVzGktf+6Ch4AsweFVde8FZegnppkUYHz1zOg+uTwqvwZ/u2pqr75zOKd
H7ikdzdsQvcb18L3tVkJtSjSSvf0NHFsleJ6Y+02lJdkYmLDY4gSxhlDJEBnswjFamd3K5u+zvXM
gDpC/UuFgBiE6BqNlsRn20ADPpF67QU3i04C+nAb08maZqzMGOM5B2c+xpqHkXEX+zmtOvXgQrnk
hNeXu5fvlaQhmwHNOXo2NpcexUq2ftNl64SD+0aOrvAIuKC4Pj8OQumhu1Kk2LD9ySUotW+9BWRP
SH/VzBs8zmft34Jq+6eGopKINLu9fQFyozy/wiSYMD9snUhrYohqL0MHiDrAVvMSIx7gP3uc8TKa
SlMUDw0AqGwEA68IVP8InKwrlLjlI4hZ07DHI+ktm02c0yDJCXb4w/JEFeU6xQEaU2hOfKSs9gRS
iKRR2Y8rzCGmHUxUv99lUMjZsTKS3QYuR20aSlK0Oa7Wifgj5CQz/zaWaynN4y/vp1G9Pz0PgMsY
KA50dsFnbCr28PeNtZrxCFfM4E29uKVeTaBRe3jJ5qwLarMzG3JxIPhrH4Bc9wWG7qtOubF7knze
JxGzpaXC7/0MeZAo97FnMJ3t7Ei79T43rP6rLY3he3Apn3Dhclb2cw+DwRywoTCrkWpjjf8aEEN4
Uc4mKk1829s9Vc/1IXYLeME0sCAA1pCoOzU3IIBdXKicDC1AKLk0AH0a3sCNCF+Ivzga3E42wrC4
Ek/5tZmAHYzt8ovB/9C8Elh6c+ntoM7yFyr7eRDgiW6UPSvQAgfdDdnKonHO9ugRAXyLjEF0lB+M
r7MCz6CsiSWFC+soaaTLZB1amW3kFkKyjzjR1rQ3qbLp4V5PyxgmGE9TDxNhsnJUUdLYUrccHRzy
nnpDBqwit6HtR1FOTsIXIvTJIeiMk3ZKWf5BWu0dNvcUbYT6fa3om1oc1RDqsg+1AFIQQO1pgEfU
GMroxyr90l+AEZA7hxGC1B7CWrvuxcaK9SfdrFLehks7G9yHissNdxAPpTarEFjtr4ZMzXKZcFPb
Fo10u0peOYbxM8zXGH3cdZFaSl9oSOY8vUFYiEpm2OUs+CPfn65dU3TAdgnSfaDr1lLbB3sVfIyx
3f2KIF6JlJiAjRqPK94uUYcO/6naNO9PbByDh30TWXPFG5pR2/6DC3eR7GJDO8XmazZ8nBmfB7xL
E6FgO4lOcaTQkWYH/c5EgFs82bFVNhwp3vQbg7144cPQwDJsyg78sxN7RtGmIPtoEcyPfKAdb9Xj
ImnPVir42dlhwKqtsmAa+E4mGKtBUtVuT/SR45egl/6ZyO6MAYJiMVCFSgTF3bNfvH5mNaP6wR4H
7EZikR/PUniqrNTAWKwOhzA1strGTvD7HogX76Dgd0KqxC39i1EYCyETirOqumQ0QesFrVjcq3VJ
NKPpP6koXos+xFYlnSo+DpA/e4QI+TaOOityn5NuHF2+OZGjiGQQ4kTHskZkujz4ZBq+uYRJ/QJe
MPYydC+tMplSlJ71rFX6d6NntbJboI2k/1JGOE02gE0XMbsofEJj87sSuxLzInL9audNdIzpS4rw
H/h11IbpYyrEiKJI5z9oqYxT2ZVUvSkYN86YLSA+9KGlgzUsvCo+QAiQXEu5n6Nb6LSIajkthYJW
p0qv7OJnVB5gneQgG9S6sL4e3igkkCuLePHYGHmwmiYskOGHVzA8KiZSW+TQwwHlWLeVgc05lF+O
8qdKcGUVFN14kXs9x/xiFURDKjjsoNeA4e67lqOTob0BUrW+s/0ZMqf1WMfoXKA1SXIe9szr/4FN
J4GYZM3omHCx5wtz2Rh/Kv8HAlRIL7Tro1swlBfVPstY8JQWYcLatNWHnmj2zCIDKVPhjYAXRdc1
+dhUkreTf3bFaopXecKo28lBgRptGFxKwRW9Sia+/cKZe4sgVbZ9QKFnvTY864Indq5hxWl+0Hlw
3H688g6Yw2paXcr523Od2qooEfpspo5YQEzKynxQGr9sOjo714u996FSYSdYTnhtOM08nVkRRvtO
54OzvTcClvf9mF4+dReHn4ZeewUEJsrVRaVtdZWehmawRHbg7R0iFkE/8wSP3uMOEykiIwLsgjNS
NBayqko8NW1HXbJU15mr+zu4f0Up/JH67oVXqwYCQT3Ht9GdLen1NuVdOtg6Gar0slb6c/gwScP2
bdk7cx2ufcAQKc+/1bmRYT5pRr7bSoqvwLjzgucguBrgUoPTrkzi4hpbfPlikumUiHUral7W42gp
C+wSNX4wP2x2ra2lMjMtD4/8lvZHWcoQDZBFDtfeI3ePEHj/U1v+3A2GCvneHP185lj8IKo7XzKE
JYySGk4f4sTiu+hMcvObNsitBNVshcJHUDwOFhfkZz0EBmXMrcVQXNpPBRo0y+SKu3bq3l6Qr8HH
SzX9GNz+TT9HiQn51oRWNhU6x4+Ikx6WeQ8IJ6pL7kxS9bHiOQ2apt12z13Y4aDmfS4c7aq9pB4U
wfgDLxuGU78JATlNKqPUJnRMS72z50EV10qfkcuLxCYa4hTuXnxYGWxmCyz4KLLft/d2wrd6xHkd
pLFdbV7b6cz9F7RMDnydy8XV6PDSG05kEg9GPJmVJxAGSIVrr71rMMcNbl+rZcnET9Hg31GiiXK3
GLel7Hjjc7DOh/C8Jty3SGqLrCxikpOylyFdSJ+z84P3NikneHa0E7UzD3PO4UssejIAyTTRnDGf
OkZu+zyIPLdrI3W7jjy2iLsZNYKedbUK90UDMOPnUhAAE74Yn7CoZ8sY1+kRn704R2h0SKlN1v38
/bQgjIuDBSG7CnShqzbTCbspxSuE1W69SRGo6DmjP78DDyfyxnopE0fwb9D7ASppR4Km+5vBOPdA
9DjAa2ymFpS4Fba1FzZIfCBDRUfkLnwmDbEKP74fpn16L2mZx3ke25qr09mQfzHeoy3ieskOu6W2
XnDwsHa4W5Ussxy22TX4rbxYQBi0C8KV9P4VqJcvv88wZV7o6TjCtDsfjOzEKanG9vV7Aaca7lal
mkHEiUMSHvgVqV2NwP+sNVZHYKEqzPL3g9dqPuMTkyAkympkfAXtO8pdbY/5Qaggz3R07w7EFPpZ
qUcMh+6jM/j2pERRcWfRuydEfNumrdwWUmYFpoVLrkuVxXDEEb4C8hztINE3+v3zDviM7gMVIKXB
x3u46yCIiHDS6k9YeFCoAbEdkOD2k13Bmq+LMTAqT82kv10KkRUqkNzflcPesZYeYpC3Qis4UPpC
fRpH1T9OkSs58QVEOjYrXZUBr+FWvt/ycUHRpG7FAKInI1SL+5xwasMa3baxplPYpyyd3c3k/7/i
GGM5Yl5oHf6RlPqVxBTlDkaDxHDIacL/9s7fwU/aPBxDs7dzA8DUfLfePWtAmgTFtv+7GoJyfKGa
QlGiIOoQ562wbC5nJQvYu2sMrwD2gMnhvBLzOcrEhiS4enCboDxeZD5TPR43SRAI7UFOUcpEjzTf
Zp3eD72DSGhWkjSdZsq/pb7LeeQC9PxEjXjTHr8Wo9IAwci0iQDAZDEasV2xt6YwnSedTbCHBARS
YfLpGMSgqKQlCqdwdNUEkqBpeKIECJBymgQXVxRvI6Jkeog0lKo3fRZiitUJhfIXC4wcQZ7toKJL
yszcpWehrnEuZgzHh3EeKtyGZtjaSm/Dst3aMAAEOrfLGSKaclKVR/q+ptYvUYZNBUGImuEZs/22
j3m7cwUNeG+Jll1G6r35zwBGbFE4PhFWO4rxtQtVfbrLR7Wrj3tSrFKNxalB1qhb4HhvW5P4Bgn1
f677VycXJCko1+wLBCV41kA4fDYc4jd3AHuZFycvJLW53jrGB7KQElWCkD9CVQYGbtVJUgnDZK80
w63z6+R4uteIQ99dfRBT2TYm63K32hUFxP0UIV7cx8XYpc/xgpv6ylvhFT1vWi83L41wJLQ2z+Gp
xh57DZr+1cxjwATyl7lInK0Q18eQiwgngLrbSx6w5dzLYq3nwRiJTHdYa7c47DnOk97GowhljxRY
5iCzk1GawewkRoGjTx625rQHZvB1p0OXi+O0CPQfrE0pcLMsHeQ/bBpmA2WSITU5QgwUQYSVzySc
JKKLTrcYkCpBzQD+OTOkkddbfj5n795QmyGG2PcGPgptIiA+3yvkdcs1ntCCOS5/N8gPJQ2Tpy9n
wIOPFGKlc0HaWnG7wHcEUvsjX2kDWERAQ5sEG5spvbJUdTAGZaWqaQZnAN4QTpeBiAe9uexaboUQ
W+yXgmx53uJ9ifGMSkojsXFQM1q+LPeq/MPBbDABPGFfaXyqnC+H6cSNYS1+2JSCiVU4DY6IXoc7
lh4j2QAGfjc6KPg4IOwgYQzBG2jH+Skbup/kqXSZDIOAyNgLVEGGyd/gb+k1M1dgMSwoyM5UGFFA
3zHNlFakuQ+LefCsLB+IkC3RoN7B6vr62zp9GCI/zSpGfEcmsxBw6TW8lszLqIvUawEDsJK1UxMJ
2iKVnzkBZzepy+HfKmY0EXRYEF54IPZyqTYx9IX+DJGW43CgHiWfKM1e94FniaxaFzfFxDBoPAIk
avYNj9ODvegKQ3FnNlf4MMNq0GoelISzABdj3+gUt6bZIo0LNkTG5iAJdaDasiJx+eWFsXOPWLj7
LTCqYZM3wd9+ez2eC+TmH5fcPE7UM/guM9gzTEQPuo+W8wM+qNIqUkian5YDEBieMJMRqc4roW63
37Joa675tDCUMafoQkRr45WQIs92KfGyAZ6WBTEmuOvI/LNF+g0EYJJHI2V9HS77nfleknEduEi8
7clOsk/pJjwMU7Edg8yGXbfemULv8RDAAFAaWUhLTUkY1WdufjrAxCuQBi83KYjuak5yA8CUbQdO
0jlPE7HJbu3DaGcgOU7hlQgA2VM3IEw0CwL7X+o4ULRwBe7drpGUXYFpQLhmc4riyD8dwlaNh+kQ
4wtFs6jS/zcAkiTNAkO7Efm/f6Fu/k3+6j8bhEajeBalC37IO9m6jklKX0gtE65YPYTQilRb70ao
wIEjgeeA4kP+a6YUK/ETDb6uHMpdgF2qn0yMfgSaoMqozIl4obVB8m9dkXuy7u/lqXdqD6mgqGqO
v2jUQ7NNbYtAgxZ7nLQ6ECcix+cDeRVkgzsMSm8nHsBfzYNn8rKL9T2BT4krQVZXqkzYnZB5whC/
XCnQLYKbf5IuKaffN4dw5d//1nw3haovIyfLk1OCXUPIolNGDY+xKPoiVihC+/qSnTheUO6Pyo5c
TvAGXki5itSNdvx7ptxyuKKHDcn4bd6yLb4aYdoIaXL8/SGaN9RAjdBoXt1xjr+TWvmLJpN4m1c7
meIHLDMn8Vkvfj6U4Q4et5pVwgg9ZTizuh3Hugsbnvs8dOMw6KXg8BHY34avzoFm3woImLfQ+nYz
hdqy60mP8ngtl5Hnp+/iu8Eu5Y6+/GKCsYHm+cd08kZ8IaO2msO7h3f8fMhw5iHno6daoo3MYqhq
9Z7Ud5BJO4HlBGVsQIHppH7dlwlFnH4donFVH8muI4ELjjpFgjPzWSOImXKCGY4LqSrjzwcC+Me/
+pitty8NJZmCQDfEEVDu4JyBlaG34lrKOUYMyZvcWcbmBDEZyd9DVRp8b2X28v3FMI+w2iaIRLi0
2BhHNGZcPBpvn/KMrBzW4ftqKYZZkExstirUk6RZkayr7iGL9FazyvHvfpNRSfbnS1Im20Sm8Cb5
IP+z+JQhtLtizYCp97VQnK5F9x90ICt7+GMGc8q7b6xtJhYk5r4GUHzFgTVXqr0VAWTah6hRpxVr
BqXO6OX+RX3a91fBYEn+AesmEfhoZ2qheD1V42jIMnUguJokezEb3uwbvewiNUmueQdz4l49BwpF
FeVza+Da9AbvOELngLDVoB2w4Tz0FwjTwkl+7W8E4nCvpFHSo9h6aEqnC5Lu0Y2enzF1BTggjsdH
uZnnYUQTn2aTk1P57AAsPIbsTxcJaRH/A7owFW/GRW7C0nrzLqYRZnsdPNhANX/s+82MMIR+ZJA2
1eoFxi/o8Yt+QCb3Rq1f0JmlC1uJ2K8PnMOLqK24jgB2cu1b/9u3exP2Ml5GmPpzO/HYupv8UGKO
HKFr6b4gzH1k9XoOmrleeYQEfSVoBUUlU222Xx8mRtF56PoLuFBcBJaEXy1lqGVG0YlBdbhRS58E
aqwsDgD43xNk8cmDVYy/1ba6lwWvc/V2FggkwjnoW/Ukao7+aQoafHk+vrYQuWCXoKX7QLiKEF6i
vuEDxX0GzloJWxKTz/Mdt5get4UZnciGIpHwWYEV4ump2HI4qsn0RqZzUWFwLqhVk3+m/ifGk8Vx
1wcYXlZLrgX1Mw/WPWL1t5if5TlkEZUcdwG4/vAw/dx8yqeU3lpNG+jg4J5xemLK1OBvo0p4zus9
LRWJC1/S820BEFI2UHlp8CV0eqWXVK8fz0QDV8nLcyaMlF3sgV5JpFKU+xkZAZs96nac1Cp6i5Yo
EfpNXtV+ntu5oa3GcEDRJy0H91LKZ/HE4vfWWiHkdDhyyS2qkWgP3s+gVOAOgFIppoJREILt15BK
/PV30DZKtU1SUHlFklBn5Z5ciZxsks7mqjZXIi4zN2BGZetkQGtd4rRR1/BzV2BPj1urZyuspwdP
wfwJWZcwD+Y/yg+D+gwUFRCsZeswibpSpbN4t2ZZNzKMUd5BvehzA87j06KtVzWe0vg7JDH3+h5B
JJUILPrP6oS6pDlVTxeaCJpXwy4sDZRbM2ULOZthe5lfGAwsxmoAPwdng8NeH0l3o0ThQCubG3kx
oBayvCfOUS0DqcAqsTib2HfomboF0/8d1abaEAt5erH1qsmS0Ugagvcee5MN6k+c11xUMolX5H8B
8ChnZWexv/iS6il9T+Kc1fD7LBP+lr7rFEsC9zEfrMLpoJFzLjWSzqCSYvB/HrjTbG/+DRIBXaWP
lUEFDrR6WeyvOns7t+yeIzEIIegZTmbPluVdwuMlOFmXkK0kil/A/ma7sB9S6GmFnE2s4XDsWWCL
mnqb7qb1Hi+wXgdUflUA/qI3IoYJe4cQlr9JQtwtvgOvOVENeNMR8LmMO8cvAw5wjJCUl7ZlIJq1
1CElEPyJho6yhc8LIHprED+REMfOtqb6SBu9iX4EMEVdMdxg0QnICH8dNjBWDXIUAu+cfjEOmcJ4
OipFEBGWWJ+iNORKfm8c3RJsfsdNlYKQCAKLKl4d/ZMhgDjmgNLNMfzTBVW22oa8/UGPb4sP+DEd
nT8VYVEBjOlLR1/pJo1pPg+ltmQp0Oabd8He/2CIl2uZfQGWDGTEh7KMkmJkVnPnIIduMwTbZAUq
TZLUKXiIwdlwS+UNxtvhIxffqovRitpQvOL5I74QhTFR31e44r2f2KKAz/ZbFNm81QzxzAKLClpF
184b2O4kTHNDwI5BK/FLXTsE1PbX4+V83Aaw5iI47ttt2HmyteW0/vS+D2rXS4AXtL9wxL1J2OdP
m7vcZSNpZ/ymG+Kt0/jqWLgAPELua4sp69iE4wkEzAmEKvBorhr9nQwLs+byiUlErNW5MPVl646P
35MwxpqSqlpi9HpZdbmO56cKqiLifZWK+oXpUNrqTapjSpBU/nxb16IQerQTmfGG5Ju/qu1xNzca
v/ngNkzFyJFzY6/8Wrb8J6EE3cHC+TObPVsieMbjeARzaKjPLeaHEuDDU98rKo5Da+xZfnDJk573
4n1jCbu+pNz1Jn2v5j17CFbhqvX2mGC7ru733c+RB44Rh3JgeVtubZB8XeXjhjiCo/QxfI18kfcQ
+lG+6T8p1kQWlDSGNighKLlPaAO3KUDW8/9cPu6yW3UqvZQd8OrG+w6mFsX1sj1i4SI4faDCxWwj
KMlwhtHCmjgbRAYtlBzVVonKLt28SUq+/mA6/9fOtGhmkuNtTSu0FA94+3TTs50qGSKSbu1faUSf
mDfkL5+SL6LfWkZVsdQHXfNzOQZWKLXcPyPoztpZwz3DiTVdihlgfJcuAkSVh8GdPitZAAy5mnNi
GHysPnXOYvALDOI0Ie7IEHNMM58ORm5DAWoWxkim+d4hY42fXTpafRa+befYMKXrHawLhwYsTDlq
6G3ztokosJadmLHCtwJtA2iy9uOKse5GS+OtJeT0i4HAI0sMz0T0gzARUEcSAmG7WRphwONQCSo1
wyM8cP5iqt95oYCpicxFdYv/b9v0H0tgOSvJm5/TAQR4Rr7IJZZaKYS+0bDJNRhvy5GqtvTWLuI9
CQ2TTdwgTjE8zs+HzyNpos2ydKAkEK7cZE36YaBw3Ui0P3ucRW6cofE9s/32ItM/+q90TcR1CMNl
AMxNmpSQfXmIvDy2Ao32Vfnpg28zoPnoAb4zNCVttkSz2W1HqRzfz+M6DgPzuZB5/chH6tWJwCwk
xNOiHZdVSwFJgRicTdo3ZmEZO9zPY+zowWrLvj5QqJUp6egPaV1WPt4Jx1S0xMD5/R3snMqL5XWl
7px10duCBVpTNpZcBfP1ATiRyJIh9MUEo0qpkAVPwyfOVQR9Xc7lEAtigBN3SYf0mnkn+SVo3WYo
qSu/tlUXaM0pW/JEAb2LcyQ1Z2R/4lTF0tDHXc9PE/qow6BCweg+c3j52G/xotKFTD8niufGfKD5
pPFqG3kwPTdIYpJovWtzqcRVOhwKHt7cPnGq71a9Q3+smn33+L9wrdKrbcOKNdrT/TSZSxsKpMNC
ie0qUpPYQW/9ez7trcbBeJ6QuhgWCzerqyhmGBHe6jNMSYou295BbEZ56mrOUjQ7rOwV51KNVSd7
Tk7b8xZryJL6LcpHa2TozsVFoqnU7mHjlp6Mm87vhigtZmPFXYLhZDbGMrdRUQRQkJWy0lor8Mvc
4e+RaEYC8PJZxavIYN4VG8PUOwdlR61yyIk38Y4gLU/qdjXgyy0tu6tWJywzB2Wb47Hy80lvlolh
gPNUsRPpRl55ISmklhAAyPfr8cxoyBe5grsdLxCymyjEEBrYWhkK0i11Ap1lAtL/Vs5iChb7ZR5Y
gxFE0J8eUHXmdZ3QuVyEzMZirnbslKExHygsnVDHrQlFTPFicELv0EjbYd2FiEE7V6dVznG+5c2s
xjB29enlZGzZJJ+/qElSM3hiZiVieAo+yw7bcQvcNGOyF3+VUch7yj+HChu4Wwb0w5Thq7KU8wnT
ZcqjLE9+bUGgn4r0NAllxoGEm3Xy9eY8wHw3wmMLG3NSJUB3cNYvI+wTOZthc74H8iQjxjHW0I2u
lBo9jdTk+uTfAURCLB8YV8d7FLjivDRVdtNVNoFn0XGcYIif0DQ3KqDTspFQS/KH8zP4ZeEKRevJ
02ETjJLAd/H38aaA2/pqmQpOjxlKYVIyf7e1QBS6vrP+QK/GxbvLgIb1tt1bMhDhfc7lxM0OKtAG
debNS6QrGPGsoV1S4uDQ5afCdigqRPatvZiRPZs1w+u/QfT3ki1foR5G+6MvrWEvWz07frINBs/e
jGweYN6B7IWIKDvb1s+ycYMxxqWLxEZPJqsBTGEm04Xuf1IMjCJbrVQ5Rn46UZ7mvYM70tO8wH+K
meIAtsW75r9flV0t3qyTWTXWLC1EFLaXukNfASiTLhe3F8jeQFoFX2HEQP6PZl5Nf+gdSJnlcfA2
5cJFnKIJJ/SpphxgVdhbpdwTjqF8iD0jihRcWHjnqNq5vZFFU5ERSYKgXKnzsw0FRNk58t4gQSx1
rYyOGnwTmkb1kdbPxWT8uIUIHNvA4AnYOhLiMMi1+q2cukXeTE5dUbAIETFKZJh4Mq93qlUVqDs0
tp/Su4EqIN09d6XIOIgF9NS7lpzBy96nP+MjZWPpUYx8CiKf0LYvn9kuGFsjXJolQUWVfjGgc4g2
Bdgjpv74a4FXsmPihUav0g2Su/qE3uaqIUN8CYrqNrzjQuLOYJTj2iiOXXTTN5Smt3C+eGotorwn
yeyGqt1fSnyyJqbrKzvddPkEOiwj9y5f1v5eDdJORx3zOQ0FmyEz3Jhe6Pyh5lIY8U5oahG6Ssve
EzEKtko+D5Pn5O9CGXG7DzM9edd/04l/Rt5qAOTK//saNbUq/Ju0ZrPjznLoBXQKHn8t/UfjG/hU
wAb7r9J0PqnHYxVY+L7LUQOiyGMhO267KkG+IEM8qbPk20phjfk73pwfTY6eps7tnOzGAACWnGub
IUB7/XXSDHOqyvSrUVPaBWeEdcGDsnQjy//6c3tUF5u0VN/LCc5Xxi1a9XKQYuUo/gfXMgg4AZmw
Etj+pIlbMvBQI94VwdhkxD2L5UThMUXfHmQPb+uBRStqDypQYxIBeLgOEnbepwyYlNd0dj1r401K
RK7eMBLL8Yz0mOIBR04ZkO6RqncOA6MoSkAWw/66vcGMBWvY7Lw61dK0UwxXdt1VQc5d4pvsmKu9
GlQ4BHsKiMwOQGNAxEcSNl9fOLzRBLaciVSDgOK8Ebxhvvu6ZJwZwncWu4EQIlii9RlqMoPmJXfw
TNDeIBzJH+eknkLTvAnwEzr7dG5sYFnBinN5MlS/LDTlWjQ27tSz9a7EWf4o/84hAPI24FWpe5tF
Dr/EDIppDik7x9GnYP+geXteQkeUw4ttpFpHPLFVIs1WOGTWUDwUl2mvKAI5uCNol8ZaJNjY+4OD
GSvUW6QtRQIGWyDWhb4AIxWWYs6GxxxS2IcNpNaQbRTxZkTxaOiIGMt2u/6mr+erZgoXwp/arcNk
uP1k49ZcUrBDCY8+EFMhTB2ak+9RWVX9TD5O3/Vu+e44+kADvWqOLoEWVyIWSrZ65H8+QXOw40Rw
A4rYVg4XGFJPSCCOWBKeHp9ncF/jh5oG5vJfXnTBwX1M/8mSZfEGV6XXCIkn3T844JnIi0wqEn6C
keD9HzJL6SDPgB3sNQt0FrKFNDd2Y5jXYn86UmqlR6c90Asb4aPagFuUwC+xzUGAXsxzxF7cAPe6
34hW92YEcGVEArDSRvgnwaXa6ugetFb+Q7ocylRmunHTjHp66CRFPI8pK40OSnPAJar7hbbg7Q6p
ju1bt0Btfobp89WA3lxQky7yl3JgpTT5ad23aEWcU5owO6I7APDHsLEoNt+DhgQ4xUOXx0+rakOk
1thBTnsDXF7qzh4iqRWFTSC3UTwXA4EJZ8TAAzUUM3SYxhyO3tZM3TGQn/fQOf1oDod7yH9rm1zD
glcFNEX4qb3xkNc6TUi6Tm3id1wzcvHFRQogL4dKnX1vp6w3M6xpudDHT1kNq8Cjo7I8Oz5SG+eU
v2Y8HJ9iCNkSCX2HSdAt++2S1yQsjtNx6exMyw1ypNgGdO1m50K2fRqh5aOAr2cMG4EmX0eT40Tf
O4oHQR4E6oju7zv3ZSS786W4YW3omUXluih0jMPW4587CSQ/snoytnTL2T47iCaVOvUoFenDVo2L
LNDPKWHR2rLnYgHJaH8y2/Mu3rWaCtYMcOwS8+iueDe9YY7/psJQes2gtNt7Gc/tuDRs0lMCSGW0
tmeC7CYc/x1SbTpTEE0ChG9eCssQKzJu9dFjwhbHVjEFwf5w/t91e6eMbhDbaztXzbzoufCTlPzk
6uywKRyavK2MYGPYfiVRhSdRHQ9SmX4UtU9JBaorEr96jtMtC7cgDL0nrZ/NxAVfK8qoQwdUulXx
TtYw3EOh1yA6MCm8eLJUrm+/sJZ5h62XgZKU0vcf4bh9cFvc5dVP9NrE7Sdo2yt4ys1rzLGrpYj3
fpFHiULJqI+p5aSJ0um4BOR0vj/SIdPmo5CRfNpGyUIAsZ0EClry7YeYhJtLN8y10hCfd87ioAhu
QW1oqxwutatNMlK8zRyVP+DOMkd4HhxCco0Fi+Z223Ui535yS5QoOf9GEBbJ5qpT5Ov6/BVF8riS
ETaxg8YjMIzZFPe31N0SFEpZKHluLNFpYsnaPmwsSm+8PzphFis3o0Pj+WybsbyS84f2OFESQPIF
a+mZk+dRM0BqnPseB9LIRBC3bR/hs9kT4jQ066TlnqtI81UBOnO0y0zG/aVaj6a+knPw7VBJhVDz
Wu5nfwIrjf0unxSZMfvKPotNzh1+GafTvfO6fIIxq2GA3Q0OVt21g1G5zkMlRdyZB/+cKZWaGbDo
sI/AY2lQmXH1rJ41W63bGAuLYJXdv5TJnqAIxpZ0gV8AIk0tPrUo3wgNxV0pIieBWyyF139DpflQ
7AOA4y5jBVnvRtKnTVjghVYQHDy3j8gzxnt5A8HloCj/GqhDbQ/KCAZ0Xuv3yevIcplrLrt/3jxU
3/luT0j4hy1xCL9mkyOjzhrZASpWBcU9EDe3h3PIV6yNsiiv1gO4LPxzk/3OotT5EiVXanowzAuJ
8H+e0+cKGb64aOMxxIjBfTkYSNrX+MU2EmuL8bl0pKYzSas4epOtlLYGQss4xoCzqKlph0p3LSsV
N6Yac3mwN0GAvPibcis/HnixlZGG+mkNIWfEy8ap5w8M8ffydQY6sYilFNONNifi1J66gloFzEXZ
h6WZv/PfhsHLkDAkede4mGAnJvDtC2mDOG2noLKQmJY42nG9whiCHFNbyKsvEKsonOfBkBL20lfh
n3Z3zOFUNxfAnvqOdOGHmH4wyROxLwwrd2YiBtOv9oZy+WSLGjkh7oL6Er0w7+Ai2sf3fqLkz7RI
1bLWgjvqZ8/rrKo4b/ZrZ3cDFiDymoe86zptXXaaB/66Osj4MGzBADNejQP58G1+Mt43M6wtIquJ
a/maEl3ZNkmGfLRvp80+64jQ7RFJmRkvdHfkuu9zJxA+ZVDCKwP8uPVu9hPRxFDem/atZ38M+D9V
Y6r37uT3AO/dpJ/aW7SkVDEBGZLLtD8q4IZycZaUcQOBStmPR9Zss5z2K1+rWYLDzaXi8EqeQlfo
FqjoEEHx4ZCIEkaxCs36R6BiRd2xb+vXtzDCbC6Jn/17iIkNAn5I5qWkx+rSYe2KpPvtrngeD0AU
tsjcAr3iLOXNAr+x5Q41VnRScIOfWHSw0AkSnWeTQTWlAkWw+Zaf3o0Xc2nIY6NIT1aXoMRSCf+H
3tGWCK5p6MyDYyBJoS/NBWCIxJ/eI2J2B+VVo6Al6tH0MGTZQQWgMzZ2DSr+aDysdyBlUKlcAbPR
Sf8M25rXCcNb4k5NJY/9BxgckY0flf/yg69vGS0U998RjzIctzpdNCeFJSYCnwMhucLMHm3k1VrQ
sh4FxqOUqZzi9trALPVJ8KGv79I0HfLXUw6SY+KPFvkmDgX68rt/YraMreVa9nptIWUnNFblpF9Y
dFPeb26w+RwpLM+s03Y3PWpIoS/mR5y2zfvHZKG3sRPpEzoMm2w2LegDDCDzSAUnVO6Ud6aP3hr4
sFBE1z0f1qVjugM87E6mWz7FydrNabdzzWwd6wZC42jyL9LGutESBcwgjWCYL9DZNOSNx0+IQy9K
Q8FzV5RI8fgpnr+z3W6T10luIOzqnWwqJ55WVY7FQNTZ5kb5GEbnXf+3OF2V+afRjSs54P/I0zAt
wtbcabQVH2U21WSrsyvHZ57zEllckvGtcEI2IPAfs1TtPkzuUAzwKAND2wtKUSRjLnE4x45MCu7E
GKi7o/A3JXMHC/cJ+y8wyKq0nI5v7SkfRBMpy+MLgAaCXb7OuluZKz2dLgDILtWLgMME1SUY6rQL
je0Yzkl2oW0bTBMSKrbbC6YF2tF+7q0vnkYPM2ISGpa1M4K6ekpKsBBIWHx2YzwarTm5N7de4lu8
i+qCX86MeuWmtj521J0BJhhO17swmbEhzJCLq5bkg5ooAbAadUA+9s/MYFagUN+duZ98hqLKzwa5
SMlzK4XmQClD0XZUUV4fxyzd/dju7RBNE7CKfm15DiFRqeETWv3dbsQsC7sUdhk5jM8KlnMf1Mq+
bhRlJNcEZ32ALawK6YZWiVZxIL8UCxoXlW1tjgG7wqN04QJpswMoe0Xjz8F/uy1TkskE6L9DCaUZ
OSYMuXeYgqIulQsSG2mj6LfycvWm5pD5TTGq4rOXP2TFI+pRsMf2T2I382GZCo7H+GobdYGvBHQR
aEWaUWRPXyLpVOMa+GA5grsWc1NSfzjpUDmxxLS7harxZcMLTGoKsXF7TPBJgCzECHiDvPzCByF3
D+oMs7kG7OQbH1H7iH7q05cTxnP0NpGk1gnigtqjqwvdPvaLiVy/R+vPybNrTCgW52eXILdURGr+
e4j0PYqR2FH2BRXhxL7AZTWtSlqmGFGnFmqQM6F6+7pIELV3G3vQGxpHhlKzZjJt1wR6S1b71pw0
3XNnkla9Y4JKU415OOK/w6CC3WRTQsdM1ZLdiWuhnjWipy+6g5pYwSkDiwYa+3HMTPZeSqjQlj7X
n66i+WcXir+iRa47f8admGVQR3qSCtL/s1EcAqLpnicEDKYMOVk4N4Vf7qeIIbuoPUVpj3Q8IYh4
YKCUuBnQLQIH4L1CcbmjO1PBbl5MobPQW1ZsCki6RpoSN4S15CTsuPNfAGO6GwI09C20M01nEHJa
xp9Gb/Gb4KYJkkHub0fjuqZnwthUOJ+RcaPqtljXIws8zGbtM+J60pAU3H1x5bdafhjoM3r1l1r7
SSPLeY+9PjFRs0nte7n7rVslt81oezd+oWm1UzgBAyXUlbNAmivIAaadOa5ftxH4ea7Bk4Txvx/O
9gKmLyWtss2BP0xf7MV/COqqCsZ2Aa2hUKEEVtTuAQf9sRttEQVHbc0xg/g2eWkPwZUJ8+UPjwQN
jXxs1aPPcCxD9I+pphRed8+STe2B1QhaJRUlYDjQqDd4YKO5hOm2a2WHawZRWshHWk9F/Y5D/I6E
YDwfG3ILn6NdKPEEEg5cfdQNycQf3ctvL0qAvP8A1c5SxNz+Nz2TPzHMBQvFJdChs6rSPEUy1Cxs
rz3UMXZBomYuGInUP5zbgCn4QqxYXTO+fC72grUq2DeiHDBrFwAz6RQxFbAtET2DI++SQIr0rKz9
6wfbYRAypsiZ74LSAKfnH+7TXJQR2XTjBmJLzENq7qI74+w/8zqtAViPwWRuwZT/IdAKZj0j37Mf
hQgVF4n7kRovvq3io1UQFKTrqvj8v25Rc0gLUJ9uV2OB6Pybk095WzL1mbxFS1GCNvV7OdsFZYrf
Joel68gNWcxfSkuBxtzv37qcrZb4bemLnTOD1vJzL7ygXqqWAW7TLTPY+UGVh5B8Em2zW3WOUWVX
zAoWgWqUGN165KrryniJY02hYfZ97SjiMm5sYlWPD6bt/MHIkAgDN6xqa4k5c/k12VnVloH/CrSS
pA9Rb1EbKTj7+Wh0ZQ0HGUx0BmXJMfcDRic5/zyeKE7hKmWKvGgrZCpxBUICH3fI6LUFTTUv4NIo
7RZtyjrXW/bAThY0Vz0mqnMStl+5I9bWsfI0idzb0iBc1n6bjuljfSO+IqKZom/jr7Uv7M3v8pr6
jIh0LltI1VaomZx+Uz6+Ct4ArZ7OzaA7tAci5fpftuYUUHs+7YB34WHLEwgPoPNquL5xNza2jX16
C7QX58CWXKreFWNvTRBPIlmYsdvUEe99qCqG2FDHsrYyygF9srX9wrWu84ZmZTZuGih4UF94TUU2
2EW6pvBWukH4sFYQG8P7ySn2XJwFFk48SWLCHlwGKtB9yKCwH1WOPEzhjTxFIPFpjiTOPUOlSvym
3etCgCpbR3GRgXlZVVntlmOTK6pBDstpL40UR4RHyQFrJl9Y1eA2MjNstnnsoywJYejEjHQNwIpx
JZilYM8dkEPCR7snEUsqaAm2Iuzl3E9d32umL2tpyWUWpdJi25/YXV/YTS8WD6SpSthnea7ck9vN
6GWuT6hKU5glr2kPvLUuPMXc1ON6B/75v8KmDBeSYAiCrU3Y52Gep6YpNP5/L7IKMVI57EeszV91
e/Hrq8L5okvYJsutiNwAl1RJ99+9oEm3faqASdxsZGePE1+CMpl+6N5cCch7y+57e/MUbBSsRHz6
tEnp3qHrF6Phzphfm0ifyBmRjJ0Y3EkZmL/WirNvO32+5hTvDSMyJSQQEkRV55G0eSl0QsFc80EJ
q4vhiXiK5e4HFv68WKQefNqY3iwNgyDyROQYmtbgf70CiprFUi8z8NcDofCUWdLlPXEKpXUq1Vk3
ZAcNf0uc8UY5VDDZChQ4egPuJBd+FwMTznQRFY3nNCNKbgj+tLwsntKTan0RTp8OMca+T75LwevL
7kPzUd/UhzigS4qZrGm6NDBGVVzszQetekCZklg5MurJqWxWbRat1AtYBcLN9BvigrICG4cE8Kdx
x7LRQqA1KNQp0Npv7JoHyzpe1rYO9yeZzjb/26rIxYF11sqKu/XeSWRMOwSZ9bm9bBhcMR7mermN
QWhUryLimM+yX4ml0DKIdbWW+Hw89SxofTswzPyNbJR55sPM6kNQhyg4vZeO+Qboic56fOjDcsJa
In4/IiD3z0OuZPmLr/xrVKLfwbLFzST9oaDQEJwEVX2xIgunpb0GocYlskrQSxH4vfYPwFdb5x4i
W1IUhZAcPtJcVO4Q/gD2emk1/gngTmrejOQQVLBP1XPJlqpL3KEWY8E1TKdyFvIsd/eqAnJGhQ7X
w2BdLdvxEWByrthR5rs/ikLjtj1a6ASG8S2mLHU/+innhquMiDbsqA6xW3TM8Nqn87AajTCZ1ySq
JD6Aa+3DPu3Y9lk7ur4uqTPgPGreGMnAX2K4lUOM8X/YLmzg8isJuHpVQkA7SOnSS29zDHByerjP
jRrwP6eWgBxT05RUmXSeAzSCneGFqL34WmnyBxvAEF9R6EZmzTwbAcTrjJcARjy/UOl6QwWQxKMm
kkSzlTTm2/6i5NRs/u/as3ukZUrCh6Z9v798y/t8rgG6PU4raG1P5Rpo9WLFo23mRpw65aou0lKm
7+lTqKDHEm71uhqXmleuSlrkpj2aAQJCs/+vaaljbsLb4b309ktQxzbSZ9118sWt3REY6QpRomLu
klxIdjozEvnM038XdLuNjTWRgaPxE4MXT3EYfZjm2ZimFwnHUZbeYr8+jMbU/BUl0ic4W5vSCFxX
yhRCzZvx0AiW0bvGhhYofxR4XfILwmzrSfVVOGrlCHIaTNKAnelXE4eWHeXYgoiaa48EbVtzJOW/
xeU2e4LjVe+rLE4viICxdOIu4MIEj8zxPVotnexFMeP//6gbRzeZ8NUIEIohHXSB1dljl0xhgTAd
9dRBcgsusOSh+W4Z92jjFCkmzFvQfvNkMgO+bF/T/VbDcG1WRCdlUVQRT6JPvcLSTvvp8OK1S2V7
1Gi3bmeVqErPbxO7Q1yqJ3eJ/VZsFuCL0+i1SPGc/weYxN1kbiZmrD8bqT7o/dB4oxNDzlIcZYIJ
tbW267surrYsGzjmC99bJMlA6Vu0TE7SRQ6ykuf316Isi+X5XsvH4dkvNpNQCeWQr2yJc/tlHjwU
jwuCH57p2mYzJbGKegM82gHdq0pPbLiaSNHoAvpA711auzdSoVhkNMmicWewFzXPDuxgs0pRkV04
qHu1VTtZ2nKGNIxUOrcha8ddSu98qgS0t40b7Timhbv4lZAuX6qbDWHkH4btEPpJ73OWwIM8wGIv
CAmIH2OpJtLhVG6acJqyHzKVyUP5C7m6IQb4Wvc6v7X+mi50WxumiPEBVFyrYn5BA0wCJC0zupKn
3bpCH97EBxl7+pUhFcgoRFVCaD+iwzorE7fzQeUKHoRgnxNfkDHY6XNUvHt+OcISAd4Mz3sTb4lV
TFiSJiChTTKlY/M8AHO6LEy98g/EGIly1dggo/rO8RpTcsi5A0heqH9ohRKkItXAZ1Pvd6+1lyxZ
4eDrqMXUhWq5PQ1jhBeo0FGqbyyTx5Azsy8Zv9fWHvmvB64UGVXbTgdPeCTSB25lygV+2q0OEf0i
MEQQMVOz2dPVX5zezauJq9z/e825aan2mg1QD2RqI4a4NULZPXXYj3JzwliQ839RPeWCT2hHuof4
AkW0lKS/GFgyI3vLy2B0JssDlygVN+I37Te8OoabBRyUyO7VQQaRoKaYiGHmaVPdErcEikLv6nQM
3FTtLYA5PadsBYaUFs8CIugK1j1Vbv/WCRVhezzDj4VTRQwHuH5NDMSCVUj0voaNBZ73IASwqPJF
o0wfhZogqY2NOoYgKl9d1WN4sIjbHwQw8w+0cPC0qrioFmsnNf9OZCi5WenhIfchhruESbhKu1U0
WWuG29qWG72R9Kd7qJp34smZwN3qUxsYt3lxVHB/BUYejUVw6+VpMzBfXOpIExSlC1gUVArNeSVU
s8Z9zULFIc4TrFY9izaD8+hgovSoWU/jIpPCMoOKNtyNqWqIg83SYbVH//gILFJDfl2F+bvRa2j+
xP7OlzpX7+OsrmFXtvHo7nha5mVqMvF8oCLDeYAf5tflM44y7oO4jDzVsc5BcUT+wJ4R0nG5ddp1
c4kWN1d2FZ0nDE7tFMBH1Rp7a97sZxaJm/2kSs6+KaDMbeUu24GLpZeeCv6YBchrN4DOknN5gTZ1
LuGxvx2RnemPLhU2Cn5fcxAakz3DP+VOcnG5t6411+P18drlWUrLj8cyUknD6Jbi473NO1vhOwFR
caZ4pZdKosfheqK49gMrmDWUjRSFzc2rSUEEt3kbmfcXGT3/Bj2iTEF48kxOrmFwaA/6tXMbuSV3
UASM/bQgKlGCDUuFxtJUEC+z/KNU83UuAjoTD6WF5WVelGGUJJLf1J2zhQMncjwKRcP8O6dv13/s
6gRtAmguZPkVniqKeT+r+vRkHpUKk2TqCXYXmyfnyGeawKc05N47k+voyTInj17p9pIWiCzUQMSw
A6S/Yhj9X1hOhw81VGh9m6YAuiIb9ZVDQEsr42dnHJpVfS9h8KTrjSSZIodqFi63s+brzi2HsM3l
RnIv96wCTFKZmauZR4cWbceGLlljg5hq3Q4hYuT4WaWWHZ5v+BwpIGPjiKtCQ+KTB3HFTIm48UUq
/2xIGpbwsBLmyU24gJfKwa6KG3zuK2vsOe8RkGkbS3cgUKJzyPt20Wjdc01h5cIaNuBlJPkYmOjA
ThaPsNJZlrZNOFDZco5htG6fGj1eQZERQ3REUIYfeF21BCyEI/P4qm+HBXn5uiNzJCYefhtRVlTv
TcgSEopCD/3vojhXHy0lgDoOg6gtyMHUmsekagFmWJBYbcMyoXmBGEXczigQ5jWfPJZ2PebD8h17
EKjnvZJwEITbJ7oFDl1B0k5O/oHKysyif3igAqpHbVQKowXYMqLWpn2LuRJDmWCiLoqn+P6fm9Yi
w70S2vFgK2JYzMqZlmKp3z8hgHZibBqZCGDnIATLaDz8u44VfZVjzCdmle6Fu5Lty8Jin6HVwqe8
ndHjjc8qqxy+04gCQxiRPJmLWuipGvVtSc4Xrsw1EbBhIiNFJudatebYtVTEAU0nfF+mQbNGul2P
vcs4/lV5gWKQQWUwayvrJE2ZWuOeYWbRPBGvCk0NbQmT2ZoFY7XGx8Bk247wTdQKGH5DqSRfNkmF
imPQVoUAxakqFyMUWuI4legl6mazlKjudFE+5rioyq7/ujBvgUb1s3VaerfOMgTXny7HIWEcrQdN
cjI1DjoVM1p4tKoKfyI+DH4vlbQ7adD3BXnmRhB3wYr5SejZo+JFZUqKFALP8qTqERCn4h658Fg+
tjjk10ntD8TZCfYivfXJYxD8A1MRIuxWK9lIbqAkQ+/rGRFgG7CmyuQDfdokWsf7uD9ndUJMTT6O
7WKoAmUFhgEptuvyb9AijvQ8nM+OUvOtsxLqQlpZJFXAUpzK8b3IB5JtA4uMBhwuT1xgdWx1NNGP
lDJsxyf2+mOgjWGP+AY8kCEpaBSUg3YavrUuDkoKKN+fsRLt4fjNWFqPaflOBc/WWArwBny+vkaj
OIeTOFjN37TTg6wLI6XGJ4AZgmHycZssuiZovwR2senZl0TtqNHeT2aa54FUpCdQ+e0dWAtKMuvf
zceyNNqD1L9pp2hZEEpdJbCA/s4+cPQDpzwssJ0AoMhC1E9wPeIIuyFjCJyFzr3pXaiDsdp79+aM
1fo4ggOKPuk2YZiTeR6m/n30N0yu1PnhLPzlQp+QX/Khexe0tZ+Yz8u59vQPpCJ1NXFKUVorm0En
A/5NROffVXXF1nAlhAdmoojiE2HMmBxdFYp69NOXD0ntW7YdJK9oS6J/Ft8M1BUvncX2VRZv1dXJ
vRJqHV22S3M6Cqmdnj457O7FfyHT5uiEH/cThli+g6P/fRKjTG9c2rgQVhlKkFkZnRXmR1vyaumz
+UKOwUBJFnyWsg0rQ2UgmPVJwW0/d/2hmngsWmIC9gZsUu09XnS2a3n+EVmiYcPWyqToidCTJ7bi
GRjfLtTSo8ByBV05COYVGqIiMKoamZummdS8A1ooFiiZqflrxT/fk4jdO4ShhnrDLqjRCNLp9ayG
+sPdYTfvZN1X1EBtuHW+K1sCaOy+YP9knBGXodr5Mij8UZpTQqAMp87ZnUqIYRC8pM5xlkfXtN2w
RFq4CI6IfXuokuIaz8QysY16NrLuZGGeTA32uRigXwezMuv+8n4ElnseiJe+Okh5GJdaYjRqcNDS
VSfu8pltjkmvO6/Y0oOSbA6tLl1SYq/dxCDkKTr1qOOrxLP+Ei6wpbRtn4uMMb8Io9/6rgAIzZjS
jsrw4zkZ63I9I28PY/h1C+pllIe+P3iTDPg8ScerUUmn174rJ67vfKGmw3Jv8CEjGVjD4fI+ZAip
6SQeYOD/J1dWIcnLW9F1FTIt7tEuySrqG+rmTIFNJwtLWpjbXoGoYgCFFeZB/sC9q7VreZInroes
L4DEDmyMoOQ5YwNIEu+6z9NNRiI+1AXkypjpOuvmXzPX6OgF/RIC/uetT2MzVW/7yzR6JgkCW9M0
C7RBqHaRp1eORw8bRYcp2yH8cPPC2o4Fa7EqypxT0/I6lVBe41tjt/EvP5Ww7jchEEOMmEt1pCwe
6bUvYS8R9uGsCwpbwmiMnTRaGYsxYwMHSus1P4TswmntCgi3DTXYFJy8nXHEwATvg/JkoKVA+IJk
WCi5kpoicqBh1x6FHtG1iykSJByEQq03cXYkNC/bIT5n9wJsu6+Gl4RWrs6Yima7VRwbe1aN2BnJ
MyAIeqe6347G/V+ATHRSiwDDhfGSIP9u7cwpao4+sE1D9u6NXetbOsxd73NLYZm6hXa6h4nlHCYT
TOl44tJhqhy4YMowDmGOVP2YeFP5/favDPucNSeLeYF5qTSTX3ijZ5qRxDkiCu9ijq5z1Yl03J7s
+QjOWNkD6tarw7zbU3R2YwTRU2tqrs2cAooUOh+2BzqVYmiMO1KjK7WMoR8MRKyO4xkZtYLYgGqM
IJ4yVSBHUJKR66dJ2yC9ZbhGQ+UUvnx9cOb8ptMZdZSKX4n9GDiCAc6LdtQpsBOwJIDmECDo/ypp
DZ93Qgn9E8ywQC3qkT0wP5Dsv830ZG05IDBuNNAiRWnKxeX8MTP8MD67bAMFFVIkFP5vJMxwhq4J
hFjEKLM5S6OzHf8PIGcgtnTgencQqbWzkzYDkBtFxKciPSDS/AJSb5VbLVu96TN+IJYlprzrpliD
WV3Nn4Rm5PJDdQotQSnIgUqAdNRgHr8gNzEETAdLoiSL9OibjzrwmGZ1Mn85rcQtyuVdm9SgreRc
WzD+k3BW7hDIoQtj8gfuZHoZRa6p1GIoFohInPT4NXUS1dz2So5obzfB8hX2P9kUOUimQIw//ENd
sSCxUzHL7gDnPrUzrewh08u/Yj84NpAJDvcXW6JJHGPOUFl022sVQxvDhRD4Vi8j7/ph7ZQDPNOR
sH0ApRQUtxUjwAvdibwhO7zJQtXU0TONHAe00etUn8QlBFM01ekEWtvZtte3nwS4NOxbMXW2qCfW
j2F8dvuLZ0sI6fzND2JpA64vuvXH4/K4i9KJm6Yy98yc2pJ5V9NpLbDZz9vAGMZv565BxoHEoM3y
6LA2qaBhSw+vNscFm6ti2x4qxqKv2mamqPVtZ4qqZvgw1FKQOOiIRfDeFcSieN9ubA1cZRFMVWB5
iz0qhbRolcl42AVsFmVWE9luDspz/KGKgqmwChZv9X7k/gFHICWY4t14D7fKyV5I75jkyV1higBM
vfXSr4ye02Ih8+ln7xh6n5wqwvGBqFwSHHJFYP5zkeOWHiVo5Q4mUVFfNwmqX7lg9v008h/GCjcB
umN/tdykjvK3gLZak9Tcj+KSclnvZeRvbY76Tga+d6Vrsa2W8DFZ0gCWnD9ReiMVYLrSY+OVzHWe
fWW85hEkuAEaqNivZflZ33E8qtOhW52UbsQjkg8f0nPolRrufMCpyTBRuawja9MT4WeMlBpYSkzk
LEslZPaMuz85KAjCVJlSzsaQYQe8uQoaVPxkLY2DdE5U24Intkno3P1iig0Ti8xb6Txn2gCSB87A
/211xRRVmiAHUeN+rOXu+1WcV9Q7oUxfPsYwgnBZOq7a1cl4cqnA2xFMmlqjUq82kjfEaWBeMd8J
phpeE42DNThnBIJdnY6YbPWJue+zX7nyD4aUqIx0EgctP2iLOABnRxg53pWFCzhn6sYspOv0OJFz
CLX0lx/w/q5iH3zNs9uR3Ef8gGKiSkDHrlIKk9ZyfA6m3sKkEjfz8WVVB1H7rt4vAhHj17hTYfcq
caweMIEroophdcecqbK1XttC3uSDYIumKztaAPFbNARYll7V0bObBjJ+wXpON2+HfnFyrfUugmX5
oOixqDMyQSZUHYA1b9B+mX1t6Epzgmh/KCrH1JMgPOs54NSwXK8pwdD/jMH0jr6VI/JZ+ZxJBas2
PTizCrQVtM/fxDVBjnhGGRZL4OwjCILqqGH+6PUqMW3gLPRcV1ZCYZlLkBg7QU6QwdHsZjcPtgoQ
CqjjXhtJiC8zKae+NABpl2xypOYFLJMIMsjGuXAm7F6QQXhg/YA4X6d3paelg+LWned6RBfy7s1M
wwC1BMCG/kr+BdFcb7Vma0sR1UkCmEbsMl+vEFxOAShrhwIGsLBN74QM9wa3et9dsAC7yDBzzHLj
kpBW1tTegSoiTuEVPEiIVVlUcCW0jopAEhFTl/sralCX8A8XuVGX9Ci4KsFAbJpjrghqWbmzNIbN
ADkCnNEKZtT+6IxV6Yah2aqy1291MVYDWtwp3EwkEjGFXuN4Fu/fkz2I2cVqSCB9TD6diQDuovtj
4uj4R1MUiSdJYH8vgA8uFWLiGrmRxIlXmjrrLkyRSqZTRTLQgly1XEeLsHYZ4Oi4LSI4zPS4wJC3
TpZNYl8zOWPk8KXdtfsRYFr0abogxg6FU0ZDgbIhDPOdv9CUEYTdp/S2jGRVxeYy6rNcJJbFH36K
Vle1iDCgG1ZM5oR4CnBT0wKZteLXUl+KoXA6cNTW81UMAM2J8MFfgUsy5Msxpi01Jblg1A+89H+E
N5oakDX8MZuqSutiORxacvvxQorf/S5Zq+dBqDt/EPoaTNIV+ZGCoQ7fHwaWrl9rQZGhyTXRFc8M
ymCfUYwsytc1H83hyLctF5TDq5tkw6j1RkoAtQPK8eZ0yss33nu1rmbcB1Kpz3B7wF3FoKGSQeQB
sG3co2MM9dx2Ji3NHztcPjiYoG26lcBHECxg49qKk7FQXbDkYEB0QYnqMFJtx0ck9diaagHT0Alc
GLlEFbj7z3AL02f1sk63e4xqSKQXkoahRQVgtXswyOXcczp35kiao1j0NLyw3uyovf3qBVRgZanZ
cR0gHhYMVpcmpOkvthkyf2dYSrywV/f9leWbU6vBSrBR6bOXMmbq9cpJRJJf64LpRSWMoNUK2she
5VcXChjwd54CW+QfEirkQqfleLpko2Yyal74IBMF1keXKU/5Z4fvsaSKeJz0XhfoO6Wyw7yY6AO3
4gPoVBm4fIdLT9XAuR3DsZJpXBB49ysCuvfz+v/H/74rSlwHtl3ZWJS3hBUsqiCCpum0N7dlXeIk
/b/mqObjW2YoufMlWx4rWjRSX2JIWcB9ATz7Qjz+Uj9EIIfS8P900fr+tBUqXGgJkyIoeYXoUJQG
DakM//k1lAseESDZYzh95dQS4ip+8Ghn1gjm/JdjpLdTe6pK31NmBFhnqyL65yYLCu4UScM+ehNO
jRbW+Sk9QzOOkdfyvnD76Mn3edCptub8ZwsbO9faYevPKbPFGtzF8kJ92L2knPteXkjNWMcuLQT6
UU82EnX+K1pvW/LZRCGUDgjTOtQSK+4XkjrYk9j7TjVOvDdPe3QhWO3Z9ESS1LI396Y0GGP5+uAu
HuvzNCVLiu8Wmwh5hByAK3WgIahDycgkNw96TzDsGihRi3lxoV2E2nrIWIK6XwdsVPLGSPJ5xmVP
tuj2gooNxdfZDMGGIU8Vd8425NrF73iRFWyxzrLiqPZYqkB0ZeWoU/Uz16MvYhrCLWrf9mGBPZRI
uCF79bEFA7fOaGE7RDRBzACYc0iByLr7ftQPT08VTuRt0isHQkL+TeI3qJZ4QFy9RYrxzCSJP+N6
CZRLcD4odSfqZdMeFw4lIz61sm7BJVAHFBOgSphqDA2e+Z6aOVmiUt1zvO1FNFtcSE5q70fRSAe5
2zLzOJNSgQemlvUUyDMMBBJoLVI1EwM9pLMqzgkzfUBeDuOomB2XY649MAuEKGvlNgFA8ZyXbvkQ
2I7mj1Sxacf67JdObsjGrVaAPnphRsQXupTxp38qdlPU1Jl9sMk/BcNxV2wHvG9aXujEf3MyuiTo
5Ac/3fzEwWNtFT6847I8ec2Uvr0m/JmAEk61POSgNUUphc8flcfvh3sO9q9pWl3GBC8oZ38uUzHe
hnDWYKy5ocLoJbIAnAtHkhCQAa4IdqfHcoDH09Xzqtw27gNS8sioIT6NayUD7RaH3NU+xKIOZtX2
gjq6CvL0/W8duqfzNhpuVjqicBGOl/F3zFGX73DLtgTseco7iWCzJ6LOlkUs2HcvkrDQBMUQYaCd
C5a9ZkihyhMUqb0foB78jINkTuFsbEuarRq8MOfxOfetnbtGoA2IkA94mjr3lbdxGfkX6STgyllT
F3GKH3Xygr1bC7ye8VCxYSu6Je7J9L/u3wT9zmuM8T62GCUSuC1Xkrc0AT7w96ZcfaZnZ36k+8jU
QBdmkkwOXfs7krpE9CmmqH4Ru3psQzvFdM74CPQYTKst7vaZ7C/6VPv0Zd7jTYn6fS0I/py3qJIX
oGhDxTbMG9oR2BPOaZ/g03A7uxZx6PM1eHixwbpyzv6Sdrlb+yC0tryLMNxhhAsz2YVRg5uHn9Fa
GJoUZyPHk8G4W1Fl3UFJZ9J5tbaYg3aZRZXlmxUzq1onPDxUEcADCyN9/lX4UTOJkTt2xOesDyKM
OT+Lg3vlcdotDW7VAtaYbDOb1AdHWuTZcjiSUP40g+4DdnOAfHkX2TE4HOpEzIp7X5RxwiLmOzYc
4QtLvOMZW2XXAr64G3/vJX6did/g8IO8dcQJU+awOpusgbv9QGhT0A6aUCwJX52v1lshP1Mb2APb
3YknHin3v2RJtQWw5FjSUTZaj2oW52P7o+7Jt8gK6bHtnJ9qfN94go31nY6ptmF5cwwoj+w/EvMU
VgpCyif2Xfsbt+DJS8ehodFkQLifGbLgA47VBksrfeBVJMHznmGU5KIBkSRd6DErEyhWIIE20/w9
QK7TtAFRex8EtJp9YF4yzdXc3QaOhjj4Hu5vvPG+34/fv03DMelYp6fsDBAFKeM/9Xe48ea7R9AQ
zfI4FufHsV8F+7eWIxtClh8xUNaZhtoUf4bmtxk9gHtn5sLf4fnYsuf0R3UYk8G7yQkx5iRj85k+
9cXfZkopOeYB2obh3eDMNz6dEqtOi755ZVK/10Cu/l+eVahKxpQzetmnFHRDL1HzFdWGe0m6pF4r
Dzt7jXg4G4ZxIfSJqC5x9QTA54GuvNgEPgqVWfk9GU6xdh59aiKrMX5Lfn/P+oQVZIJMXTwYDM2w
WjomjwuWER1I+UBup8MYLK8620gTG5CLDAeyIWbp49qR5AUnG/RKkLl5sCDxLrk1B9WTj8ZS0F/v
obZm9GXJWxKEpYXdhuC3xG5cQtWPMR50WKUqiAbLU7qyljP/Rdt3DCzWfHR8Cb2Mi4CHiSVVc9mh
mnyaZUSDwn0rxAIfgbCWQQ1k64sRBCEIDzDHcUAhB+JpfEeNE+7zpzRd/2FPZKnVc7mF+8m1v3PO
TtWaHRnQnp2G29qdQBatdaghkqJbbcJ9R7uhZayY+9FDSSgLArKPmvuAMdS/po0BhA70Q0zsV/9Y
DGLgAb2edHYlTj3QcunyLyL5Gv+mCQoznbQ0/Yqjndle2lmn7AU1s54TNv/w0uto6OEH8/FUARcj
gP7KJCqWXPzYxPO0zPFogmBRj3HyfqSpeflL+Gj3CiHH7NEDJcczjASsLbD02K9m/5UcnRVlJsM/
uro4go9afKZeTTxvi+42O8XzA7cqpMkZD2/Kr/oFiO/hq7DNrxID2K5YDA7RmpXzpdQqO+YIrjVA
9r8RDklx4ew11CR/knnD1X8AGVs18WgwkI/S9O83A0zouAZ387aDH9I4JzA0Gu+pjB/XCJTVs7ZB
KEagYa93Vg4exktvvGwK6a37CBXZuy13QE9woa4gpRcKsxYTrCVKOaIUNiQvQGLlpUJxCGJL4B7J
L6ysatuqqIzS1FuB/mWCyK+L2eePbsJ1QsFkR2E//2SEOxZe8cuMKPqq/CXWMLeQ1q+5ED4xkLNI
zGbZczvfZqQBlaY7eWhiKkCanrbmyg75tSbs3mjao3Qo9M3xxBQuz+3lmBKABvGhmCinI//zHN5P
tvgMU9sPVVBG1R+XUe1iK5iLbIgnNh5C2s+3Z2mbNelibYbmkfzZt0C9WQoTYREivDiOlEHlA2yK
8AxV3NFSRIvsoXbnOjuJTe8HPVPr9twX/SvHDQSJx+U47xZ7lWk8kd4SI0FnYjkRUqZQMTc0v38D
EqNt5qWlZC282W9UsWMugOkpz25BNxH5euu1VJVDgLf32fzw6LigdHTkvu5Ehs5M66DLSyIx9VPW
/6PSg0BjYwJ4aCGSHt90UQ1yufpvA7XwJ4MY2+PCyplKo+VmQpZR/lmCQPXwEHyt8cmTdDHZ3Slt
ozBmXtoep3jYS1DCfhauEI54+R/RpWDZlpx0kE/XQD5e16nqmC3ReYrfh5ISKGV6nDCI4lK0pJwp
Dn5QJ6jDeWjBAbz44LeOby4sFh9n3cuKmCD/Na2uoGhXUo/H2omGE/WjeqrtN+fVV5HsXNc+YSIz
u4VWdpjylgA9HwPvoGZZjSnylgi4uOZjFujrWNMzZXWQfnmRSNgsKVk2fgujaQqkTvWwV72ZqxT6
k9b2PI3pcVYViHdlRhmSmpwwPiv2LR9z3iO91LaO0CcEEtxKSke348X5TcChmOvGCFHGt41yVC4/
ItceXNhVn1dGxawfSBsOznEUbtHUq4WesOFys5cAygzJ6VpUQKM6pn4WUp5ckmK2fch66i4xelZW
jTe2NqGVHyx59yvN7fSsS8//Mw0u6MXM5nbkORWzxvb42clTj7mcns7YXE0SzIe5pISiOq7yRLza
8LtLL/5TLjlczDWYT5Eaiwg9cg0mRYWRxMKhREgbltwKlyyYm2iTd4JaYlkg8QrzWafoOsYw9EID
VjRK4PkFtZEYUrUFMprry9z51u12+YcV0cRUximFeIcMqOKQA+MFFFTyKFaHKzFlGxzAbbnUeTMb
kreUOKNPAg+NF6c+mtfr5oQt/4tYcMW/1/D+cbpRa4ZHlnLFRF0YDQaCDKgSMh7Hc+BoJ/s7+IXm
Z0RLaO2UjDvLQSvRwkcS7iwKlvJRpip+0EbOk0idXURWTNGahRX2p+04Tm6DtPnKUSQQgJGQdg6o
jd4sL8OLS+C6w0M+BGyeGVeyAwHi4H47ju8oB8X6dLwdXqdbmYYoWP+GNKS5QZUxGSSPC0ltEVds
dvOT7c9dG69f77F19ywfJHkSfmU59nkXAOXz/WTBQIXe/2PIvtlbR+LD98fWn/zkszkdZhyocMB4
WQumw1w2Z+nV8FuTpeDRF+xNTkUF/E1iOxx4A3n+E9ZpskLqKmAv4yNdGy/82LQvMJqwNWxv26dR
CMA09HhYopIuphYmPCRBNLTOrlTxx4jHIBTADI7PmGDTJZP7rhoEOjJq732DqMy89GLC8uvZYgmy
eZuuydR7G0LVfQtahwP9smlR9tgiBB0OjeBsIlM+2v0M1T7fWdgoTBKlpWjR14ujaUOd15S+ZPNp
3MepRRzQv7cvY5MhZ2cqxzXTF/aVJIXosov1/8yr2q0HpkkwExsxcmINCBODRZlrb0PxYympiHtm
B7OMPf59HHYO2Lc8zyuKqH3O/WgLRYYkQXDZPhBaE+Ept5cFGtDI+6jgI7tFRS+nSw7ObBqGs1E0
tn+I4c+qp611j4MX9xbUSZbVT6kOpwikgMx6kBwg0RTy67b9GoHxiyiKPtvxzsDnRvbBI9vN6jQE
IAfWsrVtgg5WYvvTNYo9gNT2lQtEv+orAACYXr0L1qZXGJcB1wS/mSyjGA1JmmJfnPHtpTzfBgqt
6aI7I54vU14q+oveNFY6AO4jgB68Qgp7xjk+aygaPRvm6W6kpXM3wRsV9W/moJhRr65e1H646D+q
oSZrje5727RAdRJgsJ530i8r4iScqD0XP2Z/Kh99+OlqB55N5AXcG09NvtdznrmKeamlY9AhELg3
V1L/oDyf6YKOfHw6cCNf4NfIgMc3FMmuSimOkFeyAlzyhMnpAoccQ5xeZ+7t12W5VGUTJN8NtVqe
E5rmVB0BvY+lzdM3DHoD8/ICiMZHOoNcyrnP+xhVpVw/fdx+Bj/WMwb1LRppTAJL3/iJWESNA2/C
uptqYg4cYIrmsp540Ghnug6ThPcLU4jg+hjpaaZRF1jIEQODPo7MBr340RyfXWrpZE4kCy7pYkj3
gKaTTavYov0sc5F5D6lomL2a4wKwYtaTeYmz0ciVyN2qdA5zmzjG9rAFu6/gv13JY4Qj/Uv/DJpB
OV91/G4GeabWhftyiJ7s/4qK7WARaw5ZNVZEd+bSdl7lqbDU9NXZhV9ZXGJtu0Yji+HpgnwRF24l
ghkYSGe9fTla8bFIouSDodXJynJYvprOhOi/v52MT25Ewcp/ZNCSjZNRJFDV35StLsxtcMI/ugxw
K0Y5PNqhYhBvgkbE9yI1ftxDfo1qFysjHC9mosJjCBeaEHhWXrr9YM0r83QHGw90KO6IHwIVk40S
wXAXOt2278CpGeDClpnbSxhVT1T/wk7xzWjdnRQaFI4KFPnRod5SgrWHXchwnVDGatJxnNspGsQr
3Wgyg8tx7SZrm3cBh73/QUxhewkeqm0Ygpzszs+btgHJG1dIYTqzKkcrMWC1MDyis6rPivA9KiEr
olBGx2IpGSM9Qu/sQmRlcA5fV3Cic1U09eDYdg7ZMgS62NTcbDJRIrtZ0u3LyAbQSs55wILeMao/
hcZfY2P+77WwA3NswwSDZxHfJxqclE91hw0sBYnH96c/c/nTqwErVvMS54H1uivriCqI05RiBLma
iNPZ5qz46WSYh1dmjyBD3dAdWb4bIET0yY0/kQPwdHVwzrHRUnJmKpxMugsvnMQlEiR6EydNsFnJ
mlSwZOEHU4AcY+nY5JS/yURfGIDw32opwtd62JJRcbdJKAr1VRqOR51unMARXhuTt28at5O+Y9vq
wf13SfDLt+hOLKy2FQ3Dwfx2In7LW7gGpm7ZWhShfwb+c2n+HTUZ6q+VxzavKCuL2XiOHiR0LZI6
hrmTEusEZnou8i9YyeQuvjmlY96k/siJtwKC8d647G08bOtDXdWH9jTxMrjwZKeWmHwDI+WFKkAK
bQ3yRprfUGz+1VEytTGn2I4Ut3tLvhpl2nLW6uJ45Cb05Nm7mKzUOanBZrm8P6e9EDwFzQ6zCRom
GJxiuLr93i67HMopIjv6G1Y8KWGFw1J0YUI+GDQuer/I14BL9++e4TGcWITmbIAM3n6MYrWXvSYA
x4a45QjHbf2Cf3EjhKW3sZiArRNMhzAbXN6NmRUgKMwnXuDZ7oGAi/8ZVB2TPMvk65zAmEKt3HbK
NySvp9DbH9pf5rl/TYZd3jX8omkyzMyr+Ixwz4gK128yeEmhtQrcNNhdeJEjp/FGBzWzQP7MaUIW
4LJN6FknPloGZ+NydHgqXZZzQG5t/rK6S/+TUK08uK1JHbbPkn6DnCfLSZnO18tZ1wMo1Zammrw8
E4usEpshjFfcCeoqxiiVMqtvgFwR/XznqAmeixn8Two3/x0zfRMibgG/svaUyAJ+EEmEBLxHd+79
Fx+BIdBd6aCE7KuRB/Q6E+EDk1eXr5r+m63HSlAz+lzGzX9EiD+rhMsFPFNIE4DLvlI85kXO6r/i
YPzisd9FEbEwlv3tjKu9I973k1+dvn+edFz7EOJOTq6/90YhDk8R6w2c5CNd0IFOAAv7JNDwJ9c6
fR451T0+Udnb9XyliyIHHSN5cpYDdz7udbfgZYlBY7DB7w/EnV3K6MWQH8vi/2FsJloMDlLMN0/w
QSmSrj2EJb8LdMWO/Edye3AHHq5ykxlhfd/z6SJ0TvlvIhe6KT+VcxPVLS31JJ1hhXtmqBlZ6eKt
nxzjrpXlGPQkGwRh3ep9oNjklosvyqsE5NFsKrPfl8KQdBn3vEE9H2yDynEVbGjAeMnvMQyH7ZLC
j5qSEqm+RdwC/sPWrIqyVgqKbfzdZcXuT6PGEWRJG+JlhfGIiudFhgafGzwfpdxfnL11pceybHuB
XwMnexklA7ay3bDzC/msFq0guYkgYd8cQc8c9vGfBCXGUA+SAbburDb28REU9dBJEhDi0tbylQ7H
py3v1EHuVtjS4E0W3oQUVxtG1kUrruXcWSsQAiD8UFEs3IxADxvZWXFS++df8jGwN266wz0tgtxq
r75tirYeGofq+iGs3pnTCVhN2VYkKft5dvAI8SfYsstcDIcCnk4sYD8JhPYnsgGmVOgGqb8fbIjP
HTFqTEE3bWHIZvxKN4kRJB/Gj+nPVkb/deEQ1hqZq35mDBp/ZLptGCk9lCIaLo1HbNXV3YSt92xg
TPaKmv+VljxJF6AyLPK7N3Iy+hV+2ME91z/uUrt+H8UJEPItui/PLFxG5+OD9BlKgcI1m+zSZiUQ
FiekB/48d6+CY0GXYh0Hbc6BiRZqowQm/8QTaWUHpnJNzLb54wochgNpe94XHbBGkMSuSVdo1+uT
n8Puxv2Ptqa9yBePF8oXn6JHkroP1B2zKTOIeOf2JCWC5dO44BehrKvDZUWBbMUeLD52nJibWl28
Mm2S5sH558ao8letvowox6D8YQLG6ZvuO6lZsemlNgC4fD1O5D06BQxYA07PN1SsyAmGPZRKtB2b
wv0r8TjbWjZXwrhafakUh0wedWlsdjXccDQVfAHTUKICQBuh4kznaEPFqxJXT2plbK6V3MK/0Gy9
k2vBUl0SgXL8r2QZYwksaqjF3JuRWmRnw0z/Xc1BIHT9uvffuLWdqNDr9Xymceol//VCHl3Xa64x
O6v+uIszYm/fDZU29Kyln2BeUqnAlPxvQKWRk5agfXWtsiAcO3zjlqZmUlBaB7JZblev2Fdjo9ld
thzyx5k2OkopRHlOy/3NQkTkMlSM4zkG8e7dshI9sqyKcWfZtBsd7oMlqJDWrcuIwe5LUhPOvGjl
ns1iYaJX/piX/VwfbkrHDFVwU+/qhksiBte3Y5JWpirwyfKmkF1nMk4mz21v+qinWkYYNKuM8UlU
Hn+NNhiBW43Wfvn0PwzqZ8F2ADu8iAk9hdxN5kdqLJ7oG1BQLFE40uzzZCp6qfAzE7wGMXKzJ+RC
2kekC4sC7Ku/Y7VBICIX4fk6GlU8lPpilqLJcm6HSbGSsEcfvMpnNUiGRVaUFsu2AzQcdoFaiVUU
i7ouSlews9ONJZj+X7pBGvdjE9z3j5XrXozxBosng9LXWtIlAfpJuiSOBxNunF++Hy9ewu1NxOKK
VeRDb6JHHz6GGm/dSs3LOdLGQr818w7DEApblzxbtkripXHh8VR49XNYbA0n3qRr0mVPl7BJOQ+h
RF5iADlUIbz3kI3mASOsIQLQRe/SSk7zV7s/BzOYGRvtpv1Y3Cmrx/48Sa2yDFXLKxjQDe8SJMQa
vL3OFCI3lBiZyobJoGt+KnXlhem8IMZj7whrw58CxRHuX/vaf4PMrwHgq9dpRksv3+CaHr/kxxXF
gG9gXe2sqaE/Nc7hYrel9vdi4FNj6WmHcow2nziflzcrVPd4sWABjuFpwCGj41VmreVD2Sf+mMAG
xJNInnUk1whukCPXaWOAJMlGTC+hnpdY8le1ch/LF23Lb76qHc1aVAdmhsfEScQT/o2rJenrX9wB
YE3EDuKsOTCY6RKcbFbw97nvC1Gp/xCC/a9/p66EiCaEh0D03kthRm7T9eyLV3XHMWo0FJ2xsSZN
Lj8Pq2Z5RuC3GkoU2uuY83hRMO+zV53SzTkpriPZfysGqa8eJt5sCRFMIRvt9u73NRUBXUiFa+IW
L4mFbZ/hYqH8KSOMSvNkkha2QqcX/ldXagexxDIdOq+smmN67clxAe3ZsCkY+NJpzT6K9Eu7hLON
17iOzJ4bn94A27VEXKbwxYdYF9nsebKUKJE+4g0E6eLuphBY18H9M1i9Bswj1+ZiEiHKBg9UZJqN
fQxc1JU6Akj/nPoqH4OjtzI9wMBcrR6LLA77hCHTDCQBp9WGcEJOwC5Jl0fwH0L9lUmsC5F1V5S5
O2qgr1T/UU5UdVbqaeVLFt/SHq71Bn3orBj3XTpmReOLADvZXvLwc5SVvvVMTs0lYVdsjaD11bXr
Hd6M6d7+qygNPhGU31F6Nzqndyxw8sxnsW9A5YeDyD3IwbQZPmbnYE1FOHLTicvgIocd1z53vy5m
2DS490qyNLo5+5KpshCnDKBgLk3GuCFlRVV1bxtV3ZzHUQzj6ePLOu/SxNp6/Zu2uec41g+Yct1s
U7V6/iI8IuT2IgR7yltmy09SPrHuQxPZ1MsTPJTE6L3FKb3zuEm4s01YkPOdEWaY22/LndCNEVta
JsxqnqUg7q/IL22vg8ECFwlU209QqjtNMPnGgavOJbsaGGMTRb4fOVXcM8xKQj4lmW5RQXIcqt6G
x0Im4rHKi7NM0F42CTAdugkqzcMD/9H1KvQr8y7vPWAbzhHtZiOKo8XcWWOeqmzJBO/BrPFz+5J3
1rim10bMMvDwiUIcV/UJrV1exLpopEaRi+MYkacf2UiLK2LpaZ2D2MxpaiGXdOCdlB+wu5qeNq1F
5wcO2rFmd564VMecyQsvDgZhQXRXHyZ22v5kGnaLJJB+h8mYPV7TGt/RX5vqzMuIDXEOIkFsnzQ6
yj4n6VwimuY2cLOfN0NS2xSvLxd663icloZjwkoCUqnKod2hG11EWh4XmwHFq/CNpZkPN3J+ibqL
M0J7Dg5BjvVhS938Qi+zKyloDw+9rihDavKhqoVnQgvxl48rjtwCOjdGTOtw+ePhlcBDE21ODLxZ
1I6s86xuOZIb3WQBX7eh5AR8Vjd6R6ERffWvVWwG2zL++S0LAZ96irAmGu5HM1hOyUSm7I2vm4dj
d3TQIdhnj3ZNfhKYuZSqa0QD4B9QtylK5V3XC1Gps0m9O40bsdbBHawHaJ739RoyGWMZ3YhxDAux
fliwLmSuqcU67cGx1ayKZ8VfDsHnXtq1KP9oS2QFQ1DJaG8Y43il/YrKL/9apxojBVpXkSuC8HKH
4RMMHFjD0SHn1oc1GjqXq92soQIi0BokM/XxIjryGIYukvQlVEionxHMZxbNTtvE8Y7vlgBUoh1r
9kxCHDY5533QWEwU+tHmcBRiC9Gf4LUF7+2QQ3lDsPlzg+iCUgHdRTktFBF3qVHF5OkNjONc9LyK
7W947+85k5KsEs4TUX8u6D9N+wLgBBsMclP5qtltarawz3KI8Gvbo22biN/i1ycp+728RmSWeowH
DHoqiE8FZtKsrmzN9D88qnImQZUFJ7ntZf3paFFoCszq9K4pLuqe3YZv4x7S2VksGbbt74r4WA/8
P5p+WJkynogX3NC1l9L2sBjvuqL7X7g4/LHt1FbfWHppGtSFkYsV4pMOBU+J5XkZoxER+b6GVlpj
nkRGrTQKZ+cRK2HR59WrutxD4CJxwn1VGwd4BhFlMYO50SgInpKfX0+Dki7W+2qMGnbgj03v5GRa
tdWJedky4TwMWOCctifkDYVRV7U0lFmH3dcWfy7XzfNVSsjCXr0xc2wITxEnJJUbrBFVBNWESgJd
2dCPoItZhoUSjzBg8Et5n4DjQKC+CaF8OOArRdzU8IyF7rZ4BUxpAxRlYb7SpZRx6Thz9yey3qBs
1Lb1RdFZNIIPI/kSvMdMJHCrXslV+BAnN8rQLxSJO0LQv7eFRfGFv7tVlQ3U8aTKW/J+jOYh5Oei
AWtAlS9ldoYyGZUSUjwqGtew6GmmQWfxD/0PoWtZ1KVV0VJqug1OSIteYdZ9FZtkYfwfkuduzH2y
A3G+WmAAjED6zuckXxBDBMC3bxn3r6sLmqHzrrCAvrNBAk3BEGskNB3xkjr8gYyXkPU6f1PkqA7r
2tMupw8Y5isfQs2XvRo886aqzhszRdgOidFjsC3Vn6Fa8+6qq1r+qHU9T0MYBpFgD4IRNELmvS1p
/Itmj0Zx/QMsMDUeF5zOjugdFCsG/CA73IXYL4l3wAzvVmPcV9z/ByiMsf2Edt+Jon5MYwtcGTrW
qYQE3/VGai+FDoN0FtPI7NbW4vThRysZztU65zXDOzyA/mgijU2JK+8oECmaruG8ik65aDrIyR1E
TMGvlTEQJUU0IHNs7R854zevnPzRJ+TvQlCYKFzy5Oil4pSomJFG17IsRgUMyM5xpg6Lxuo/J5q5
/HWX/ux4SKZAHvtEYINQBCHEOEGZIOyhLZkHI6L/sPpTKEPzJ7vlm/4bafK3H9SVg7mlEtN0e9qu
37imgL+WiKP1PvaUBRTcdL9YsK5vKR37LaH2s6PZqxk1jxq5VxqSAzZfgDJz8lM6CsZnmzRy3wgQ
Emy3BhispZGW0WruA+XwtTEshtQz5vSPpeoD40Cox6Z6FJs56YngLqsoCggkDqzlyGh1hWU77Pz2
CiwMuYiA6ADkPKPOtIzw25PkacHVhHpHGGaU7iaTokGQx+yu4sCaMk+GaMOmSTeUH1RJbF0NjhMS
eL40N3fNvThuwEoI/1IocMqAYNsfnFIhenMTUbKm3hV0k3F40+8qdgkkojotbKPsmRjm2/uxJ0Ym
9etEVjU9RytdmhHEzYF7I8KsYVPPkt6GcC0E1W2uj+tfPm8tiBEqPsNUz7zPUJLUOmT6FF+VSasm
Ei8reG869tTJ57ZY74nhtmzMncYUboT5LCtSe8ujBffNEvNITQ5c8EMTr1H30oIxYbisDwifZsgQ
q5TlhYgsuqGKVvAMz0x27BuCDPo5+eiBQJV//jMxhgCDIYbw1uBMmLjV7bMBMvwaGHLIyzst9s3y
C0lb7xWNIfVHlqJZ81INA9hApV0k8jmumLi9W8YLuA6uhOyvuy0lY8pQHx0zsY8ejp5ryzDFpd7N
avFYKRYJoI44EE/b8idTGT7itDRF8cRQa6ASOHHi7yF2Wf985Y/VPW1bSZEjmAIlKh90YiMQ8Xut
9xWnkp5uXNx/rxE1jusOqNCRbZS42g6pGtJFIP8Ai617yi2DKdr00GdcxSlMmubJAe+ulHDHwfwh
YKec5Bs/LpbTQiIy54zoCDVGrI2maCBs0Zga5p6S7FatmVVsyKH2Qq8e//1NFZ3kl4pU6lRsSW4h
p0dNHu2YSMY2BqfQ6oJyGv8gKvBExagQjAB9Aj6NBs8Joj5oKUenSRXib4NeSrLkPfyT9Z1gDKUk
P1zYoB+E14UBN5ODmS+3gT9quugZSdDyPSF0yg667p2I+AX3lIOCK5DXS9XfsFXSx/FCuwk62IgF
VJDpNiDrDAP+K84/21yn7/17Pt1l49d6Ox3BENVx7ioauuMz4QyW/rRi4uAmJrAu90XILLIQ1fiF
g0uzPnJkBQWvnVLJbhD7skvv4+aUqRxJ5dxmuTc9wFVXi1qoCz0J3XAlXlc9VLBgm04KRMIGlKtk
5T6VjS6gO3UqQ5PVluHfr1mbryOoQtulIP+Xy93sE3YOxey6PN7vt/m+Rpo633Pn734jPOljQQDt
R/Fz/XhbmYnMqHezR552bmj6xaXCihM40bkrW1jtG1Yyv3IgLDmdtr8qCHTWrqzRBf0E6eICDLqB
y7SwQByMngMZQyDiYyyCHPk9aE56A8nL9HUJthMdH9825AIZo8wOT8ba+PtsN5y4/Usg/XFOLQNH
RDnX5RHpnib6PkdSmE2fFY1yXQEBvvuc83tjgV7G4sn8rjGJPa/fhRYcS3hb1c9zd9UhvHqP+78s
5VTgpaLPbgikrQGUd6NZKd1MVHu1sG898NohKoKOXwXTpBNbyEluUFRF8B4Ok+QazX+VonK93zGX
eyK7iyQQG44vO2j+s1egKDXnWlc5b21qB8k2pigp9aOg6VV/v22x1xX5bRB9FEcpGllpumqiMsJ6
xjAtCAHcPHOl2lj7F590xV9M23DPku7Ej/wgvq8mMSV+E2JSBAFr+L0VTeyoL7BfwQCYnZuo0Gb2
vbcWmTHfpKeZ/RiB0qRrpbZ6opBtLrNGrTeCrdWGbLw84shZKh3hkMt0kfj0IhodgM11sJBvSL7s
Ji4OyqUHSIto+XV0m4aeH+Lwwm9OFWUXaS4s9L7xnaJHc0SN0K9AapNrT8GNGTYjVe/UEqkNcv8y
TTkLXhRatBjZR5qDsq3+lRMA0ZT83YqZ5GpBWL19oKwo/6JG2vogSOF30O+XZSjAaAzJeCVJMMLb
AxnWFzNjDOvqMHOtxAsx8qdqMOrEZIQ7AU76V4gqfNvofg642aA7eDJU5x8mhedZyznhgrKAqOIF
k64gTv2E1/l+nvSA8zOE2SeeyDCI0x/aT4Jqy4FF9jMOEV9OLIQklzKCaMiSkmdWQhPllrbHzTC2
f9XRmwCanRtlNHxGpAAVUR/TYLCcaTZKiEGmBHoax9XYfYXFA2xNTmRgj0M/wCRh1VgzAnPO15f5
b6mvKh2bUQJeMgAwJmpJfn1k2mzCAIlwRGIVt8lPBy1cZQzSsccv1dskS4O0NHPtsSQwwEQHa2Uy
KoGDCHpTRUBHBTUCHChlsxhv5+4NxIhxWQCQ59j5m1xci+xalG1AxuqPVeT46MZ9Twr7IkJ1ZyJN
x1TTnQ06XVEsGLEobP3CP8W27c/2QRvcp/+pIaI1+you5fOHQw+gV/Idw0oX32BEmZ60NmluyE6U
PAIyICuUCxC4h48WpuSvQO3M2gEZubKiwsStrdS2eV1ktLBRwGVEyZ/hMpcSXOO+vkztjbEmDgt/
saujoIc1gDi0N3cIeTLWDR78+wkW6wNkoNuV9F443J8cty7Y3v7lFKKTdNXXTk8DiSXkZ+kE98E4
LkqJuTG5L2hzM+r4REVX18GqCRlCeITmkUkRwjF+deVzOTf0+yI7KcauZ6tmaqHj/EXqhc8qla/Y
gZs6+tA3PryPpbNWo4xevx2x4/E89t5mPOJwLlYQS/LR/Ah7UhYw8RCmRpz48b3nXmapQ9gPMaVp
7o3BK+EEidPTWqy69cIY6FpHDfA6u3v2nwJeyl3t/Onhk2j7n6/m0gZHZhhPhe6ThwlHD6UcJVUH
sgywV6JHmYrREyIJ3MyIapOfw4Ky/3tdyTmkZ3+QHmSHmrfZuTSzaqYZ1oaFRELO4LUgMe35+KGC
SGH0QM1g4hv/5HTDtvgYeCNACRGmMPoWvtvahwU055ThS72g7fdsEAfxHLmOBvpwcT8mUMsThB0+
VwYlx16NCVxZGp2EPeMg+HqXeym4BVEyFDTY9dTsHXZt6AcIRL2txDOnCyqmpG3iOIvj8wWmJwGF
5ouXjKlB/JX06edmU5kdLJVJTjM5u9a/24BFCGwhmecR6Aj9wjx5nN1jJ9I1RfwXsDsgzZEemOeC
PEsjFchmKO7jwmY6XMrgCTb/5tSTW3OYvJ/0FE/T+M9aUrbcErQhYZro1qTcZ6YoyNO/W1E35ytm
kheYjyoumGgWigLobqVB66gVmbszD0/amvGMb5oiDDXetWX7dX4kabjEz4gsj/KT2jxP9PAA89dY
2HqUCnusoGIb/goc/TasiGhPUpT5F84GcxVtGr2+aDRmb/Kzxg8QDv3JegcH9QtgWZO48xjqTs39
5WAjDMCr6r4+I3XYmkpSqKY/BUTQfVOdBctSxE7Rb9+whQp+DDnIJel0C1Mz9WqCI+BjaE81ClYN
w52WQuCqsTOdPHG2mXPbwiTIg1dDJ0RhUnFxqaqJuf1UAt0y8Ec4/Qfsj90FZbqQmNpXrkaOKimn
KlfLUeJloXvfRf0WQae6Ucn/KpX9ZxWC472TGrGdw9lSKP6qjt40rOW5UZTRvUQGWhBqWkewt/qp
0WV5pP0IOh4Ul+/5rBehiCz2+VGaQLd3qTNRQbJER7YoyM//r2dXtCA+/sL+MlftkLMHL3x0Volh
EI/xcCmqPw26bSdQqdOqnUrRSW6VMP7oKZTMZpTstohitrfc/v/U29Ypk9xxX59cnWd+U6c3p7Uj
SiYjLKHNYYqEioyK7m8MywOsCacKdb/2Qk/iTn/vqimP0mp+4CV9pmhFc++pAgqcgh2ZrjPQCfHJ
ThTeU3KaIRZvdt93BvFGi9s/lv6M88uALPCGJVJAIImi3sLqUFpIs/khIg8P/Dg80BFkqtWuxXmb
qg6WQc4ujCamEB+Gc7wlOPIy4L05FOE39ErvsD4ECCUoIQzZUE5GKG+U2AvYh/+gwRReCrXJxxha
BihwYM1MGOzXSX94bMmbhNshgft8rOGvCCpAXBimd3IEhsMDYf0FdH/iPUAg05yHgrdQLynIxru+
/iu74kMiHql5v7yBOZ7wIzsyEfuHYeX6dkKzMNZULRDkB3OW/vdkAVwU9J1vS5AF767JBWWRS0Qx
aGuBY/lhc2C+1D2tRXY6y9vrgbDntNH4+AO4n8eXQcplGUba/4CDyp4V/NdV2YPv1VOBAhntHCiY
EAunFf2IJVpDBQlgMLHCNPQx2MX3XiKz0+7RGORVVHahT/NGnoNg/hrOjUrLbNtuNJCg6ZGI+eY5
fvJ9wFbEdo9O2+2suE8xwrr4QuuuSdEPJcNWu40EMcaajWms8mUL8alK8C817Hl8OeeQB4yJoUd2
msnYyw0QxJ0e6MaQgl49NG2/gAzOa2y0/Qs5s30CX+v4G5D8cdrLJ5w1xFAzcdA1TwPVKj+kZ/iV
yauL7m47GyVvF/TsLtr0mRywnys2Y/WbjBxeV8G8NCqpfQfJUEKbKSnH3a+YpEAOrDTxXJQQNkA7
R203jm958rk0NN1Q0gdfVJzY5R5OW97VlUDiDIWDVoFYysalZdSlnw4GTM5ZH18DkebgJGC9HGTf
YMbBFeutIFf9amAhBSeGjiD4axbDUIt5SA5XuH02zrJQo9YSMpPx+tpwSTK3ZDA+PdO3k+gM/eho
vqbsusRHw421tZHPpG5kSUsjOdKBdEwJl1MA7WgD+DzZECqUWxnKvKwaZ7SKM/sBa+05a5RxdoLP
F7HMzXNQ+CPnleK2wz+xn8CKg+6NA5eNPIArsbvKfSwrtBN6ytQi4TNnYyKi/7Ohm7VT4Mqkhmq4
KpEUIdIrTwIozk2CLxGMPzCer8Xf2J84BHVETA9yXQ+N49gcLb+7QfQd2TjR0DNY0BHonqsK1/iY
HrlxcradZGVFLdNVivHTf0pO5Dnhe+lzqqy+OveW0Yx6bpAodCjIBIWJKqellNpkiOIj19d5EpsZ
Xv2z3Mc42iHW0E37oUm0OMhe1yttoQ2IzQ4DbhWzOAc/NpN49HOTIBiJCBMpxMS8axK75/KVf6R+
zqlHB3rY69QHDAwoiFuL1o++z/f0uAuZIMmCMLv1XWP4YH+z2mte+hrwFxsRB3dnByWwVCIWGr2w
3XsFUmzVMPqA53bRf2vSPmZa/YeLtHGXKNvDQYmCkLNL77ftQvJDJzsFg50xmmQewEIEN6XwXA9D
4BsOYouAisDPWFQiib2a3CnksIsNbRJIRaMRccPeXNQc1GNvz1Ogb70stGHQmXXDv0ShtH9oR+w2
1DY1miEdvuJgJTh+Bak06L4NshZSwy/8DULVTiAOcPirV2tnv2O+0EJDMAEBJkwyvsa+kDCCSI3R
Vx7euK4CH+wcdKgRHc12ZGIVMszzm+0OVRUeG+JORDwCBxEjYt68SA5JwwYNghZkBz+OIneRTqdM
IN9jMvnly9oQMiIIB76AtDxco3hw1F2MbOdSergITg+MHS/yhdwvugdhDJoJ5c/cP4ZliDuyVwcl
zZ2DLXVskNz+JBLFMhgGT35P96jO/LIxHnzaELFS+Ovg9AYhYrCxgKQRlaBm+Gi71hd+IbTXgNO7
VPRlb8tFBsBsJ0CeoRPYyfqkZRNblbx7YFTeebBHb2U4OTbfwR3YgN/V5Khtu3JNBwUGSlUhwmOu
HgoC9WDNVtmTTlH40OWNi5y28mak4rjdkxRDPgkABxeoEz2ZEigv/BiwtM+d+vc+foml1adJbRKm
ULusrF8fqKNK03pRb0zipBEfiYHDiCij/6UtuGTnrmtJIpkc5wthZGTfSMuCx30W0cwvFPr6FinO
l6MYPLUbgmCn2PQiFS3o6PVbfPsZi9fuULYt93VvVeD6/SAkk5hJBlEt0xuAOWFmHgOCF6vHuu04
3IWq/n9Y8eoKRBj9W+rYnNOEfi5HwfP9lA9ri32Srej/guCyAY6ehEUks7qssM7mK+8zJP7zTtol
Ks5m4Men2qZfLOtGChWgwOAkBCzx6ZaVhpx4QyuBKNNAIfLU2pQQcieiGqg7966fN+P7v2dLGXRZ
L71VFUTyYM15EM156T2pTVotiHFctN56Yd71jgWLuwjoTBVa4YHE4opypcSlvHTpGp9mzoNa99+m
aomFDCVB2YEu4/no8dIa5QJIUcX8o12jMHSYcuylcJuFl6KFzW8tTzpClng4/EXXBlu75mlGJ/HF
0XRwe4uCfeaZYn+RB//4qKvL+L3c4MDlcFkBA9mzSpY++tU03iboq3xrImPgb9iyVlZk8RFMxZsV
F7EYthtZDkLE8NEBrZxHFMyOvcuRkA1dHeZNCbeucBbQs9TV9cEBjz3WXXE0kJ0KGb85RdAPAVoz
8d46TponrXVOq8IcI0DnTajJDcrxm+1/buA1dG5zcz6P71IZ092kYypicHI6eyawh0xDamsX4+ZJ
NcAST/eRIGFQXMiH4TLwyg7JhWCvndYUy/AZSOOVRjho3w+rOW6cjBYpYu4082nxAYMqHKV++qHe
3ysItIdr76jOHjYB0iRVPkmpDtfvJScTk8x0Rlx/Ms9sZMOqludwXR+GTJ/XimDGEN/n8G4xgaTI
SzyviZ6wKNgkZ5dJEseSOQ5SEGXYr776jh8TdhxJsZlfHA8PNSLmC7HSekf+Ww2Pv8lRw1UBkMVn
sSKU6Q822Rb+0H/P4Uw5MsHdb6896PaB5nUGapHT8jVHjesNk2Q7sKqigJkYQEXs7sOBVpVK4EQD
tyL08caMgYk0PQdlo8l++haqL9Bu15MSk/2ohtmxMNW6UNGCPId1UnzDPPwAgav6lRbtCnY5udpR
DyO4skJ7g9US0wcnfCh2K7Udpi6pa1eHpeTec4P6sIZtHpeKwaPaszTeII4qliUAcLUNNrcJlE94
IjMStK1sgLQHc4F4xL9+OkCwsSQ4x0c9v66CcDxJL5S94O/DeqxSvMoEwfkE5BWRkqpRNAM3Tgwg
yP+pk1cH5EVCKV+Myrj7O/9G8YdQ2z6ECP1LIhwHhYteZuFYm+0hQMlHI5idBuGso4ceGsmnhaa3
ADVYxfKAgaL+BJdlw7LbF3eYw5Now2NE9nLiWVWW+RaCj2dYt7g155ru3w3+c01uI/58v98U9aEx
UvhVxhbuWMYeMN39vFzwQZgZeYGzE16EeUl4WSIvohpTXpdNPZO0qTYvzNtB1OCwaYlnP2AeCimu
emxPrX3wkGn85hhowlmLN4q60Cvk/AsOwBIfjKvxYBsIFh8uSDXrfEGETEsBVKpEDaf95qOtJsm7
jhpQM4OVazsTrO/f1BfeQ8BDUK1hObztFQnJ3yOvPRJGgj6V832rcSytC4VxS3AWuXId257SXZqg
hbUg03dtLLJTJVKYTpt99pvAim1aeaa5HLe45HSv5a0D4g/ovbIfCeklHm3nPDBnJTatvifIdLbb
twIYDRd6eyoIEbIRV2ROffgIj0vrOtREx3GmWhf7qdEb2a8kw6kS497C4GUprxcQTvw+53Bxz1g6
3+cI8sLPbCgLNYRhJXnd9MtHvydD4RH5VGsbD48gRVHxBguKx/G87esbyqMvEC2rbfKvIuxSm1xP
3QfIOVhf82DiMLvJvTUf1lfgCgIs3SzaTkPT6dXVLZK/0QAgCRb523r6aE0/RBIbRMy0LTQCotcN
SaUjaBtNetZflVorniDPbvH0ZKylVZ+sYMeFmg54KwOZi29RoO9TMHidu1rJqDTUDWX5CURBuofj
x579s4nfn3lDxEJtl/kzi3xnOD2D2aQ7HfFSU8Ky6iWupFEWPvAx5pRu/2+9PS7Fq2qSqclVUaqE
yWm9wgF6h4iVIKfPvQWYfIArbczoYOGqBNL1mKg1E1cG08ECgOR6ryXTHKSoU/RL74X2fsnz21Ao
vxtICRC21geRwx4Z2ywh9FEvUPg5d4ISdAzrihlm73oeLBHQBJzOJzFu4uNbbquMto/lEiCp4w+o
IKqpE5hE5MO6jqIz0Oh47cXmZw2a4+QkjrhZ/TpRdLM/betpTUA4Jqnfn+0oHAZdRq260wRBx6vp
omvWdfeQPPchCp0GzdrcN50130fUpwqAEAzs4YLWN3pR80WXZiNGaTnshQOeRDHIK3f1fpnaGJCC
IjuP2WVvPryzMf+gQc2tTpCnkQBvgl/9i3ufAOhDkVeX/ep7EgSkeTptCUT+jj/ujOpIKWGFhpF5
gcamXNlmKXNrfJLjqFkKrS+vkvqD/XAlVKi7j1wyiBskPvUa07SRfhcul64hHS1ljoq2ovYd4Lxh
o3u9wr1LEg+d4WuJ8qc7qZzEjm4epLlASpCxBTPWrr88K4Sgs8l8cWQJ0KdYhLYAXASGYfvfbAiA
NxCCgHjSNfRJjb2ZUqI0qULix3dqJBSwuJ67Y5iI/wVVx8mV9/fjFOTntKTNoLzcOiK6WWyIHije
zN2HXI02ZdUqestKa6k4IgA/bXs3FQ2zKBvSj6k7MP81BkV0Xe9yGwh20POFAsppn7Hl/Htwf1xH
r8+srF09aU9FeHzp9ckJX+x1tnpkMG3Z1QZ7K98xRLA75ddcnaMTeyfMJ8gaxXsRPSvTFRhmC3ZE
xxE4L+S7eMVO6QKRvYZrGkYSc6CStrYd0+lwGDWcVTROi2o6jgWuchq0k5jf9OvuRmCUIUafxE8Z
iegiIwFuPBp/76tq0pl840aE6xNEUx1JdOhbIGu7ks9Sk5YXGUMcyZQdnLRZ2uF1AKblOsnAMWt4
cbJd8BxMfswMwwB3AoWnw+sf72/Ad6Tvtt+3urzyPl8JuEIScAGItve1nk3yuVG9D3oxeCaYwhu+
CLQZ13I1LgXpX3UOzsDw1b0c8MLy+Lwa3cVQMOo2kGcmeQkiKboAp32FLCUZBO3o+u4FJ8lKjVYB
vyeoRH+okus6CpG0gaxvgLYKoRRoWNzP3ap4i1nfv5GujGNJnNvjM8T8GHhKs9QZCwLrqpua2hDZ
E6cDdk8ti+Oj6iaAo8smRypBiX5NngtsFnEJTicayarJWV1C703XIwP/+j2K8YQQ/J/tUqXuiXY2
9ykSKua1FriXM21/vun+SiG3xLO+FVLavUq986XyUUMXQKxRH6KHUnBUKiEULVcg73O82NDS6Yvr
bI81dIFBzZtP1epQlGQNcplZlKUX3BgU0ANcIJvo1OOjlB1F3SL9Dd8EIkiaYkkP5EEdDfWhdr4P
Gc9OQ+jyUAh0gRxvJOI95l+JyL8xtfhJezW/DoK6RzUx3gepfh3LXhA74xbA+p2P2naYybWZKwzh
QiMt1xG0c6zzOlNH7CaKtqcSQ2AtVoWemlqiDjCYTROvf+tAQiTW61FzrfdYmeWRDc5c7DNoy/fs
/C2YVqqFKg1dQwCFSv+XgKR8sWVrf0k3H/WnKC/iighi3ZYq+n6WSfp90Uaq7Gu2Mbkz/M7lKu7C
lNxSNrVPfk9PUFFhocDgGfdp8HHoRzd4/RvGC6/yedO+1Bl9KgCCL5ZR7d1uyGcvlZDMVAWcyKYX
ASKhqWhD8wCDyutTA9+MG40vWupGQQ/etPcwomhlrXQ7dH//l2Bx7nljuPvlqQfJOS+dc89BFPlE
YqB7gOjPyi9/72ARAJrZGI2HmW7PhV+lJQk6Pyu+GIB4cd5DftClmL9edQNAfo7aTY4rmH6cMnQk
J9HWmdVxRH8OPf1ytelDLpJe5/ATtFj2jq1JDHVmxT0T+m0yqmzynXahsV2hn7BkENGegdH5HR6j
TPBs9z+9Nu6cfCTzbXMpoBzySBEZimIVnj0+USG9PCIe2AKDj/YGizMQ1QUqVp0lvyCJyO8Gc8/x
LcDcLC0DZIO/pWDoiMKWlxIDHkRygf2vtAw+YXglyww5dwgDfs7u11M7uXWRYIWlZRlg+f/xQFJA
/QeEpfKwSld+tu/RjPP5fvwYq5wFnvg2Zudf2QKWa58PGz3QiUeyYR5C5+MN7UT6pMOtf8LbAsWx
+lSWHYn7QHDfDaE8AvWhAEwv0wvZhd9dJfGitEefBvriICXO/fqLe3iKHZcCmegvHzQ77eje06OO
ZRnw6kfw10058mFLulGoRUp72rqB2pGk0YkIHSFBh2L1NBfsOk68bo0MvQp1LEgxbKXF82QRH6iL
gSBk8mM7ofTDuM1s6/da96kAFUo/LU8gY7RxzWMXwxKi1GAiGfIwRz5/W/uu5ZFFZnokvgRlGNgu
xZZfmzTslNCe9TpDleOQ3wmAjfOXlBNo82Ow4mfRe/V1mjdryOqLZsZGk7gsDwSgauYQxo7o2xgY
n6NT9037H18TiVmwVpJsort9APSkbnl8X3VcOlxEsY+I7MJ1JBvL60eEY1rEdTnxTn1YF2m5ppZq
TyXNePAcI/gu/WQefW7xHiC2pW3gCNQlaE2LwS652rpQH5xrqciM3IDneOiV5mApwVNbSuiE2nb3
HdOxS+yDuzP2hyDRd6XBoDotcHsdlCqof+3rQyiDUkabsAnPo2BpfJUevnEEdrjcLBlTqh3wne1l
Jl+Pk3n8eoLeyTfkrvxBTSamsm1UUQO7hKfO7bd3+VP7livobrUuemOL7pWIHTD82GRIyxnBTPq0
yKO5NnqAwQveTylgcRhAdFaVpumlMDiPqog5QaqUa+C2XsRLN/CZFCRJd+RA89QdLqUifG66wuCW
fn2Rmt+PuuSP9dNVFaYeuiOWb8blxH5Bd6ezwuZlyR4RQ51/mp7R9PT+RPs3fKvn3YJ9OrmMZJdd
mi6mBd5XoNheQ32dSMdMqp/3ScI6G626XkrEbDSyIs+qV5UcFHv/BLk9uxEX2dRG3P0w6AnfZpdZ
9mTv25lCDSpac0HgIvP5S0zjTYwB0qPuj/2OLby4FpBiol2hEFqpdSKc2fdQMn15ssRVqG2HkAGt
uVWoXeKsOtoOshem4mcjaq27namjWOxGA1/ycnK6IQo2wy4/AjVRXwQ+G5vHgPvofpJCllHeLwMP
6lMcuFmK4KS7LsNCuHTzWemWD8wI9Eu0hWK5MvvOlC7VUE7jDQzjgXZePYBMmxS0nwXATMYlDWFk
3Js3+4Brmtmp2Na7lzWLo6/MZaS9TfdcJklB2NI+3SqG03WcBS6ONpkBumM8Bc9RbFjRGmVXLAi2
uTFFY4cctenOxHC8VO0rJKzV7i+mFIdeXOJtuFgL15wEhHTT2X8as1bGwkw99yT10smfBpFmQ8+8
ItrD0SEEQM8DS+oi34pXYmVm0gkEk0cv9FtRR+m8GGRRiSFYP49clUDnY4PCJqJQatx7p8U3dzFD
WUBdcfqYz+gWSbvfB+Aqw9svCU6Kgqgj7ioQktgKtnxpJzCQ06dtJ6mP1cDgCnJqtSAA6yRFOc5f
/ogP75s4MFMZhe1nPxTziL3RA7cbVNEmgABnwnIROYKGH3F9AP25/Ssr0MKQbOakN1jb/+NGAIjB
MnoP2ZdvwetkCbmCXPBKCRVlv+qW3BN9cYlpVBzy7llVANoALx65ij3QaN+A2XQV6TVuTVpH6K+B
0sQABjKEuFtBrqyxVPEV5grWCRnOPQAN+5i7TQX+T4klRtRBT7NsoUUlShuu0QAaqI+1KFwkS2po
1qWJ5m1YtpBTloLev5Szw1VXr3Qi9WqSSDDjoEq3vlZdBBOyyfqZmwwKbFumyi/ZxiDgQ6oi+wCx
RfyoekGR7rgBdh9I2FEQVjyFqvAZDNucSrU2Ng6OMKwQtrNpUDYxq/ujYQGHX+U+rOc9D0dYrIbo
9JymMWG7GPwrvRTdCKMHXN6r4qhzNLW6hMDZT4F8hvjIMK4G025TnwbgEbqQxHOkR9tMVx3NASv0
2SKz8UTNoTepl/4najyykNgFe1g0rucNX5c38dCHIjd0FkmXMweETjiKUEiLJlVSBuxAXGU6mi2z
U+1ATIY4Ci7UzaeqzHQtlbnrZdR4crn5tJdHQtcUY8gcJOwgicysSqoZEnudKPuoBQTJuegsAlMb
k82kB7NDtocGA7kz3JJEyaza1iLHKO6uDOD5gFOeflv8f3YMWkjQGY+CpAjOaLcSF7CZ4JiF8hNS
q1j0LwzwBgByuf7eIdhQWMRU0v5WcHRqNtvlE5RQN1gKSqPzdNiP0Rz843tigdYHTJGmxM/AdyM3
oIYi103dnSOel9NT7wQ0Af4BsGU2QlMU3/lhSprLbb8o+WujYxuX6mfkJuFbd6tPg2NfT/VDGswg
syanCnPomDQr2ykJ5VVb0TzI/QbVfeZ27VELxVfL0NnjGZqgTrL1IFIZU6Z4IdA7FPBwDyxMt88Y
8d52y+GTjZLLpqTCBoP9LADT9gKYYJVrFIevt+K+BOUPOIwboNeFzp7hMWTUyykNLfHCM2rI93WP
8WRHMRS+m2A5RG0tb9PdJZ4QlwZyWIMKBle1c/VYODG+IxSF2qjr0kV3SucmvTVi2ilHc2OZYgAI
c+CkVvD4DzDerMMUKFZAJZ2aqjL5WV0fmieDNlOI1j12yZN2r0tQItv75ZdgrzllOkiWQILr94ir
XIzLy4NoJqGbqqgRhb4UOwR8zKhzgj9d+wu5fd46IZlfgeE0NweapaBy1/SdhI83+T/8QuWgs2bb
8ap4YwgdTJd7w0EvdXM7SYxZ5hWKRErlOAmjH8Ah0v4bMSGTwQ+OISffbED7EW5n1zdxHpNZaE0t
xg3JAeudbDWoS01kviiwIAoTJGi9+TjvzLO3ujnPEEzXrqq+0qG+d/5V01KJi70CCGAU2reXv0+P
QgAXhhU6pCSmU0Sa8UldGGSq3YCFbLwdKMMYFcD4Gd0H0nt1mAEAk6kpyAAaZVrXJeeVp6QkAzuR
v9vnxDb5aSUj/CgR53OAlI99HjlCC/0JjY/dzjvYG+9xFpaUvs6cmUOxbPc2vCLkT7BYMeHt3Efj
CxHfjA26QJf4JIM6nXMmgAaRHUnwDHjITrhS3wBgLLSPHZ8bNPYB3e2UbrhNNGt0JekD3zZnf2E4
V5FrRIUx/WfeK64/doEkllxazcRgGgmYfiUruNwhX868IgEi8UfbOfX9jaWHCSC2AseF8RNmFvam
DgMeNsjtKTEjjFOFy4mJ687n5mktCH3AwiTg9NhvyLwuze3m4O6SM7BGXxEM1/djMM6T4+6BB9d5
+nRAXrclF+0cJe56QY1zbn/nRM6WmULdhSHe8YrlSIJjZZZKxy/NB3StQLK1shGjIep0XSBzPG/d
pEEVl18yqK5+BUjl+JuE8qyfOd0XArdPk72UngDPMl2BXiKrfDrFSwwES6z7fPYi5UvqHm9Jyjxd
IwoGf4aqdIsUSqQV3AXJJG1wBOydqxvVJOs9LB3MDwPzSGS+VPmsUCNwcQyUI2M2gZJrxK5PnHD5
80vZkkzi434W3fVLLde3vWP9W6ujQQAzquNBqffFjrY7fJwAiProKANu6EfMAeAR5sE9XQhYEREE
HT/EFF5Yhd6tYZxFIMrdJGrcwxjQHrgy5RzJ+Wpcc3dNFJXZpFqgOjp1rExSqyxnz7HRi5/KQGze
lSSYAcNXYVENw9HqlQ6mT1+hMWHLXVtYrapfcLFhnqQdhoNd1gtbO6z8BFF2WAJuLEKImIalxdoU
mgKz6EAEBJgxQIa/82kw/FrdleKq9/kqxWznd4s0JCBVpT9tkMNLdYqWhRgWiQRUZrDb0zGwdVxs
sMrAnCN5V8ArWR8eEf01NWan8wcRPF3SlUvdBmintPb/4BDgNuVRUXVuj8wkwB+ylF3WvoVRXu5g
6zonXgHvnXqMlwgO9A79IKZD77OFk8X51SQSTxW3ZRxrMidACMEv5KupLRLvLylrDI8U5o34Nqkp
uNFj0wpmeVPfankfJc1zMMiR23Nbskthzpw+i/TcQIVLbzs9Z5ZjqluJyWUFjvg5cXEzF6XmEQrV
Ar+Jm/ZWh6V3McIMt6H0WTVhwvpz0l5Rj5uvXzMkcxTO+/RyT4V78GQ2dM5MnhmeuI/Uclj9PsPD
5WLXwB31DfDi/Y5RY0g4TcS0kg2JMOKXrkKA1trjj/AqU6XMjOl6IRNLvjY+keV5fRnnz1YXs1RS
uSXdGqksrXAo3zT474wBx5UepsCUOQLQsrSdYPEWma/y93Enn75KIWRgyYQib2Ua3LMXqQR56c4D
ZbXCPP4qlpmNgFpwlmLLQP7HH18xI+vFGqKJH/jx9F7pY2208vFEEpEZYEgSQ8pLnAEH8RjgfYRD
cz7Jo0q9hQEPIkr1ulAKZL1NtnM4LyqxrC8aGqDGLToafD+MLDIxylUgYSAVRYRrIhfg2CdaPOMb
IsduOjXwaRDl/l9Lk/aMSH536gSTiojgxWyjq6UHOu88UJTwV0FMJxcPb7uMobEY599kFhBBbfwI
6DOUJGbCvOeGDT4i+77A0VdhkxyFYhFTnrYCNqC5O3T+Z7B9hwGY+VO6GBlLcfud4GXwXYqm5Wg+
OTl6aaiaMynHBOZk3/ztDtB080vxej0JUc4rR2LPVKSbrjHCa92uEitbjnu2v6KamnqDt2Yo+eHp
6rJvKGk3oTHnWYrJc8VMPDLjottFnjcEB+aprNRI7JtKbDsEEm9vpILwrKwTf+uf29XNSWabU0l8
vyRM4SQD4X1tD2An0O4QDxSq+/WVUWVfx5SKnOUtaJWNDF4eZ/7gq3b6TIJiIPgryef8dpGnjtUj
rQ5u/0V9qzm6vh5FOEqmffbSL/QQOFdeTqvfgu1ZU4lQMARckvH8ihqB+90aOEU/Hd+/S8cWEskM
nc3Nb7J9AfClnKDsFiC5Re4qCSyDDNXUyLqjDITsWyMvJsHPaO0acpMzoRy0RI5J/maL9i2Q2cKi
JSmM4YOPd/VnbDrB4evQV7uk71LrhGXuc088FHTO3AHhvHHNHmmoo1/FF2bGGkrL/tN2cIAN8BbK
/stTaSboOOV+QKcaFvWDVHeRBDKF0cLpR6PRlPEAxB7PK8mDZOAmNhPGskkKF00gO8HFYpQ9YpZv
GryXMcYwuapfqiJVZKsLKd38F+8H0QIfye2OyWoL890iVRMXDeMDOwsueuLdukr9AOBcaRbFWJ6y
dpbvqVPiDwvuP6UW+UFAv9PbRgsZ9RpA+1kmZOOxsV1xOWlJSdcNa2erIi0+GRAqca3u5gOaU9a0
34v6SEwtS+FVtqZfV+Tbp2bIGa6JyOWwI+HQEWZmurTjxWDW/E0yhAayD1XzLxkDCetHI4SZtDGL
1R+YT1NVRR2+/AC3IC6hSrXaH5vbhRuyx5kgGzVa4VR9JB17pFosh1inkruyc7mDOkgDzT9/6RUd
FPcDQJ/XnYatqt7QNmLf3FqQQhciywbBvc1Z5WTazluT06zBPviRGqRjJ03NJK8gmciaVCFZoi9K
+hxCGLT308TrMmfSci6lub+OPg+9XE38V7anzZyaAxeP84GAzm8ZnO1u5fc9i+Rc13MY4ZkpWoix
FDa6f9R8s3q5EoPbMfwsvekjli7hC8sRqKxHXHDLPr9oz1+Rtlafe9ztcDY9VSeXNeU0E615QBcm
Fim3U9duVo/Lr+Xqc/i9t+ngt3dPUYUGIT+f38OUHENjd3/v3uorWukhI0FKe4+GJ0lTCRR0Rs2J
Ty3oM9mBmjyI0QWAzQ0Vk3Ek6/SZ8wUKvzZqTDpS0daFp9xyexP9NDzDmzdWRR64Kqzh/UCKhBlM
/YWWZbAc8bkCPl+6ww8ac6VGYJoFABZIqVNHII6iPw/HwlpNMpOqw7LuOK2qQ+OF/oc99+kFYouh
mIZGC3NH8DerESo0KYG7PymrGOsjRfejFj2ic9NB9rakLWKdneNojrZziyU3gDNZokMq3n1WWnKU
FJ416RMqG0DrF+LTOqFGZC2jV59G0jchVu8G3vK9zUA8HmaBuHabKWGXymWAOBbV9/UnZB4CmpRM
9kEnslSZtNOsYh4ejjoT5L5GWU/Q5BjrX5WQ/8fvpTZN6Mbcjp0js8fdu8Ef7qTBn9EVHioTRNLR
fzhfBJMfLK5qmWz/VKViMah4+K0S37cCOB/o/lVvc4giLge7zcOl9k3wJkjMppoPGbfJq0o+gCPU
wR9mgjSKyL1ve/hKRP06OGcF7IADTPTUWeKp2XHdXFSGmYW04WTiTZ+QLQXftRZ9BAuzW7i5XmoV
hsAHuXMJBBVXvDhP4OhyR1Y6U5SvtzHu0+yyeKIYJWK+BZ0wYgdTSq2gJ2N6RAAIr3G3fzTmmibF
3p5MFgUAGD7hoXA5MF1X2NTC4uB+QhCv82VQnC9etJ+GnWkrtIp/yF3pcI7qycJ8Wc0ANFWsjy19
SVPam3ptOS0opBlv7fgEwMdVDFPiYsIV5kGEnBjojeIT7jrAgFvj8k0Ijt4nOHjm4EfxkOxPrOip
GUdxvHrcbsFYP42vHXZdKh45hOhF9Gy5Pk4WL17EDhYA8fHduTBQfX2FqFO525my8MDaTBW/44Yj
w7vm960oL+GAMyF6rgOavHEY9neV4yH85pJT4TNQIaLPwNzqbA+WANk6s4quEg0dcN1149pzblPU
GC7S8QSyibdBIOiZYGR5cO3+tEC/M2UnG3sMBpx4+1/3oYKAGUMA8PnkNRJFjnramqxaC1AZqvQs
RjbnqNHylkzP2N0x0sbx4j0oNNOXDopGZnJ2PSIBD7la2kuTldqyEHXp+YUtv/eGjVCGQNMSwmJV
m/AjlhXMEuNKkFmBDFNkurQsd9+ijIDDObR40iEFTe0CIWAKfsRRzn2vmJteS4+RzKRXBiju9tLb
MU5c1WYCBHm90Die2e6fVPRs0tGBidt91Je3fafhpnrj8qzx9cwwB73tjCTLae/WPZt+8KC9rCyD
POT52BmAuoBB62kXIEl2NT6TOFv2Uf8g/TZPCXAvsW+pBAZikSGLOXM6N4N1Oe8bhVM5VQvlAYNV
EOPz2nQIL5qHZG76SkB9YphuD4TOLHtKmIkE+ntURlTlpkk2oa679LJX2PPSuwO2N5J2JGXGZ0vj
lnFzaMjX6oOjR4HAz+X0EfAZhEBhUjZc0TqxLYxR77Wxy7X66zS4e6wtxk8oUSkWzVTY1DtswV+m
JKLe8mDupQoJF23bjWMVvullGW+FYP8IS/UZ9QwNvlfPj8AVzwY6YUi1hXu1bzvVN4rkmQ1d4h/J
m7z7FsI/m57iMugyGQu7Z5aD/c9bDuHmidBC0EUGZRqJeOxeEULH0DQM7uNtQe+Pf4iylYjeBEEy
MEwyg4ZRrkpQldX8NW8gSu5tMScfFb82fRWawIlmzG4z0Ewz6FcqVqP7/6wqs8N+GA9oTsuLXtrX
xE9vXwWrW9N7IsSE8jgja+qP3WdmD0AWTSAMrx7td919pzz/SPh297yjFhO21Da5NHcIdaccKo1i
9tsm2hCj3o+3fzMB7odD0J+TUmMof5JngAjKCfcQfHKWZ3Dr1REPUxMi/0Cn5Ozmq46dloOxExty
/WZsUPOMLR0xkjCeFgHJd6U4J2tf76Z3EnRnbuEziD+LRItGJq8HrTUXX/F2Dp678EXvbfm++m8+
ITjHkga1fZirs0OSclWzWi/jaEpJJ6G1GwR3ykPhCSWrCc6YhmufXXXy2YjSbAEo4UKqNNsLSK2p
KX79XDr3/6/ZAdnrmJHIyVbJ1hpH+00a7Ay0vgEfQ6bdLPUW4K+ioTL0a/ZkVaglpWVYFnC82MrK
XYq90r058Bk14JvyABNJViLFfWhRH2ksmLMY13dVxtmIhXuiIKnMFWqVZaHhp0qN2E6hnHr+xcvu
/iiycE7FZlNUAaxphYpaanRe6fq4CY7fiO6OenLuT8pmsNgiyIKx64F4SI4lC0de+YoV/T7LezUn
9fz8OiOLfBeaVg/AjuVqhRbTbu4tx/01GNeUS4MrTWNFRUPN0Q7EXgh0dee0lToj2P0zd1azFX8+
HqDFB21ppysSF0oaFXRkg1yqpjAyHjmuQ69fRdgIAU8CY2IJ/0LxCOkprXzgNMzQgh2LdcnypRk0
Nk6ximHRhFzMKM18zcMceZ/iJCOeDYObD9ap0PorcWkqNUgUKIH5VTYTCIzDF1G6UPIRZU6NX6cz
b4UcauzUHQmW3G/F8j17kENQjHM2ARwzFUQwKAkE87Jtx1QMHR5ponF85yixlAgwxIxtGWQasyUy
rVH4SA+q1QkxlFF88Gxx6EOjMZZzycUPvx4TuCh3AQs/2cVpYz0HVFDbwwN9wzyKK6PrJ91iaACw
EuwooZvP00wM8L/SQbD9AfVC8aFARNPpLVnsonUgRa4eP50yZOxfpyLnngUEt/ZL6bQGnHrrqwVU
Tj58hjb6ZrW/ycqVslk5HE9dKfhlGRhV6EBbBtpLV32By5mi5K3n7J3bOg/wpaewZe/JrljyG8rI
Vh5VaDwqcllSXf3mwipGn8KZUsm8CM9U+vu9PNYdjCsaFMJAzp1ZbT+1zwDMaX5hTbCeNAnHdsuZ
SsE4Vt933M8t2EopP5jL9LuvFD/vyeSEyzkNvLMGafqQCralFh4erOmma3N7Ns5OfWhn/JUs5GO/
PSipAOCFrgqTra+olKCbSIY1mr1Kb36emeaUJs1r47jMKlozj6INSJT29Riec+mHRboCDxaF7C9u
KQ1KbEGm+kihRt1pieW0vWaYCXjc6tNS+HrDU/iEsnElkGNO63gB4MEeZwih554midDv8V+dZufZ
y2ph3a46jkyMSNrckVFAbxHWM+mwlSxAHzfryprWAayK9Rm4lGJuQlZ4pKXVOH7tRol4nST1rILd
KOA0Y3mkWrCuho3/qCwaPV4ZZHS1x856ersWvOjGHJaNUHnz8LM647+uQsvx7emOEHhbkKx2ra9W
UsgEQunxZDKyjsQG+3TlEMIXpDpDOkstFFGLrFWudORfobbKanLcyfra5hcPMJzRe3g8Uogo3Cjq
Hy5jtnUZOD62gZ9SEY4vFG7L8XNIgLzqBedlKPTznESvw+tmy3hjpGYKCd7JCsxQuZxdHC3JDN5k
qI6+c3ddVLYbfmTlev0Laxd9lQrQya6eN+ywqJ6EkiZV2sKJP8icCx6Tz9mJZxodQF0oF0TKgjSP
QYXF7kUd3jp6ydPkq0k1CT1GqRS+Rx7ToptYaUrCZendWUjp30uZ7w7nfANKLsgPWZ+UScMH60qR
Kb+4qh1/uvk/mv/6pu9O6mKkVhmncK9qYtNexUUaydjuJiTOVlVp5J+bUCCT6aEVu6Tn4yoUWKFI
KZ8ZXDViMZoC6ZiFz8BDXro8wkJhqcQtVIAx6OnAWAL2mCG36NwKzjeqKeSVLDrHxaf11d1UdlJe
PGs2jh//GakDpjWwl7u9QJGgHwslrHP4pmNhsOgxBaiOxt1WUDD6+gLZJBOrs0eZ3ulkz22vlcCC
SqDanjNkqXWQCT6YCCrWHkiFIi7YMdDOy7atvroNSb2a1P0QzcRmf5B3RbrFIc0+lbSMFlyM1w3z
ZSd9PZ8hbaslztwc3QosBlzWfVhVozaeuW10HYrGYomDy5FZGisw+x89VfcGdC7bVAipNpyEcVgY
fTSQMBe2rSy+ke/Td++RA5wiNmfq6XcSZUf1M3tepHdw8KZi2IErPY3n8yL/g5f1nN29041IN/4p
fXQsgCTwkO2mGkX7H0RW1saR/HLBZ7ujc8p89KR08bxsZ1z4DcZpd1Em0THh3ilF5D8P8iC2KP1F
QaKtU8AsrovVx2sNRs30T0DnjHsYiaT/mPX4cr6rRBu5oTd54gVMRvKpsuD3R7PRY2CRdNveFS6B
QU3ol7VORbc826DUTK709p2esnQ2xndffCvMk8QQr6090nS5q7kHUjqdf48mTKwaJnf7krQwA+EU
NFR3HeV9LRySEy1o4aXgDuzTqs2lWpbzMLSqreLO1CB76Tzhha/Z9kb+zIhgZPUo6b3X12ksllzW
MCili214hPiI8hFYU2vCmprR5sZC1G4w53egrtu2l0RIrbqgrVBiPgVir3rM6JGJdcMxbAqlffjc
KIIBwQ0KVctohgog2vrFjyrT9ivNYHOcJnLsHRrOJE/VraQLW7qdW8IxaNJjkqNDYhdI+SV7JD03
NfIuKcnub7kvoiATUFQzvzGY030//0CbQMuPC9lOEAD0yvah/nTtL3q1OMJ8prTnOwH+Gs4Wjj61
OlBe1c3tArBYQQ51crNHiZrLVIXiQ/vfeosuwVIikYwGSuc0xMfzJC/5TQsvymmbj2bp6is55bwa
DHTQhlPpnjT6yOq7s3x+ulBDwiA7Q8DuJhyhpL2n3cYIWINASw/2K+hVINeuRFopSFxFI2OkF0sO
nU9ZID4aAu2Wh4aXIG+z0fzRbZvXywrs7y31USNs/msHY/5+OMQB72KKR3LfoXBHQCMIgiwXX7Ku
0u3z/mRd9Mvk6kO7yjTr+I1NNLWqT6z4+hMJI4Rc2MDo/FzxvCQ+SyBGmeEvUM/1aa2EEgfWDX5S
d1iS0utGvBQA+fr+yb+hmLp2oqOC8v6loUkuir9ard1PbTP5d+Hg8bq4lcdHh7JUEnNzOGl0p1j2
d5HM+FdecTHup+anajTKbjS2drseROXIajQXUkgUKmsuN+HaUw5EinPGXTsTtzgtcjPzyKvV/ki9
g9m+Z9euHOwuu1anuYov0yWpeeKKQsBAg7ToE5xOREjWfrTGzwdnhY5Jkwu8HJ03MhTKxuYtQSJ6
ZqvJuuKZQ/1ayf+ppnYyYQAZu8KdabJXU3cWFQ6s7vt7dDdlw35xr0d3SsF+JEDsYN6+NU/z6LVQ
LxsoKhXSIy8+aCaBmFmnKysrKoPXuYyv8wfp9/JFxSr0S4xAAqRtQusoEJAwDm6dp3+lYHxnIT4Y
6GgzsPPabtpkHAy42Lb4C+whZf52kkUrZqbd/G5qXvNoLic0FLk6nsp2HzTR90PtocuRLpxPu9CI
KtPMAeStlEwjza+ST9er223wajicxx1IEX9a+/mtXtYbEh1iuXRhM4x8cApB0HKZFE5I9DXgyRxJ
2889OFu+xl3IhjneMns01HPqSl0X9J26hI1CMkhiPf+F+dmUix/+BMeB0J96oidDKSnMdIvX2SF0
NDcFwCwPG2hKtVprMkeNO6p3ucPDVKspnPnUQklltylz4fQwWSXifycNmMh5oAxI9/fr7pD11X6K
vaBhj2bfvVJmCcgpAvYvnjjg8ZIUQkf3StXtHzi4A1mbwG10hUMHaXwJnd7MyCh9dSoKYpIbhvw/
XHqGex86RtMHSfvsyM7LHpuj+2RodQ9DEZHYILJHHwH7NIrwqAc+sCMBqStwk1cNKDyXzB7l7iak
Qm98upAPnLjlcINUGVpTyzcRH6T9X7OMjdnFPyO0oAhA9LwBtW5lDlKBHOYC+uF+4bu0Z4g5bjz5
vAByW8GVcn5gLIx/4Ewa8bjulX/pxMajtTkKQ7Hi/V3mxMMSZKHcbGAM66wGGzZdtlyFfpr0XPab
V9YuxsmWhO9mDdx9WLUu5r5gnr03I4YDHVqPFnWR+aJZ8xruGbvY+sDZyylwst7tOCl1dGk+zSJ0
bXzzXfe0Nw8ndwDarjqgVgn0A8fYVSS0wkjPVqBHk+N6Zf3rM1WqWb+L3uLgLtdZYqwISYPnlWt7
aschZFl1LjNWv9/YqWt17p0DF5Hpm3w3O3JSev4Pcko6aSaI5GLLFIrFKwAAFL3kpNjL6RpVu0ct
ktBNLAmVFPkdsPIu76BViHbbtSdUkOifmaaowVWuh4bd/OO2pRK4TL219sGN7pwyE9ri4KKfivvm
sEv0TLzEOKudv5tCSTTh8z8TKjkA+6ddGkbB9lzzrypz8HKo4KajPCssMQXvIebLz1vKFHdyR1P7
xC15rfuWdEZpXk7xSgdzsOzxA76Dl5uL9EFp9TmLccLkwvkJ75pafRdVYxI6v8bYsk0ZUqERWPt5
teYUwoa382wItKHEmbMMXw7NBR/Dawh4FnQ7oPl9vYhee8+H3EFjHZzOcLhiVSCXRO/UqY11qqKf
qWoBZSQ2ET+x+h+gk4w0f7ZAgHZ/onJeH065STwtaK3GIBfjXJo92Ax1+4rJDpfQvdvUlCWGuwkr
/j85noFqpdxm0pQFBBlEA33E+DuqCskE3B1+M7FNB5CwHlVm4XilZ5GUa43dLbkfB6fixZFv8CxE
8d15x4U++VzgI8l3DpH+fNcm1JFyuKDggEcjOMdLzJII7uovaxuop8N06tSFzrDaLbSlFjHvGQOT
MZg5MSVVF1erxspwOjN+8RPv5hPHKuIS/yn7OpSDSrcUBLn+8OmWc30qLxn6nOn33HKZ9czavNfN
yet4SHchL6lkjXg8OmnMA/M8gb94S+Os+Fg+UPuqEEtO8FFGbvp/Ig6mf5Xw2M9nc2cdceBvAUMu
KUEZvpznK4tLbN4P9L34m3rmD6Lebrr1xifHBx9+GGrIGqYGscoBicfhqsD6f4Uu7qUgaL8t23d/
7OKnjU6mV5CyLrvG6hcq5DlmxP8tNILXz1xNssMlbra5WzVoN+6ctUALeUsCGSrJf0DB29RhQV8y
ckHHyqxfNKCF9esVn6NSXi/oQRH1nr6wxC7P25v70SCLAvw74hKgpwpRT+s6gVmpe6/eEvfZeFSu
nt6ljeJsTV3nF9ynt49tTSsVvELmUYoARDwL1UxotNKDVfTojqMqUX++WSI3T59ksVrFolNlLfcb
T6K6rlAcQuoJRN3QkZGVARt+lIOM/XOHlf1BlS++GIIZYv1cfD/+2x95dn+VsznSHIgRXiSqIDJV
hnbjtT9pQzpaWhSCM1A/KiK2MTaEzRXZ6quVfiLtNXmkudJF41c5HYXEQ/9ubmgVBDO9x3le5T85
RWUJOhK/rEc5QEk5sU9h1cYyh2NQIWj1mqurmKvfvnu6M29RKW80ahAVvzBK0/BGmWqKHz8E5a2C
dvCwz5Sb8svtVz25y+UF4FdrYCwsaJXgoXPw8zIyz/LORjb//o83r6y8lzJDVPwDXcmaBj0NkeiG
oYprHoxEPzGW5F2pNnWWcmsH4D4En/1Qrcob2IV6TKQCh15tIvqlf//MMrJTKnt4pf4xuTsrtv+M
/UYCbJOt/GuVWRnniVUtoUSwM3BZ6LnTBkZE/bZeEzuwfiLtQ/tH6aOcwrHdx+Mk24u6W5nIMtAy
8xPmDcKZ1fbSBKuDQR94BVbejubj7/59f21GfdUQvdg0ldHwzaof/rB2mfWhgmbH4GSCWXselrhf
TJbV9QJ3x6qOqC+HivcVOQQorJ1UqO9zGovCzBQyYP5Uc1lwBhVSbT7JVReJfSj4iE02TocXv0Ku
4dM7WgygrsL3YQVigBbBDlLP0x5vpMP0qV2CJc2qwUTLq6AtmH8yMANyLs7IC8KCJ+jrpVTtfOD+
evYdPc0inkq35zp1w9CCo184KOimbxMkkLtQbUI1i1nLNUQgosiZfRkip2Y+4AZjLzzZq/DfqJXb
TWAhVUjhLwuZ5qxQX4cS1mIlYtRLcRv8fHz9+7bP60XIQAuxvsFdzb2gYVEzFR0vJQEndvtOlCag
L41a2WmXFr+oXgnLcmk0hyqpVdOJ1akcu728r8SYFBSFW0z03JqO7Qv6USuS2V4qtOfHfxzSoIzn
khmk8cSAukdwuYzomsHPlHdiqBL9sxDPP1AoKzYDF3E14CSFIabKvKYTOwwsN0TWv0/jkqZ/ue3I
4EFHOkEb8iZYI/VbI6okvoB2v0RzSINmP+g58TrNJlaUG/G4EaQykYaJa83OjAsksmwhbIgs1kjD
URKilNtJPv0YiTsYg0Va6m58nIvCYLmhphl+oUTLQs5Sly1bhwdUUYcr5hYynIrBgUKx2kmUoRrt
WsUb4jBdba1opqjBg8BaKdWs4Gx776wfzC13Z27zk8jK7BkzoSVUIiP2pEokCFXv9xktdACy4rMQ
xHDj6rrAzyTBhsBEpk8k8zxMQIW1TAiVo0iRt2xGddoQipYkiIhbUZL/UpU1JvQ6o4yd9I30Tj92
NEMD6tXWxhWfcxR9Jbr/rMxQDsboOVBMktkupI82U7hC58MqwhBuslSTEQcbHJKgUfZ9qbazMCB4
kpm444Ioq77pBHMf2EhIikxEdTb5CiqoDAqIPSf0GWqLmEqXRY3IbVQis40+cgN4hmxUWXdZmluY
28zN2qt6XWwCoc5fELs9ah6VEX+I0wUFk3hBOr03V8ZO8cb61iUOwI0EwPyZBORN9SgEy8s/dlr+
vaIqTRH9w8AovS2oNpZ2BgRAAcYaxC+ktD7zQTwOgdKgV9MwnBBHCOIXYuobnnFpxGk7jhSaKUY2
+zGVgZ+fylXwcqAZwSu5KVo4Yy9NqUjVljN4LQN/+G3/MMHM5jOdfmJNBMxMbuunZ2favavrLKza
N731E8M65X8xJqqBZLDr9awKxY1bZdQogSZ5HEDPSS0uMru8pbjhHv+rNCmujhK7gPSTbLgVlTy/
YkPOTn1MVXXdx6vPGYWPWOGSl/dxQIW6M+Wcwiu03MtoF88UJAlVhC4Lx9neOxsW1swdUS8kRqzJ
qMKKiADlO3pA0/KWwgpBupw40dNJVYnyobV/V1QcjFkYlSQV8Y7vxtL2icTGNzReUP+rDNroCTx4
yIXo4VvvAhwsAv/JL9V6h8GXLh5wP5BeP2yJW23bzemnREOELxDrR0jIjvV2mFKhcD21t/Ac4Nv1
Cb5wPgXO2JoH+RUIYuCQB2ZWZebsCzOWauVXF0LLxxUiorpI9dI/Kgw7GNEHRrEebXABql9mBcKO
HhUbnE7lOrt/y03LurGIcXsqlZTNTk0LhlmDYyvEetDzGNEBwNr/OjmoAfk4aPqmyX9hU6uS5eoW
6BzP5cpvEKGoxAj7JNdTD+nzSr3Bp80nNquq78ZnFUoPFPdcCKCFJDEd4T34mpoqitZT+MZ9EIYN
4vY5XPvBrkMDIBlJeFQu0sbVz7V+Pt57Y3/kzmPmkZeId2IkI+EP4ZF80IM0Zf19Tfctze8E8hip
TER1XysNgUFcxZPqH9IEMJFGdpYvRNriQnpQgT+TrOwFM5tJIflsMM+d0F8cdxx0h/lHcULC5kJB
vvzRMS/ven4KdcRMUilRxxn7/gZDIzxS13ULANhaiZsJ5ofEaCtzjtCvTQAG/vSY1GKulQtByDqP
d4XDAgzbhjPQamNV9hk8fjHygL8l1T9jlhi6eNssrauZawHuRvxOYTj1VjrvMwTSLJZZQ2gKvT0/
cM1Ewwmut8GXKotH1XkjJakPoRdO3KQT70QZVV6lGswBuLG8MeORKrMRYSBOii3Vi2g0KiWpPr9V
5w5nqu4bfjYonkNo1cHs3gk6zSWuraptL3jtdNp7cun6RQeP7O07U+5x8gfZlGZRGugXmkAO5Qoo
JbToAOa8ksiJnADzJtqAS+BvF3m5V08AjQnIT7xLE4ZroVtCIoPRgjje/s1/Hh6+6fMbM0GHkoWr
1nIrc+xbMVOuaPuPAacl5QS0njxpvm0ZKHUTlv13i1ISYfCdYZb77yT3+aB+hk9No1M3Sm7lmsTS
qsCA98I6S+FWHQvLqEXXU9w0vlCseUFVZy/8NoOLkukk91o/BT/AIrNGPwFxS/6sEwlfFmgnaqrf
I86sF2ffd69xrweTo3zub6DbgfVMMlHonNm7IbLDpUmLOoq6LGRBbqEacDPYg2eQYGZDtO0GZPql
0bovvwxtk3ucMiBU5N1Uhim1OpG9F4Q9r2jqXrC6Q/+9wjd4oggG9blzhbrKypM/VArU76tt28g5
CJGWGKLkqCANSIIEGWt0ncwa0NeYGbIpYp19EGHrgJ63s82dMFbPso9ITuxNN3gmpwL3Kg2loq9Q
W20imRMX9ywTFBqTQQPzD6cwNqnJOhXEafqFnRhSnCBiPLZMJFjpcIf9/TjqPuF6CynhrDv9WnH8
PEkZdzRCoSJviO/GO7XkD0HWNFKcfdWgcshZHkd16K4/rbF1dQ8Zg/kTXMD4FDquzjX9V3YdZQK3
LaWLTLDeaA1LPZjIUbOKDVZ8mIZBqCJmuddk95BCF/uiyIPXosiMCg+H23y5jME8dlG17wk3rIsy
0n9wV1SIckPYydx0xm1M6egPUzyBLLi1XNcNhSSOct4mbQk4UDFpt6sk4lPZe4BKSZcZmwgA78c8
F9YO3Y3vIa0pSFPn3m2fJEQmbzOYqz9mAvM5AZ2dpaT1r0QTT0Uc91O3VpJVIReKCqu7R4YNiH7P
pRlJRUfSgpc52JJ+QS0KrF4n1LGXVrN/wI17jqGICqHaFMD6eTladvwUF9mBIZBDPxDPDuI1yDc0
VZP9BvrGfT5lNHTWqrkG9jgivrwI6Bf3t1t1XL5oystluTgIHJySjtv53VspfszH175/rGo5FP/C
XBwYRPaLRNBmmtZRr7U06JIwDWevjOl3EhDf95w4sS3YcX86/azSZvRFtBGojD2WABntCJHDhTAq
/Nvvhf1YZFsHukuXalbLH4WKHGy+8IQoUt4qcI/6yTUTHs+xsVbVRgp45ByEF524WAu7C1reiOzQ
tbxm9AJlO94hsbwRMdX9KLaAwDRuDsPzwNMQ/ZAX94Ov+R4tN8ZZp0daZSQR0iHN8kfg8+AfYjK4
IOlmdaBv8V6+mKSj3dvmNp0L0y00bo0JbhP3nlnPSXR6ak20Qjl6KBXW84hAdyAfoDiwSRAF8Xmp
UKKoXucAw1TWT9eRIiSjETcscAxkYsL9dqH8CvI8Jvz/RpM0TwuKUEqPIv5EsJGq/ioO/c4tEUXy
lWsl10BrfXaQJ48Vbk463lqVqA25vwMQcNDQtTIDsAMhX1dcX4OFf2MawezAC03lhTwEj2tWF7nF
rk9OHTEse2jTKJ3oi1WFJqnSvmjadbRiP3GL15zzYsWsfT+nodT+FgZ1G+Z+fVJpgIDXstxAS4C8
UByL/MgA8OhoD4OHmPe7C2Zvda0MCVitf9ticfZ5mO1K/qoiVYByCCnKQICUO3fPgSvqkwz1I0MD
9TRhMR/AjLEjLUCIRseNuE5Db204CiaGyW9zDV7MMY5m/1qqEcJrTI9EC6sUGJbgVD9wnpJxfwyq
G/Sjh7B7KooE3IkZN6kTxH0C4fSpGOiC+fpSBM8YH5OppYeXKwRkwvp5JfrLy9HHeAZ22KKB82Xs
wEfwjoXDCs7vLlfTx+c/AxnkNymRLpDnp2lUQWriy0cWZMF8scudx1qLttq7ouHsw8mW6n6hIdF7
Nfc03TYyCtm2QjcGJAQXEZythkYH4uh4wse3ROzzFabPylcn62HScMVHZQorb+Rr2mj1bGQyH/2v
lQgX1qRc3RJk1mypzRs7gGhYXLCyFrs3vUduaK8MiMZ2O3s8ZXS7BC1Aie26A4+DNpXd3C6PaTRx
Y4VDXPMTOsK+jn0UvM3m5U4TjCN4X9iNsWvOCHEYAzBSwc2hJOCizzAoXL+OWf/kmeJzANCOIZsp
cdcUYIgIWqbJ/bU1mm32aDAo0RE886Q6HmnnmmtCOztL5g9WM5kMoPu3I/VU8bAmXzsSDwMRGCDf
KAV+URtzf0kmqBEeGZchdmo8VF8Bc2CLN52RDnBgVp8oB3UNnmNxAucIgMppAoLChStvARzKLJiD
lrTii/fYcQabwCvsMqNMf0wdvooTK+p4nto8ST7CBtvsvpzT5RYYrPjHHI1cmSYZzyIHuBHqebwC
D1g0dCuzHcPu8m0KcSQ4DHwITvLGjocifAyme03mVrUDL1uIOl8fCU3ycqQmcyusbQa7ndNT+xIz
V1xm7HwNOMY8jnlue4HyvoishB7QBCt5S5EQWjmJqPdDnI9+aURi4j/RCMAHINGc57ZlmsAY/62k
IUfC4iBm2I+csVz0n3S+NKlR8QTp9jkZGMh5cwG/MRxpclZDVvHOd7oALid93tmgXI2e+nkFRdgj
8pNHzV7ObkiPACwopWcv6B653RpryIyI32jU2B+zsJn+e8TO1W8CxiE/9nNY+J4ajskRIT6UYujA
O1vewRKyO3G5efgKf7b7K6F4GcBM1ztk7IYag989rJZb5e+CVh5b6VGlRxgFIaisCRDJnSAYPvC5
rj4vsc67pxL9E0hkALzYs8GCceK3VSRLpkWaPnvp1udXU2gg+03heWNMBnEAkizyVS9ZyK1qvrDL
1QKg4tjnn6gHRO4r54N0XnZAbj9E10XCKzTpmSV6G9KkNYGl/Iz3aTAojgvVkb2xf2lcS6B4mdjD
rh12QsdpS3AqJDoccZbDMIxGLDSaUgcy1eZrcW9px4J8p645jOum6rub7NfKMcJvXvVKc24nslPp
yIRjvS4AkJHMbA6pZozgGTQUv+C5Yu0zElRjh09RD+p+U5113x4S2tBMh12aSA/uVM0ymbVColrw
P6HQDTLIfDKiAJ1BKIfF9i2yr8v+6MQPmg8ttlJEfJj4np4AuzPkxr/o+jQL6gb61ir2P6y5QRZf
XE+dfMlwUP1/hO1ZNkuFJZLxriNhGI/SVC5d2+0vVx2F0vYmPgekQHwjayaVy0L8IRLD1fxmE+a/
/TJOYXGl3ugLsdX88XM1Cicg5j3vic2vOp0sggIaeaz04tlwHLHHft8u3SJaxvRAdr3JK75jTzKo
A30usYAgyGLPvJhTATmXGv/FLg1fWoDhGFzb6otqRumxO/mMAwTG8KGZh33OC14w7DR5PdQRO1Wa
x5z6GfTKPgCwldQjTVJWodCuZ1X8qAycpNYdjPB4FO/37rVHmRhCgqr7YkIhpDjfXBtR5K/Jpsis
FXVlLufiAAvy67Rcx/EiHBbfIX3nmOdO97vQpcRheIvDAEgC7cupnoI2Mz2Gel4RAUrcCcFL3lHL
A/gS7RYR0EyO0IhuS6brOFa780etntiSOmfgya/5bban7O5YOt09PcVyEWXppVfOc/BXd+be/fmJ
JImoEMDnJLAKLwC5MbYoaXSMAqqC5aFoOYKBY+o3cQQSpCGTo4rwB5sSw+g+6N+x3p2z6sw31eyQ
8G2MhzYCxVBHu8gP2uEa1T1O0V+pDBr38zLhBGZfRLrvW5GD4rL580/j/wJe3nlH6o+mt40ee9NI
Tlobn3W3aRZF3GW5nTrTx18U4/FpymSzGt6CnHTjlYEvT7TWWLHdpfqmpvDNez7XYpXVrSKg9mjZ
Vou4lc3oSSIwB2+CnUBfaJC0IowqQVtYhufNUxFRrG0fxAavOu/voMMyxDQEDwux1VbKcs6kN276
y4KRjAVTc/WdTfkWv8a76bJYXwAGbnq2UNng2VX7crU23yIXe9SYg4vD81A759qe2prWJp5KVuSW
BOgGeFrYoFDRNDIVZYn8GRJ4TIsqv/UvTh0c2uZgQ/IHERzrWOL6rJB9aDGhQ7b1fXyntpvihOcW
oIPlyExrsGxnbsL7qqv0YInj0f3mM9ws0E+zMb9KyMDhA1VVnccgXsYGRiYh/3DslJpUYvWmNu4N
rf3D10llj9TSuaR97xAZ9xNKVBnpYBHT6D9gn3Nx2PcEDc23BaoJsLGTUr/nSBIQlzQrYZgC+XUc
VDTdgxjKQAmZumnid/oXm8yD/X0PY2pOkH2g6juq6k02xv5noW9CUE7C276CXr75Qe/4aOcrX2L8
JIv62YtALbCm2Jo0jV5hXdgTuBDA9focRYqpkMvU+nTHJrMndgAUSOqBjfqRmxLdSI7Vs2KO6IzV
juNPpBp67xtjdObZUuYDpzyb1t65+GfCLIqQ+VxJeF21arEkUdtSSxklL1wYr9eKoK4byYFQxc1R
KevTx1HAmZPy+XuqQLAkM6q/ExBujWr+73WIh+athb/wopWFqq4QE7rgmxYHJnCqbtngk1Jveotv
DDUW0hH8FSmA8hzx/U41S4I2rXzppt7PHYefYQ//fiP6BQLopDu7ZB/THde+bIvC7ea/C2Bt13U7
o4721r4VSAJNZ9mu9g5nnNTPlQfHJYXnAKsuRVta4Ry6O6QgYd5d7YHzvkBmKbPaNhW+L3CM1QwZ
hb6UrC3fgFFTSI7nZO5IHjUk5DtWscuc9KIjb2VLiNawdewaRkqTb6/kGx+hrJkTCN7IPvyL4Lsw
lk7f3jGtqspgbDJrBPRJTLkvsScvBiJ/7MdcslzzV+mxG0bqSdNWiuWnkCq2DznyzHqLmA2VLGWt
hDQYPp2D/ch5sNaJNrd12VsK9aEiWUVWkmS5UGYSSNg5hcLzWAvBbK5nXIi0SdGuoGPXBND7ARNM
vwbKNkagD6b6fRlENxmIoRNs+a6Uw/v+ErVnO1CMJc15yuH2b2AKG0e9FCAAqykqxVWyFvgoI+lH
gXFEOPDPyhcjXcO4zvhQ/9c4r6wmX5ty0NwdjxMuHDDGjickIg4EmMhYU0dULAUsZ4ST+TSL0Dpi
oOx/NZVdoYPTLOKGlgidheJL2RVRLdumpjSb41a55509J12xUH8HJVWKAhAH9NVgYMTzVADxSAzF
NA6QsAx8MEydZrLu6CfcmFr3gofHHqco9R8Axur9K2od33ySQXU645JSZA+MU/C6RMvksUuYWHY2
TllXy74gvGWwkWkKp6hoOJbZOvb4xS50fwGi3PKCilqxH2pM46GwWpgILJtaGfJOurBhCI1vzKtJ
TBnvtr0F0+rFkIRujP8OMxU1n+nInD8Q0vbt1KVwUIphxuN5GW1pyPIKSetAPG2cTpyTqGBBHW6n
zILDq67qgBeYRixKdkVzz8z9JSjl05l4YFJLadjP63Hsb499mwKe7pc6jilJWMK2QgW2Ps8123e8
PhjPYm7NL3BbYBXurdNy40DGCx/H75f2gGiTt3DEyIK9n/NmhbjuwYdrra7XNZZ62AVL2eXsyTv8
JM1S6f8N+JUQSppuRzDgsACpL989LiZimpVAizMhCFXTfK5GnlR0h1TqJYC4WtbwNx4FzajmjYpf
PZ/qYlmi7yuS/dKfyPOj0ed/9dRsMELRmTXNxLFJVPNC8NLAJZK4cz0GOz0CQj6cXWTDdGq/suw7
319NwC/F8ptZKooFFAAXJZcXBs+Ys/ejYb2v1biiv6a4VV8MFB67+MZ0xY4sRQz0HtBOAGVHnMsV
33PhMwHCEUNclzkOMJJdLt8P8T4povCQ966p+l75+oDiIEQvHaA0L7hxWMxEmjLBL5gLLSxTCHmm
LIeq35t7jpqgt0M1t6m2WWV7a8Bp6LmKKnVbPBy1aVTrHEKG+viiXMIfeYWRHyG2hG/b9PKQP1pJ
YzrXErSU23I75KbcI8lIMkbDPmBTVn9jxfsh4iQfxb4Sf2foA1Z23M9Eu1/D5O5vX7Z7GeWnAADl
c+ypw49SsfYBXAYRZC9pzkaoDukLppjhJCrhK30VoMXtnqUectH3+u5TNSDJPrJFKdqX3htfi8oZ
NoHFtHlM2QwpUTFrCGIkQed6CDRl71NtFS8vy/30ZjtdQL9ZVY+2R5NONdWNq95RxrQw0GcNNQeN
64RaR2YmAuoqASYiCCpBzcV8HbpwAO76gflLdWnSVVZSrT9HlEc85nwIaRiTlLV9HD6pt7uegGyq
/4d106nBclXOjF99T6pOrLxP8X0G8Nl27EBp1PHq+AfrKs0Ku44RgkCzYiN/OKT6NCiUsxN2fAgl
C/UZzMtCvaObwX81z8U6XecJ28R/9QiIUHjKKxKUjgDG0OreYZfVn44VGuOqtp28i2D/wy8VIdYB
ZfeEWPoBzWRpokDc2+rLjiPpKhFtKwUCSqyxOkT1oa1EYRf6FuZqNOTjxVwnKsaYh8pdIsTwuvsq
ERuu4lW7tZrDyzg5xfh+36RMlDjjgRos5CX3SXdy+UUu8ytQ71g2lFQCASXw2LSArWUReCR8WoiJ
+wYa6wUhLE0iJL/Xp4iaZ8oeAjxHkgWTb3t3o8KZRhi0t0g9A6TZstIfKNO7SSxzpdGPm5wOD2ad
W1FS3VOyQGcpxEE8WFDZaAmfVVj91BNXQfZjZYUmat0yw+HwZxyl+48nu1ByMiOkNUMcMflJ+Q4+
Fp2JH5XCMjoTRBqizfX2KhvitG3vHblt3oimNcPIYLjCZoOOz6/aqlgEY86918C1wHsOthVcGNCB
5mT5KDIOeep6PfBKevyKSl1tUNUlZ8YKhP17PMetSwrR08rMP1ZE/sWaDCmDrD4m56FQL2opufTD
JFb3hB8J8ucnjz/1KVM35D+TzkUJBewu8K+PtooeiV1vE7l9QtzVakISZkGcG/mnBYPwYMayL4He
aPI5bsQ1P3YR3BnRKl69umPqJ9PlfcGFwJsoY4r7QUo384kiYXXfsHoTBRi1AVURX3awfjZnKxPw
X7gyjhElL3NASiaB+9BTk65kjnWnuUStkoicEohtRZsBmHN6IXt3tCa9QWeheKP0fcHG1otO419C
QNTtG5WPoug3D2/Wbq97uqGiN9qS1/oR+haek3E4Pd+CNggnYYjx5BmLjGwoO/sLFwdaEF90x0+K
YXB0K8MSQAY+skmkhDLET5OEJrybINfBy+VZrxq6xsXQtTXh/Jpa7+/ZUcyM5331TKhcC9O6n33T
329pzv0c7DZ4xeaY1syLAaIkuqg1tyk0S/Qm2DnCtmnvfye33NqKBYyKbT56IXqTGNIAMQz4RCkR
Nrknd9u/2qlmpbxW1qtyzf+LA1mzTwF2J/oGgL6CXlURB+xCF/+3QpJnhHxR/quOmQ0GYiXQsVEC
uE3jnNctF6nvGIvtwrKFwGPcQkQvwPuW28/mwaf7637MvcYNBrpxk5BSGysIAtyu+VdQNzDai4GD
A+3iUupnU3HgTxQDGPX/W40WjVGQxAUxmVZ+DXkPH3G8+bewC3cHcxD4dqWbVe2dLM+GZMSHg7Ep
e5kRkJ7ljI+7RM8SA7MGJaIbtIjaXmbjXGjs4LWg1svBQbVRtV0qJEwSJ9wpi1hOKul1Gnkj/c1d
V4nkddXZFTrxINTlxZC66p6zImlAif+7QeC/VM8HYeL5nvHrhfuWJ5Kq/RH66IJKlMjCW+k/OSvn
94cWjI2IEVxt+09LW9ZwnWvAcRwDtjJMC5Htzoirl7kDZrohIPKfhedO+oEgzsMuu6k+w4t2I0j9
Lg+yJnTMsEWr52+tHNBLEIfI0RwMY6Fsqphl7vrH4W7mdhW1nSrX11RVbfe6mdaWwp8f+whnemqo
ZXRTL//zTTsHzuDhHgmZ0qnF7ql9CYDgsZ627JINujemCqKzJWGqPaFOJipNshMW20amKH8skZul
zZjW5HRGT7TqklEF83u/yruF+gqq/4hu9wW+RmdH2ryyGp3iMgjraJkCJOA8Jo4pHrxlslIbhE3S
GcuxU9LCzkDe4Y4sv9w5P9aoBYtBPfqMvePLbGBP6/bwzmhjvQbvpd+/2Ltqkn9QyhMAEuYml5lk
ihW0a9sbU61EKRyCSUvP5QCrrjRkANdgsvuRBi+ypVS6A3eiBVrNj4TiohQwLBicKIrskgFnvj1b
DoWSxh/xzxe46p8Di+cdLs1FJleC7ckx/1f9B5M6QIa3/5sP3e6sC1VLXqARTqaIgMsozJ6CTacL
6ouzSCdjR94J7XVhuvDkeZIJovh6ARIqWEff8rO3hdLkr1IKTquydya0G7vspTeQ1LPhqwklpQ7/
dSn6big0hupaD0avyoJoQGlwNXbK4KD5SqeZqqRqs4I0uBhG3Omicj/Z/fhr/5xyGq68nuIYv64r
cVBfXvmCtdn+f6z3D60VpgjHKG5R154VjcZb6qNBrxMvj7II9HbggmIvI0rDVqtD6X1HJEtVfypJ
NQm3Kbmml5F5akd34Jr9VWqP3NTdGnYYyWYjwsl46ZND3c2S9/DPbZHAE12YEi+9HLootYzLPzGj
01BRBpad9tOvxBHevdgySkCIhLl4gZokKhOUIRZJItkyRf7m4KZMm1EzzYzwP1YSGazqw+k6ytGS
C5b6CJgi0X653vzwbmOjEyeVRskaOMmOF496JooCcq6k0yO0Jiz7tWyQMKWAgispw4eNC8dTUAIT
HNLzvi1H4Sz6gNag/AD6ddVd1ZhcNuIOWCkvJ6XwDbSd1wUSFh+ONfPTaxoSgyrqmzUmR9Zo3WKr
FJF/U2pirXFhTI511EYueJqelgfvlUugZmWDnwwVglP04J2I61w7txriP2LYPk9mU6MKFxJbdjfN
kMSFj9XrpEg5567XNHqORP6bD9fh4m9ZILocgj9tTp9C1ktsvDs2NsalYtUmcpm+3KhfGzaS993Q
74anH/EhzEQYfTamrFXtgl7gjcKSDi2RJLWTDEdfXWThWkMEQXSYhTT8dFW3JCo7+AM2rxTHtSe2
VaqZmikZVVmYd3vMInX1GKwGS7nzKnDE5DYGJi5kVue0JcikdHR8vQrn6bll5bJpEewlD9dtAzti
cHmsthgj2Qn/wPG3YJLEEbCgR5j06sL136Yc5P0I9bavpwILqx4Z/scgbEl6C2dgsYiaePl0Kvzj
PAO721QEMPv1N2IW1sqwPKQLNYX1qW5wk4z82Fh3xQoLJnByaiqXe4ScYyLUJTJx8zHYyxX/CNgF
NdvQpNMyZiNVIhu8h5RE0CpEjEkfU48XIdWw20UGUP8AKmp3j4vhLMnbmcRNN76cGA8rVQXzGuA6
Aj3kUQEhO/FxvQMmyt4UdkXEtSkxkyyN4pypOQFWMXInbE1wLg0XpokDhvlCXddfvGuRH9tplUk4
pOZOm6iakLFDGA7szWt8QHmFiYX3X7zBRk1gcSOqlfljkhwDHlaxG70ead4uYL7s1YpK7XgYpzAN
HlHS9FmgcLZnDCE95QSKyAqE130C/97EV/jWDgCymUGCPI81wAWLH1qx3O6u7eDYIuQi+LVVYtxG
d6krIoB/3cawcRD5o7vs4XnCwu+jDZPPG+zExQLCN5fu4Ssdubqm1kM7tIfl/FO2b7wqGsvaDhBv
ag5btF3IahcI1O/3JDHC0jZq20KSCQSKofUq+3pine46BsbT41he7nooh39Dtd3z1PGvMLtUm3gY
xZEkC2cEZpof6qVPjQZKF7Se3O7HIDgSm3ZgXG2NuJdWdDqAo4TIYpixEl5T82CAJqdM+owOq2sJ
s3n5IRzJMYCLXHjHtYetZClhbC7iSJAs9Mp4RnZIMhvkF4KpxaPRFCXI7UzjSEbzjNdu6JQH/rYu
qifU/WjW1BBgpwReFjKgN9kVHuY6JV5MZHjW1mLB9Cm2RhcbzT912lUtKWOVulzTPYuEFrP7gVzm
VkeiMfBeUM/zy9zBQn+qnl+eUrKaW3L57qBdV5EAVR66rafcA3dzMS+AXrENA+Af+eHOX9fGneh0
ZJ0NbLOoSll5E5SMI7fusLSazkGXV5OWUzkASANHLOBDNirzKimwXV22QfGZANcOM1JCRe+UyfBi
n2Oxm+y4fVCb1wdcNBRBiCyyrddoTEsWhoBMMfaeeXPN52W/Sy29onFXlbTFNPyIMECfcTK3f9z5
OnlW8jUvXFYGjrL18f6vqVcZtISk8Ygj/GpkT1kLFIEAl+fvpL0A/Xc/EXx80CrsptCK7faESUIh
Ji2w/Az/MKj2SG0542fzMnlhKprhcAR0bFbS+Qxy5TGU/vp/Hz0uzCmnwFojHIsE3hvDI7dEjWOt
90qXYQVAQezfVcUfJGK2jPt/FVsH9FItLdp47jU0z2oaqieglMu017qnd7Rcn6XswUf1jZU8QlTF
AWWypEF61k57sR0518cSvoopLvpiXc0kzYzyrJEnR1xpnMWYnZ1kaFDYFir0qr0XE2bmjAaegUxs
h9sPYThcDYFti50ZRlN+dU4V7V+ZRvKt1jCZonJt0vtTTHrkhRLE6prn+ZmIRiy1z1SUOzMdbTyt
bTSqlaVyjCfbZP8E9UkiWbA3CS6e/TkIRRMsuZn4yhVKVIb5cqdfKzT99uiaUgX4S5XwLlZMi6Dy
6ziYOXZIJbGBQ3C8wQuCuO1jltORAvn7y9cbXK2QtvPQWJ2wX2hF6viQmYWm9iu5O2q6xxr4zgPT
j8mLS/fIgyYZ6+75vANNMY13/y3Q+s1qLtP7dflZrTx7coCXenaB+Tx1ask8ydSxoPiPfpyoiAe7
KvGb2xo+Kc1SJLWRrJvUqNnfyP6tHvd7akiZGM5Ot7u52ny3HCP0QtL/z1LQVpIePl+DoKe7bMRS
yUgAxfTbyse6YJnI5UPf4EFppq0LV4GXCXJ6jGpN/aglegdWKvfHCSlo8QyXbPuMiL9qO2pMWwBT
jDzffdgd+dZXzoEF0pEudYTjZ8b0o+FChJ4hf71Jv7ZpONHkyaTOfTTPVdf7qjr8MnZEXu677Xek
e2aWW2YEvDVBfw2cdFZZtlK9PtsoRmQHqi6yc9QhO9AtW6UFlraM6QDoI4wWQosYNl1REXqTaVmN
6Ns09U054r920fybRjhT1k5Vw2KbHeEFKYfxWtDOmBtBC8JMj5T538lK17fKuIGWx2CCza2TOb75
I7JzPFvuWxQu07LwPGCBSTAHhEoDBdm+3fbgi4tm3zaUPdG/HqlVgtHD1DPyAmrI/w6CVJBCW0Vk
0lPXL0rPYUN0EhcS0T2nTTNs3Ozd9UZ8xARXGl1PMJ9xV0QmDCc+ZbLmdBOZH73J0xco6HP03zO2
oRzOQwcT62RwXXwc60Iv+4OieWKwytxsNCKlXM9nQofIhWuDjPIdGpT6WTKn0hr2zcjoia25nCUh
nHbOW9rbk9LViFfqCyrlwHYvOYP9gXfAPdUp0V44i9CsTvwgUorzpggSiBvXhL7fo/CGQmDldKK3
ITIyL4pYaQDYnIafjXVNclT1yUSOX119yiBoU8WPY+IjZhd9j8lxRS7HYNXObIDRTQFVQdJONHgc
f/veE0bWX06x9iObS7spWTiXgw+LYDsGoNXet4/+USiiyG/oRXOGGcY1+p8Vx24H92qXNgkmwKzv
TEzFWkUXoBR+aGU/TLZdSZI3z89abZ4RwZw9Yoj3tQqYeThyFRVmdy72Qk/uw7XuTlXLCXK8xJsn
uGfyLhV9YjQcUlWGhmUSKgkEo2ISA3bEtxUdC8FujKRE8xuTjF2595gEPJTQYvOMNt1F4U41Wkyj
eYZzQinzLQuDKF4vDQ3jSzgBfigxsfLcbfE2zILugyH+4foDV4AhwG//LVvzZFndrIKg9TBJwtJ5
5W1EHq3peL870MlaGqgMHjbQEDCHKWh58wc3bkx25sg9TUcoTrIcfqtz6R4R0u4EeJW5i7uHvIc6
vl4hTiePWOq77Dpzv/ze1p+E/JWKtH9/8i73hElSFz/C1elM5FtpumnFF5/qNWNHu672iL14ZZkS
+lIXJtdIb/4nESkOdMrZzXhnviQUUkJhQPkBIkqGdN+SreOrqxNmCIpCkX3mmJPrtx3ssq+Q0RP3
7nR98MnYaZr8lZz4mceMggXsT5u0BP+HjB8ifMdNYsHI1gPhIKNK+O6P8GDnnXb0jco4KVtqm4eA
v4hTjHVXc5QQyXEUSa5o8+PCdjVof++CRP2lk+Ui4pjq/K3KjMfgaHdj7ScC5JoVBB5EApu++Y2+
VYZkqNSZEd9yFhj1A7lCxOpIgQQmH0Z392qK7zjBovSStMBrq3CxGYKQvK21GJvi4Q9r4JmWwH+I
GpjaHlPnnC1q3uxei43AkCez4WNRILdJPJKrxPzDaBUtn6EvhzrskvMvrvWqQfagF3Xmjko3HKgv
1kvzzRaAKRcxTka+FBC1OEsF5wR3FeqQhvn8ZQjlC4/7kGqnlLMp7CnGEba4PfnuqgL99S7p6KTh
UUSSBuW/Grf4qA7kcgMIYmX/TsdG6KiyWLHB5j3F3zbzk6Zi2QtyegBDhwfqJ631sr2WrJg88JgM
+FpKYIHFo0mAqpRTfICOANaXSIH48bqME7Y+L/N5hfoRTYLoXGC7hR8mog+vGAysoPSUKynqR0Rz
4wVnWOtisNCJxEW83dX5zM0lqoARIJx7LYghm0wjNHCd/H88ag6DGkVpBvYlN8PM84mb8pC13k2q
Ix4MWlx5kEP9/2gpAHmaTrhwc7hoxI7LOMbtLAj9za2hHjWHgXrzq9S563TXTfQFxRgIV3eGBjg/
oY1VAm26JIUvzVyV/HIeRA+IOQuuAOgPyIVKSq4QH4h6QI7Qfj6od9eLtfhJcad6+gOohk4GDJ6U
CRXKHWerIfjmRDWVirSZ+Zcewa4WVyiY5Bw/VggAp13FSzOTUMuVjQFTpMsk7uvd+Eleg4SI0qfy
jt+wF/+SuTnW0DzWcynawd7dGhKmtqVCajl9jWRO7aX76WjcNuh9GuOLfSIUbqvNwGuXeGwDNzVW
Qf0c9SieD/XDuc2T/HX7m8Tr3i1I1nuHTls+a9cyn7j53m9qVGKww9JnTa6NvsgUbM7JXSZ8yZEB
ZbPd2UVT4vcfc+Li5gF+jr7QaxhELrqCSjBCDIvdmWMLd8E+5jI3FM/M0FH5IEY6VQh4XRpPvm7R
aU/oC06xVVCGtMg9OgCHAmIRmfCs1ZdOkmMMGVccZibEx9x4NESJBZ4bIhwowwT8ZZ4oV3mPcFO3
3E4BG+qTInYVyN3MQ6ye+kziA2YTxqtj0uPFBSSHo4c+dCoQE90hHg1t1AokCzMJBLPj4SWnpzSi
jRovFR72dZKP8YgpJfcR4UPkHVw7XNF4tTzuh7Nq9tdxci/DWzGKNxAJ+yxoOoWftTMMWrbAF5pB
/BQAIQqrsStRsfsE6r5JMUBihUyFKPYsbtkINTx+BkVk0sO6oB9Lhovj0XcQmoGt+L9b76fImQl+
U/n9vAy2wvmFskje/7RTr7hf2bVhgNGfHpnGD3hA9Ds85eHQli3m3bM/MxS/DH3zYGBk8M1vBUxU
jy9K/OwqH6N/JlngxKCtAV5Em2zQ4m3ijAjmujM9DbEHcZUAnuh++i0rHOSNNFyISzpxqH2iVH3f
t3ROwBQYEm3p1/smLBydFNT1k+HaW22moGm//SyJ80Fjzyay7+An2yjBGEmrVyzPbCrY0err8UXT
GWf/LW8lEO0ytEUqu+sZZNYJYImt2glWUaRLyN0ZGziy6EFm8liTO54RHFHUAbRz2A5Ys6S9wDfo
pzMviBDnlWDNQqVSDLU5VejDmH7ZaKRsxoW5YpuHoPsAQMLA+Rqm3N97XuginamurXcPguugcwsx
osyQCg5gfoGGXIA3egiyjspE4+P41muEVfafc1ydTwkuzjGUAZ/3p9DL1fnDreVAez8YSV4EV1eQ
9Nr03JMi7OoZdpCWQzlvA0uWd8jDFYGwIayPURnyC6g5iNwPqnAGCvUSInBgXUUTtr/fDz+PNcyc
tyZMh6t7kdB9Sr07RsgQQWKifdyWtHbUAW+zoS1FHENF5RDkUjndZ8xL8JQMSI4F8MYw/dYh2zY6
gXu9tb1D9t7nS1WxmUvpDzE/Ua4SR+t3GDkS13qATpoFrywprPS6Y8IV4/kspqr+IeiYp3f2aHqj
QBKnHUatRxEzp+nATmbnQiOtqu4wl2HcuRjy1pM8lk9G03S4iww6jJvFEAt25LrCGdbri5Nfm3E0
O2uldOUmean0FszWdpZW4DWbToU1yDxr+wv8zdt0cCnBi7HqWaEETZbzRtY1xd5ZJp7fxI6EPbBg
8nq+hnnExGhwWIelgkjU5nbrwaF8UslbOupMR8bGgmcrxkDvsnWGNFkm6wUcYR90K8jUvex49T/D
ppFmp1t5nhfP2sCjMABA9jH6/i9h2aV4vBKSroi8xC8/khJlH0cem02+zQH0WmLqTk3jN+M0wwx9
PR84pHvR+QasClNNbjg5Hrh2P9efoubXkIOb3aPPjTjUxKuosltF5AwO3/EvTXqK9xh6At9RLrF5
MkE9gh6Ko8pmEUhJl57Ad2gGhhfdvuxa5tgtMxUKA8tqVx/uXpN8k1MewXRg76ofx7/DnO/+Dmjb
Jk4TIMj9Zpx3ONaAgvPzoVnqQi+aBPcc/ybxNdBYl9Y/+0yNr+8nCb9dJwXiaO6CPNI5bn8c4tdv
T69KN1GL34ta86wHiUKdEDqhdlDC+eepwkOQXeczNsg35Gwj1MrMc4XHYjZ3C34/SVXBn6fUHFkx
LqRz4DSq9/JOkZlPmxIpAzB4DJCL7F7jCgQGAgfcQ9cMQ9kMpEysU24lBj+kSN879LmT8XohfJlu
aO/esqfn38IXRdqsmwjw1dyjy3Dh9dHhhF9F8+lE3+Q8K2Q8Nz5lkebsK/Gz/GT+SIJ/OshjigTi
FQIyFsOt/ybcLG9um4tq4Xtjdjp7cHbclqCihGC0bRGBzpqJ9apJ7UeMxN+XV5zv6fjT8pn5quu0
TJBgZO4nnDQDkDkAzJ6iP+CxovCtLm12X1BBllX1GCueOItxzWC/Y+B3zUBdOauc3Vgh8KZDpufb
qho1O7ucYnVxja7ClIbNAF7AzVaCaRRP+ZrsuhF3iJOtkiaCgz1cxfEse3gUUbo427sOSl4XBjkN
+48UL6uDsefwdKUEWeTXwYwtzxmZmY79okvp72R5PKPRvUovIueh0WP6NMCIKT6sINrPHyiIGNUA
EkkBin6WA2rJTJ0hC6+m38/o97FwigCKKvRwGq8lYHdgGFsoPyjx6rOgnssW0NAIW9DAdP/tajSr
2zoaEOjmVcoCvDNeNCny0cdoXl1XmQmtMJZek4qo/UX3g1YEApULQyHFmGWh8tZXCZ2T54a4/z87
H+jQcdOe5wh5w+PQwOIFaL0A0KhkHbbjkmnv2k+tinsUlDwTsblNInU9O1Ulvoi4TwEo/sH8uhsL
CjzzZb9NCKPPsNUvh1YwwjiPIwLz1UxC94G4M1RczrE/IK6dipcu9C0wDZpL+4z+BfXJXOMAWTyF
nlMqsODBQmi3/6X00ldF2T+2cGjGzX6z9VePjkhV//+Po3zoYpI4iu3vJv87tQ+T17omgULZO/sh
jWF9FKlzfDlf2dEgOyNUNAbPXL42FYa54fI4z0zqJqY6PAlNnth2P9p/XyOZa/Ga7XEGJ4TYYx5B
vKF46itCB9sW+blG47V7V/taIk/Ln9i7VIk26NiF1Vi2jfPzRWIaYk85DlEj5GzwBkGcH7W9+mKP
+QYWp9KJZYydVBBoMZvCtO5CuxPcCK0n4HcsBL8oPTopKwsNT74n7IRGBTgueb3JwH9jd0+sx2R6
Z7Dm693ep660c/PoodIH3L/F7rfSAkLCciepoeMJUBPTzr+eAFZJoaRVOhRUPsLvtMcz0t3dkG/I
+qcD1Up3kgB7S5ZuwfCpyNPmJ98Fk5QZDKyyvlCDgabgjI412yZAoxFrxqpVdZEbD43lrKccwZNW
xWXFxUi/W3YWtO7fuS/OD3ujspqy2NyN7iDGNF2p8Dnrs995mPfDlYk4hexoCbVdH7c+NZCKukoP
rS2OK9Vv3Z/D18YTVO0cEsR64yqExF2e2A1clArVKyFvlRxodDWUtJiG0mZq9ze5NFZDjWt254hT
p9z1Z+KzQHiJz6byX/oN9x10xQYcrnGkJIMLb/holKrpf92JLECSgMM/cwfDRHOk5nQhXdCvfoC+
GB8Gd8T/1TLPDyL291cKUH1zeyp1meXbKwvPetc00/gInBhc6+A7iFm02o5KbN4Cl0A76yIYEfy5
njlluiPmo7UsR3JUrFgIMZIXrxO2O/ADcDwRwUvTNh2FjDRpmKbFsT/KyPjJDlCeImttRm4u3tzq
S2JE3VhaOF/k+54jjzF3694O+wiCMgUskmjkLWd8wdirsTNE6LOcQZR8AGu4ss62+pKbpzHo5yMi
mGmbOwowugT2EGLxpfp9tyP1t4bjuu+a7pTUq79pRaXGtUnwDqjwgElsSe5ETvxIZ9lUzJjRsr76
r6CglBqt3KwXvJoSrfk+rTX4jVeFY12RGlel/6u/THRYZrhXMH/xlY+o6VCF6FelWjMo5VgnTB+C
58x7bGjQXUiykXtQbsMMluJQR1a5gim7sLZLn5Ii6sDDAJE8f0UtRYdLsez75Af5/kHEbttxUrQu
s5zMOKsJ9vPtIWF6rI84UNWI1dXHA1Q8fw4fO5b/zwBLiQ6+GkOLKteRX5cWnBzZqERcPTNWx+J0
RmHNsycOCZ/gRhjDOmRDimWHIvwMygx7tD76agPFNZwJfn58LNfFM8N2RhQhNz3VhbjswC/K/946
XKJG6wxDTw6D6wYU+A1wBuWoeH585xCF/iP2W1r3ZLkz2NkKpvqNKBRVM7mQPHFSzbGaXacMNmc1
RUU44YJuCRtKewhEVsoHuGONXK+Zr9Wee8yco7AIQ4/S83tJf2SuDgTk+ku7HRdw24pAofxvQro/
ZkBkjySCgH/1vyX1pHSpT8Cr5MToDZND30nbq8DhU5Q1ekouRmjyfxfLVvmSfa/aWI+lkU9Cpg+B
FBvpyiwbj9p7M2tZZAxAMCPxEjOkIO/gxIZK0wdAp1U4SOLwIml6f5MxTLxOBBILqmMRR+RQ7qU+
BMzZOWbOIFEsq93NsfIkReuMqwTZg7Fa8uI1NMy+jb6/fffvQg8CbOBTkiU5DdgutB7tbc9mcgLL
jJDZyb4Twu4do6OwLt+rjXKuSiGqjKXEdyqMZKCGZHsIoj/Poe82ArGIafMqRgkIf58d3b+TNLtU
c2Wqifng1HhdSp61pjTDttf6ird5xb/W5EEsDdWuMHYCF27xUapXnZoAhE1RyOrD9hc1dng5hC9i
K+J0xx1BP9sxbsyGsufm9NQ8w9qkx36udVpfk69IS7qD4KC6oLgb6dPdixlnTlANEm0WO5IFJuoW
GNlhVP27vz8HkgZPdKEDaaHyLQQNP6gvBeSW2tSIU1Faund0lfNyYfpf22hMzfwHhTOdDwpCiW/5
O6X+J9f4/aEkrNu6oqWLE+2Y6jDhBEAN0AHMhXo6fQDa1xwS2KJiwH+xzhU7isGV+zehzZ+3P1A9
+mPealt3qRNnXFNUk/Hndw9DzrCe3d0LOjtAhs1/I/yLXohe7o03zO4timXFbA5rKpvU+Qaw0uqv
ULlJGSFNdkbvCTk43KhD8MKaiQvX/AsBwZ0Ge8uVDZqAxf8aFjqgZifODdKS7ZTDAu+MLN6Edu1r
SV+8txniLJYM75VB22km8ogg/4jjpzpKpX38C/c3vmdlUk010nDAdgEAnnmawGb5G0j9gslonGx9
Jq04dw3jgq+H8OVjuNd6wi2l8vGDtr6Si5eHAbJaiLgesC6fmbJolhV7UrhYH/GTs42ql0TZW8bt
FOQ8pGrU/8mSzbu/MjTyWcB/4/CYzoyYf19uhSl89ciS7mkxVTb4u18GsLjzyq82PLRxI129nBok
9PAGuyJWIIQCehDO4iUHgQJa11Pp4y7Pn/TwRhw+YSNcBLC5GDqSzyyOE4aOtsJQpkFWFpX8v06/
/qac6COBLHZj8HblALJQPAf0gvhqIenFR6lLoHzLLCco9klVVqJ0bKRC1OOMeajQBQqZTqpZnDNK
7htpTptkWspMRznqjy6eHXsshyDxu8Oq7QB9m+B/LLzWjTysJqvrWnpG1Vh5tgOtWinWN9pIO6VV
huvcbksDGvTo1/zGCGT7HRmPjKBt9m9ua9KoRBhwV3owa2cVH/+uQV/rzOq5MExRkTzfpDUR45rm
vHqmw8l1ieZMc4Luyv+7SaXD/LTDAbmA1bMgAKA4+Zz3uBGjqi75Ii8HHk/aEGv1+2NBQwEGo0mw
vZYF135gEX7OCYmMmJv+IwoZ6moxiwpnirV4OdAa803yEaI2/AcPeCj6ExSMRMrr+j48a95d49Yv
3/3nYreRjx429ZcZ8hNz/GPTZR2D8kUJ2qd665Rdxq8OFfMlKpRZNP/hVjeZXzsuhd5N8mxyLRmV
u9COj/2VCb4rI7z694UYrP4LRybyYdYMxN5fIpmCfvzvlbfxtO7XyvKljrPZAjjMreItTCq8fdoS
5XJreh5goxkk/FZHLqZMHu2DmfGcOBjy/yg9PxtiGmK8a2SNAglwl8RsiwauVJgYd7cTaSLkucZ4
jywaNscr/7fpBd+ZCPYqJREaHAjZ4Ed7JSSaaP7wlbB+3PTnQ2mJpQ3tyDWa3qgeS9b7b0JF9+SW
npN0cyYm7El0xNe3K4aEv3X+GP7QVYDB8nXvSkIWlHUbmqB6G5Om96k7pkV9cspG7X/5IMs6ipqo
+GMqWSUH74qM11AgfCN1xfsD7L7RkcKMR1Ur8JLmMz4QDDN9CoYpJ6PfMNLCpABG4ctlyCBJOeKV
2NBXeM+AgMI8+SC9RvZTW/Hr3avODlczB70imBNZekPmnTxrut4mLXkM6frkgATK9jyihPGnwWPF
rVwo0S6auLjPJ0zip8ESVcji8xQjYd1VUBqXa1l1DzzcP9wTybJb/Zk4bNLxlGvZSht3zdIGaTeW
x/3git24IbFPd7Cjyjc8OQ6pOfIWKhRoTR3BB668JHYiwnw851OBE7VLNNcq4yh4T5KMSeYeNtYI
QM6GXTVCf7P0PQpTqO4gaZ7imMr8//N6qoa+lPlXaT0tHz7k6I0btHJFhTGv5ESaiSlh2IOvkOoh
0EBnlfuPCQ6Gtq8hF774YbM5TlN2E5uQOQnwZBYrEh1vpITl7+fXyZNIGHIuf46NrwlkQFqvlRhC
R1WUJuGMDyiUVgc413CifmvmgQlt62EOAx4E8CLZv3VDnMXesDeq7WMEXV9jQzFfz0EUD+22+f4r
HvEsUB/6UQhr4i+lfeya9gLDtBzt6SSqss20mU8irQp+xNxrgv5f2jPHmGzu2nJMUxBdrzCTJ+ED
vFsuf2u+rxDv+1oXcBRTYphoOVryAbE6EpyqHqUY6Hi4BbzlDgjCyf0j8AFfooVxNIoyYHn2W2CV
HXL+7VzYUKRA2+A2bNsVDJxs5Vnjyg3dS0o9PmSXT+Q8S/Wb+KtR7RF4+u3X0XWd9G+sge2o0ape
zQQadKrKVRf+2JxA88NWqO5/C/kvDI5f2IViFI27SIIScsy6gC/PFD2EzvZiLaZnbZQeBTrD7PPe
NdYfjk4PaJwQPnXIHQ2HujH6jdmqo9daBe476E33nsVpE5Mq87XvqQ7Kfq/Crm9rKotMIMrtVJYb
EhmjstOGNZxy7jpwSAP9IqEfxv1l9d3J0YdRyPhlBX+2OihTc3mWM9Ya/1sCalVTxhasqKB1OFbY
/ceJJQYGIuC6WJV80QEwcpd3+cpgyl0YHp8+UDO5drqEM2nC983i6QsmNBIxx4CovACEH6HARccV
AYQRHYksHe5GEMfpfAL48IwXCJuOxX2iaYqTf6X9xB/PRkfwSMpmA40TH3LyB2pdWMRrazTGiRn3
d6XYJzlLU61Xj/ZQOFtPlaubRSrIY5TIBNG8cBx1mSIE9oFkPCY+InObr/P/UQsQSfMsYXbNdWw+
VHebj+Orkh0HXPVPc8JqmDf12KBVs/cz8u9gm9Kr5XGPWCUkDsvwaFaKPLWz/RmdR4QAD4RTkwT6
fmFMnAdKDmxpvO/cP0/wegfDINf91+rsoBFEMF9dKsq0LwiLo624cCSmh0Pd2jMCcdC9FT8O52H6
wGZZfSVPDzD0R3soTadPbMknvEmeu31EoGryqKuUo+E9m81EksGkQOZCGgjN2LbP3ztKm4zmRDGE
UIQ8K6vY4tNqVNuYm17wP2JdNXms8Y+MD4XI9WfcyN6xXBOPCFt6TTeYGxGw4J6VWjQ6uC6BhWiq
VIsP2gtQPcoIrw7Gvh6hkMieYpXupRNqiSfKhWCvOmgIfu4/RNE/4IcIGYUgt1RdTM208PGtGWaN
MqAOGQxtvqr/ha1DDSOPH2ei2alagR4tUJiJOfvGCi12DR9QALb3sKfdQmgMDX0MElwf4NUdmcRm
Uqzcq3Dk3fpdCn6N4KRr3KJBOs8Xl7PfY2UnJzYuqE02iCRHJOrH2iMsprJ9qY6e1B35QNGnC8/y
okaW+l91uYnz9SMmMBViZuQwtj54gykwtK9Wcexj18iI+UJY6rnSX6opwiRQ4gKqDwwWKoqsxQRB
v/yvoolDsaGNETb03N1KoaHq30N4vV157poa94DTZ+PJb8QegYYZEe5+7rY9u8vL0AxTVtKsEMCM
sIzcVXucDLGoiQhAGqgbdAUgWNqAAkPPO9AuffByX+iRNC3vkepalsA7ZOylerx+eVBbOZwBRFNH
TslhqVdRkcnlyT7BMgCYNsvRP81pJYbqgQ3srLnkQxBqxrkjiBHDEITsOIO0vCUeccbNhc87tqpY
GUyf6r+PEeycK1fpAaDVTpHlWbHFhkTuPn3oYJ/xms8dYppzjMOpHNXN7tiZMsj9bDFUOfDm5Z4i
zKppuCISucN197736WprVvvwxSjyZiMfDdOGhmdTU7dCAlbRMVYDXd5Vc8sKjow2stBVOP7Olx07
3yh/JILEq1aCJQGfkQh4oeovTHU3Zo5sGraMESx8oQsh2yEjJOtSeqd/ExBxesg68u3Z0GLeG/Vh
B9cAHPR1K4/Q2ERrss3OQgSyff3IJ+8+gXoKTgwj3i6x8wA8MnJ1usI1XoBUvf1JiwzLbeS3lEB1
z3A0LGeMjy1spsqUZZn8FHE2CPbkKnWV4Bim+VnG0eh/AoBoHDkNsuy+oaQD/B4hbQfSDdTo6xla
sEeSeN+1RMu6Q/e9YnJahk6X7XuDQph2fdgys6/bGGz7o5doY7vkhXcRl1jhLuZMQWXT+uH38fYw
g0Ytnl1dsrv3LtRxri9zQPb5wXmwCvAFYbxZB30qpVdg9R3XNtxNRX6aaX46+XF2P5rI7X0u2Dkd
7lGzDXqXeIu9Xmn5eua88Zddm+qG0WsdITmFsm9KbSaGT8igPmioaTviz3qWGq3NbSMAdL6s1pTw
I/TPPoZVuICprqF8T4mvfIbz5Q2oRgi2ukYynW6BZ6GMPo4K9ACa9ZySyjhS/yvZuRzOoYqOw7Qa
/n59F+NdJiYFgXeJBtTuflpe7HZDvNGratgUYCm7DrOSE1EzD6jdPlxMwKnHTB71sXPGhQTCYiOZ
dfDncdMP64GcacdlCFzSlmVLTZTKUOutUHxTCuexK0zIbIl+5ee4zDpE4QHRX/j2hnWE+rzxTLEB
wVwSeUlV9q9Jy0iQVjc9/SitX6+vuEVqf0zYaBVURtyZW92paint66oOB+cObadTPXI3BTKs6gk7
SWMO94qB/inv25u3JKTn6L8meAKdgppc8xvYsYfQqwMzPldtRx2qB4A3+6DIiT6tF+QxEOylY9jd
TYudH0vIxtc3eMcae/WDqJGwefLFIuuE7mUiJZjaklgvAAsLSOh/faLH5WKu/7JVYac+yw7x2IFn
tSi0+YxA8FmXRzRyV8ivZd+toZZn8JEX3EkEc5Zsn64jikLYloCet5Y5eWWCD0/x7UNvCxPDd17u
69H6+fO8J8Fuoan97xKMrwU+v6waepDEqyyJXa/wNr5Ld1RiZbljA9U3bNI0Hr6pI2WGmwYvSejX
aP2bfh3ksJe311Dl1WAbHBgU1Qo16O36TxulL1rFAOk0VQ6tfYc+6I+aXbb1YYMAG7SesQ/KCsu1
RR0kRqi9lh3Mr1mWxtENJ56GlCQaLsBzv0o4XwXuu8ZJU84W1jIkL6Xb95qq2bTU28+tT5vf+ZrI
wXT/Xu0QpOHuMoY94HL8FxrinJ4/wK8MnyvyhqPMLDLBXeMA2tFtD3RmSrIi+c/5bFnoH6dVFSe+
w0JtDCNT/Q+ltGzB8RAHxDGXeXjk+dC9ftCSzrfgVNUSmQ6VYGBExzerTMBvzibyEbU8JiqiOzb0
8e4wuKkqmStpVnrjaxGA9CMAvhUYEY8X4W9oq8oYOvP8ceu9fgASLLOu/uSIRbeqUKzEzzbepXAN
49Sc1vZSP+/8+BzzE7pznkbAGWhGL6oBQ7+F5rgd3n16adN3P6VGbAbrZUjS99tq8Q9/rcDajDJS
mcyCrc7RqyKzZGs7GGTNghgx/e29TlqDBqBcybmNwxYeJfrh2+A/ZVQS84xEXXYirAP7yLTJFFKv
Sa68B4fwpaElUShWVOxCe9kZlOEQrWOcny+eMdbX5aHwwzcSauX6P580IBAAojNU5r2mZqMLtYpS
8zmxxM2jOilmbQjnRnK6oHzrJ/nBRJ6RZITnIvzDxTrRcb4FhMYKHc5PTkB9dP55VHhe88280INK
6nyPK7PPebU7iq8WlTeA44tQcPmFYWzAtjdXQM7jmpCeaf4EC/rF1CNo3/oP4/X5dqdBdh+umiWb
GoSg46jQ/Wr/pGq6fxFCCsPlZIW18PJnMYlh3Is95COQBCIF7r4HlRg6kUZtrJRT/p+hyTyl3/61
RC5Bz2HQUXJ1k2uJy7+65RHHL9UC9O7LM7MOZQYc2Wrd/sR7A2GRQQKAQbMIeS9pq6VciKmcB0Km
pRdq9RdxjtVcarCkkFfo1EURFSOmzoDYgqr3PVSGt/HWDz9ZMNZKiFpcVJhkjYSumcgemZ/SYACU
iyJGGLpWZ2z1715z5EXV+A15NH5nubBXjfJD6Q9mJ8xc1p2Id3XEqclg6Pl8NgyQ0sk3/tvLKZma
DS8tKnWyjrPKB9E9xjYxOQ26lV6l+NwHT7TiSoXCyjnYELXb3OgGSMVKOUPWX9B+uqBPufSGZ+h+
c9vPohNzazgWNg4LggIy/II5EHtyd1pswwrMGqN43FYW9KqkbDSp5yqSv/Rs+teklQGFms/+Jbq4
gbEqMRYHj/pAKplFFe+k7xw4V1yCSk2g+F3pkoa8GqAOXMu9SzZEaELEL33wELR9XiYemEthcuJL
3FVIftT8q/UPUN2R/xAWuMd0KmxVEOxDSENXoIkmLdNxrMOQcjZQJlPZbKnqic80p36XforMJXhN
E3gYGRL35PBNQ019oX7AlZMf6MDeA98iZ8zZH3EKBPaiSQuG94Kr0x7uJiZn/MqgZ2BP3QmjlF+b
iQYrBM0h6f0mbZhJHeDqtKZF580TCkKI2i8bra91uowLyACOlEmvO3sYD/AatQ6U6Abwh9n7vxjK
pbbe0WVyYqgnm3mVKMKU86uwpVDJak5XPItPsZ5OAinJhiQ2e22KbLrWL5exQz5Sk9j9dAha6TTw
MpDYRKH55dedYjgprX+nyVpSfnoabibXqy8YvUD7wmi8uMdeOnDUN6ql4ArW20lFdwlrCho0DIsb
cFqbtMCikrDYwDK6cvCVBAdDIKq75Al0lr0GlhH94+xTQSbxOpOLtdwD7RPnfRaiq9y4SA/6WzH0
7zYFoOOU9ax7H4RPKm5jZfnL1Lm/j736WdWV5F/qPGXwUkjJ7/RCYyRyH1h7AmEIe4PB6ldLWx0j
/ohbKK/pEOC829HdTMyZHmmUCXGCfvDlvS9afFc+2/X75CzFYHzxsD3fx2W6myEmJ6WCx5EKn84j
d7yZR9Qb9WJSuRAAHLEA93tkj37pLOxGoQv2/8FI0rLzvcR+CV3wMy92ENq7SH8qhvi2bQFoRhji
EqcsFGNEkxGWUc8NpLmJZJHmcakUtgwgbAzHMDp1tHeMmq/8rymDumpPT9PXh7aBPNe4usgMPY0d
txANIAkgOIWdzLXjxVxFhuyKZheBQ80cCPR2DfS9PsLgPS4k6ey8Vs4q/XpUNeTHH2LSy2eAJFeP
PVr856kTsP/hqkniZRC3SX+75WDT6Y1+tG1gMQrzaHR3COZUD4Q6MmQ0uZk70SBMe1ZVmC/1905r
+0agndmvu4zZ5WlPFzTld5GQXxatJQ7su3I0vbHUo6bgzFxQVyia3R68ulZtstTAp+lFl22LJYFY
4sDjHWhywOj2gU9IBmfpf/JbDi6Dn03mX/rF9OfoSJOLO47im+wJ7lEvZsYmemtCYlJ4/rKkhvCZ
sUU62ph+r/BS0dujkmniEwxxDA8hah/fFbVc4jF8A8+CJRIHCOvA0N1guPOFFvLTsowXN4IUHl0c
islgIYzLwKB+MgXp8HD+AcqI8b1lGw60pS6OLhoJdemAZqVKAd8h9MRWA2ujX/G66pEfPd3RMPya
Ve+DHPXTZveJef1KqUKanaWl1kwKuazbVghESJ09zEZt/BJfSy5VYdUD9k8Fpha7Tx40ifiv2uUz
tUkysDZUTvodqJyZClsp+st+VkJS5U7i/N6r+Q9RNzy6F+/XELq9CF/HZwzBxknRABtTtSCgeGjp
/GsNqArv+4lfFED+tP0Rki3rizZ8gcYpotQlJQomgmvSaHgqcvVTQWoTvBegu9yDFOGCXpzofhiu
jZTJ5AQY0tftXaotSsZIoVBqMvaecG5B3rkgI8p/pyRf2GWBDzfxMErDO2GvOHchcdeEQwB7r2t1
jXtgfZwJ312W6tu0LiOPWyVrwMqojfX8xjn432f1zhdEYhe21l6NUU0qfH3cgcX4kZo3rDtCJ+c3
4SiVeJzFWa5Mpv1Ay0Cbzv2u9UQlF+39L60gJoOQtqeUevFsxSblqGjCVR2EpDrdcK9La2cwkRsl
TANO1T8DSjSw7l8fVjFercuy10PKi/lvVyiV4Iv4ZsohEF73xS/HVBQQfoJfxklIVg6d6ebNzokJ
+imXTc4ZWb8niCkbxZiJeZA7J8Lu1fPUSazH9INI8s15AuVYZZL9gA4OrFkajnNAUkoKnsdePePW
mrGcCacJF3D7pr6e3B6/5DZavSxWSifAfzWIfF0Y2KKiu/W/JM74dhsfLStGg7c0grDio8whi1Pv
8cdcQagKUpNELHm5jW7iLZFIRWOTS0Zrcvr6yhXfj32V6dKrsSGPmJERijoDMhOJoT/faJa+Dol2
85KHPnp41LyK5pqMT08gq5QbHHMdosFBJtye06gz0lOI/1vO1AHNZXYKXC9gd45YwmK1VY4PSJZe
VBex7MSVHxI0Q2EmsK+17wuGi6GyBq8RmdnvK7KnLbXStScHQCK1VkrBilOar2l/HEx6SbUFFD5M
+zfNcHQrD+xLB9kkKPD/a8rmVqxk8RSmYti1Lu+lgpKlr1LrDKFo4jzRtZSFqOV/injb4oamf1tz
oYimG8Yxn65PUVId6EDmHNRuFBjc0IMMCaJy7ooByJI8GcLLqimiZvg3g7QHkOx0C7I+ExRFdjsa
JRUzy3PY/cBC84suGoKp4/LxhMC375sAeLFAjUidy1eogNsDDBOevN+y2tPlWyP6rVdmJs9eslYq
AadIcun10e4t7R4BO21k9slJ6pC1BMvWSBs9RopVcG21v1yA9Rwlp12kU5VBHKsrUTC0vcf47LE2
mW0UqTuZM0TygXNyen02LXSGPF+zfMpdWKdLE3qNuabAg4NoT17ouIA7Dd6LbCdj5S3ajTsd3ERB
4G4UAQdwbJj7DY94HW0IneAdIuJ9mMMr8gRMyjSREWhVPTZNMfLsC+nqPZ2GzPbe/wwS7klsQCM2
kEg6k3J/Zt5kebnWukogkCkjPpU3VJ/LRUu+dVOZ3MgAp9B/MJ1gXjsQ7jFb6/Qa54sg+Lt7/i7y
BE2dRyE5rZ9Hwphk1LNFQ3s21Gsf7ZCHKabJWWy8zR/oyrEww2GZNdgmAi7aufxK9sWciuPM6uFJ
yqvLK8FQIXrF+j7oVBBtXTfC9Lk4oc9sqA1W3QYniilPxKwA8PwWtcbAmf1gJKQrtRezr1i2yP6n
aT7JDFqWzUCLjFU/WiaOEZGXOvrE8KjbojWrZHWzN0lo/1+K3HIF7ywHRTjvF0nju5s0tYv+aj0f
F/JRC7idqMZcSFPPEp0EwTgDOvY1wJhljo13OXtSatWz38hjOjkujdRVR5mX9eIxYyDxaRrenvti
indmcMb/UbYvW/Pnw3Dw5dloI6EUlzTDqGCkAzwHawVuR4XhM8/P9W5C4obiJGAd/l75M3SBckun
6vG1S0u0xwDDugmKbv1cI4eSmA/8sNKyWKaTN/aHOT6yO2J3nULXynz4SQOZXJEBqphf8CEF9dE6
GBRsaudSb4KraXq2i5+MM3LCk7m81JPlRPJsuhpxz2nVK/m/S954Ym//mIh8efjjLp4R4O0LmWCd
6+OxPfRU8/pU1+muqTi7B1RMAMb79Y0RAo89ny6uU/hyLcwaQh5x/MxeDwdtuQuWE8X+M1EscLKB
0VXmVrO08/NNLQuD8zNgnrt/jVRuGMLLQ3ObLtL9vXh2LdTuqtIdN/35ety786wUWLSFho2Ft20m
Lp0tEBB2JGT//vcrRvCRnGvXb2B43DsHfbJ9lHTbm+Uz3219C0YedZ7M2XvDjkVqgoDZKSR7bwXH
Ekw8lFsiWHNzFOIU8nhkrwMDIB6tJW0yXdj0xdO3epM+AKT8qnKrzlA3Gqc/gGdy798CL9dh3Bl5
1NlXtZXfGO4udxVnlrMePQyvk5N/1DS0n//idUIqsfobead+eobzh3O77d7sSUbbQml54VtE4XUn
uPsP0o1LeRbylGC5mjs4nW5HHOEcU/PwcmyXootIDLMcqLDXy8WS8HuEWsJ5PbdgqufRS2I9yFTW
ZWdjWmbolAW5Un3LUQ30Uppbj9BRLJTi6WnY7+JuJaifftBqrqOAyFWNLvjpez7FFeNALJEWl6Ss
IpqrLVsTxXALWM9/XzQHq2LUDw6DHEGhtiagaCvEc5gG0oS9vvchooHzXyPe5hiGg2fsYVEsxkqI
OqYBII4yn5rpgDCUQ3jhEwtNgXXAmLSuQjLtZZc8wqThoW+93mT6ZhB0DAZ04rEsmT4umY+cAwI1
JSfYVUWUj75BXaKPa8FRnhzpfQgCmd11zE3w9x3crhEqkvuwiEKV7veVMSQA4FNdb1k1fe+mLoDy
ON8UCG32E4ZhtaDG8sSXqddfKBt6t2KkTmBKbScKFjdra4VFW+N/0+oS7GnmcyiUKqIADYYhYGFs
X+34dleC8ksZ7lNxqG4Ug9ZzrNlDnTQ+5zzEouk/Q3ix+0QYV0T/RAfa4IEGRlNRtFlKYLPJT/gY
q4evAgY7SAknQDLH4BwmTUoVAwKmMXyObuh7eMsOTzJvT5VVGfU1kSlHWO0imzPiDEqGI0gxwxJP
nqaNC0w+vSy93zg7iyxb19wuxNMTbBhfFc5O3ubk/WYI1vqH/FItLMfAWDeFhNfI3+v5ymL7VU6T
Ycp66geF1/NlsHFCAE6zxwx9GyBGG5D6DCs3pqeuwnSILhkCF3HpSMkVYxnvFr3+FzO+hVG6xh8s
dVJ6+Kdl0AzWHYgwGgxM1jQXdvj3tAMe11GjK5Z2eTjpnKZqzmPUMa8I2up6c5oJNbbDTQycIlor
EWNlx/k2K0PVD1pV6cDftOFYcxDQgN/uM0wZ2IUV+6dMLKwQI//DebN9IcR4caA4RSAkxioZhQ8B
FdFpD+7fYA1l7a04tjuY6D2UGqQzsbb3dR1qhlUfkBUCIazBPu4qi3gATafM/aHcRLTEQAZYeTlM
Dh3HqQjTwg21ZSzIcAAgon9GDgIym2o1EbwW7dEwVXFvfyROTHRQbw+lMcLtcIQVsbrThSWO/u1j
uN/U2ddN/isDgOM1ockurxB0bYxXfDXXtW2AMtRjRilcXT+tdGHLqwzyzUM/XKUKJs9HFoSYI6Iq
HyYP5yMZuE3/dcUYqOOJG2HyBqzjexUnB5tjzjmca3pAtZ1+cvzNiVOfn2vb6TK5zSukL7qsQUqC
Brp6X5lud9F3Soa5eBspV6iGRJu2MUAmZP2veWVGplWaFiHKomkzuyJOWlcUgiB3gvSeEFymNbHi
g30bTZnwvwKqBVLWZLhoXf8OFGCBCNEeq2vXIqQR1g1AXRfcFLr6W+NQ6BFB61JO0Phh/Qx77E7V
TqOtbIZQQhg/p0MXjqUD7IvEpdQLoUG1mcsoToTipw48XVWnwjXsQny3/MhqFMIf1YG22qKe93Pv
A8TX077ogf002nesuRHoJHxBFovzaXiJwbFk5DAaZfZq9/o+cv9lm7V40faDxIkOrHmIju3JNy5B
RvEvf8FCh1xjAeE1tOljgGwDqrZY9g8Ub01HIjWE5wUESZgORpCZ7O42oQkhS/1IhmpsmPqkCZGb
XEjeVLEBgTpGALRiVK0zMmWnY6dg5TNgHRh4El7DfLwrQlYLfvfFa57IWjVeSGELCLmtLYJ8ecDz
hUy+AmmfPiQ1URAozZ+gn4UgU08XJPr/vDUU7jl65zM2oGp/0ntxKVJf7FrowO+OfOZd1W3dC+cB
JmYAdISl5FWjv4dFypE2DppZ8DYvALp8tEKxWSDVvV7js843D7VXw9jxxeymiWb/+qd00jRKe7/o
HcHBlqSzCDB1ui5IxGOCxjWN1WteSYV4WO4iuZtArwPVnVeId90Ec4U9Pq2s5TGqJQBl1b6h9IpL
jW/KA2lXACbtlZR2fpOypm1FzF7zoL5avW+RZl66BSiMPrT6rM99umORoBk7obzOBqaDrIuidXa1
mwao11/9kBKkYVA6c0gaxdnWYZT1e0FHS247TFP4ZtI3cdguH2sCRmZNDUQVJgJxu1Q5AZ/5lIqK
2TuPh3OHasVVsMvh+FibCS8+ZpbRG4SYAATEi1/IfFrh0C2sTU7LY59G0DB3Yzr82LL80dGAkjhE
gaIBZyrd9vmPrTLnKOeMEaw0V5bhStXg7zlb+lxyo+nWExDz7Ajp3EhKRUAJQ+60xJ6jXxK2e7Uw
f178wKDY6H7R+ENgSqTwcUgmH2ROSR6eaf9G/NUTzeNi+Y6R3BzMHQZJWjBtEPNRmHkjWoMUZEYx
XEsEUuixB5mqmYlrxsNYFSOhmAu1UohWOWNMZHtmRsokhaPOyRuZbbaE90vSt9lgy227uOfqOsLn
uKmSpGlRLZsBrb2+0b7f0H/G+0Jb1s2IaFa4WtUEDzE4SsHVYCcWFSzxzvja7iljEztCS0r+VPMw
ePQUBC7Jyip0VPEanSF7gmRMSF3WlUGUMaNs6wGqRBl7DSz2hJkPbAeFygF9WnEEdCEYlX3Ys799
LROlZGdetMvw5AodPIKKuMDzl6SVsBg5LJyfscJEjp9tl8ZRP5h+LhSGoSBos+Xo9nICfVYE2wyh
WzVOSVDAFUi6DnxZK3qLXTMNfF9bJO9mWexWbHG0w4SzaRTXCUCxIYnKuQ2FS3uj6yMlCRRBmSiP
ZU6GL6E1kHsWaQ6XwGMhbHWRr8nIkcBylNEjT8YtRnkidZqzb3/3Gdju6lQ+A4oVPmcG2dlZokA2
47iKX2BdB83+Rn0xMaohRTfrV/u905JCEKyl6mQhLYYmD+rBEZ2wfZdpDLLD9aaukYHEk7FwjzsB
vYaKNsfQO56DhjkMu6YyEriQAiIattx58F26CL6f29YS2YeGWXkUP5o6CopkSZr9neYDN0pcPcHv
fBobb5WUN8+SNMVfbPNn9r2aGqfgeQetbiEDv5MAUyx4vkCzvkiDDA46Z9nUCukwa5PkfNKu0imn
6hP+Nmwr+5WepSh2ZzoyFkcBzErF+XwO9kWRGmkZytiACuD4QNxvc7d0e2aNOD9k2iN5w1AkfdBv
LH5q7AcCyq2YhdXgo5Ep56q1s7rFNV7fqVVxYyhfuA3omQyea6VY0gxOGaS8UnBZtFv31O7WDNCF
4fRv4J1LxlsczekjG2dsutJz2UkgUS+uNa4ueqLegL1BVyjn2QZd3qgD2/9A1tk5s6DDoqzPKlRL
Fft6OD8S0nXR7jgWouf2GcKic0pY+rw41i7oas189G9/OjghdSvJGIsJz7s75coIH8tuAfqchSGd
ktPyc+1xQv1KBwBlqWVus2UbVF40Rs9IP7jfdyW68+vJo/hRiAD167sbIXdLK+9FNV4GQIXxeUef
MVeJBqGun38H+yx6zd9H8p9f7Q6V/0gv3wM81EzT9sG1OTlZUjqwmGZctndAC3jPLWQ5m0ctuiDL
M8tosX3JLINvkuG5vUDOxMaBcd66PqE47j0En09/Zz+tRKGx9B7qLcHAAcNEWDWAZjS2VtxQyvve
cpfUYmlaXwy1ouxhXyXLdF2/Sl6YJAW7+Tch+wSN/TfNgVF8j6F4S+zB/1sOyuArSrfhMfpStUhT
cIczdc+axx4dIJSrtyTRmh6N+o6P1K9ayNoIoav80yuF3juoHWNLQR5OP2RbFuumFEWSfswk0dKO
7QCalebktcufDDgTV9nnkqNc5dWItju2nJXLVTOnTCJe40TQEOX+SB+HRZmYLVqa+xm9H2u2+l8c
sHnciAWBs2vUYVdYVDL83yQ62hSkt7PDyo7il+tVmTxbppCnPpkT6HIWbhUBYtBksutlVMTyWJov
ri+PSG/PjGL/BlKtSVHRdDqp3KBtk/YhZp+e/aoztUhWcf4bGn900+SIgqE2c47p2k3XVAHr4XQR
vQ31ss7upUCO6x9IPYUiB+kgZvfc76Yky9zrZq9DpMexFR1gAOAwmxfdJ2YJwpVjvA0UJi5EV/WH
EaG5OarSFJKNls2iXevahRfrPC0b14MFvW/unc7JF/d39KfKih62fqmkQ+/+4JSlLXod34jQuQyK
5DyZT9klWoKyrdocA1ioHlJMwhVqyWxFJc98IYTNvPRWkiCIDXnIRbwWeLvO1h87SNLhJngF7F4U
6mbRGmWE01HrpEZpNavujP74uUPcCHix6yRQD1N9vHmf7+TCvXLZF1GlSU4SKEocP/9ZAcB+I4j3
7mtM2HIdosuOwSX5ej6Eb6kqNxLj6aIEPdkyiRuKMsR2p6SLNxN+WktrDHCKA43RROARlAGz0raY
Tm3GjEmBflebAd4pPMo3UcJlhNx8Sp15UdwcMdtDMkVddwU8PXWV/0WZCO+opshUAVOMAZn3gG56
IYnDDyrk5RwHZgqbGmhK1fDPSHMBkRPssiNjm7hzI2Ko/4mtK+W+vBEA7NlrjoA23ytU5ekPaB2Q
EVn4HuAyY5CxGHS2ges8Nm9Ym4SEUlFpieagCz+ZeB4NGu3/NxrvCzwWq/jWfG6BE6xhqnBPKWJn
5CjRAnWYChY9pMIkfBVkQZAPtPE1NqkYV+Gn2xEvXzDV/Yk2iQbGfV0eVx9FfuMRAnZALGHySF/X
6BmW1LkzcXid0sTKwTJPZA9IGPKn4JLQGbYrP880YIl9x6pQifFsOGJNHwAafg4xYRAoftbRiE+z
twaDAudGybU9JHT5HwkM3Qh+Kdp7EOkXj4YMleiQzHLcvevV33a26JU70QKAzj2C7tk+9cK2xjfF
RnOCIsjGvrakitDRv3UkSHWmpRnDc+tfdjmgHESG9xuoMOogRUuhH6dxf41decwS9gFxb5jioDlG
j6hrmEI2CWkSO0yvEzjLr4/7dkbee+OECG0hlBeQv/1CKVKfYGBglDxNBU0rPEHNtU3MoeBRQOX4
ahZOtSVn3+eeQSo13WbEPryThdKRbJZU4Jpy63nRYHLaJCD92ZgRB6o8s+A1ohk7M9FPXeVmP8er
ffi5XoAjzZ80FxWdEiDbY0/QFS0SyjkXnyCdbIhv/HlJ7oMCku8YJtHDqOyr26570/hKOYf3P0R0
EqVJVEja33KuKBH18n3pPfdiCpJ30aV3hLv6PmBuicdjOs6KUj9kiog5hgOknrdEHvAD27gdVyyS
L0UyYASMhR2xDz41ZeQt27YkvCLXs9HU+xOHF4nboJ2AoJk27MtyOXqjnT2hi9F/E71iOfz2HxPE
ZCTXQXOtDEfYOUni2p6TR5WCjEJUYZFDBIwj32tpwvLGe65Ef8MIoI2FGV+W+pVXLpTfoUL+tDWD
+H9UxfrQ8wF64Yv8WCHi4yL3ixfLw2b4V79LjSW5zwf6l0PvqjuGbPoTZ57PR5t8NP1u59trjhRd
DsWVftT1s5OiIBDvXmAZg5AcmDzcV4ksDueDUWJ243E9ZTcQScx13ti9tFzGBKfNeR9gEXssKUgx
aDzCma/vgd+Am4lSlltHhdgxSlAxt/EssKJoZDnADQeGtZ7bqDnkOXGgM7/aWbMJFYh0U8mjZ1I1
bBes7FoVUD/WgG74yt84ENd3r22+ElMwdgTm8NediVr/3Btwrt4jAiEPBs8wraqRNDRE0E38qdDt
1mws30a7pmTiU9gIZ8FwvX4p+n8DVexGOibhZqWDYm7Rr0Gw39p/FJCaxm7Cy3qhxMHdstfJcv3j
5OxFigf4loUQzbQlCUzbE86Io45nNlw1IKqowflFf/PmXmWWFcmaBv72t88e1samov+9TWzD3+SC
ULUaUun2KIhsqSlOL8Ky/Ogv9azVVOQjqk6m6MRoCyjS+hRASsf4gm+PIuv5vn99ecaZN15g/O1p
JjzrCo5kjHTnJiltzDSsPk3fYr3s7ZedbAcLPZHiyTXRdz/FG7yOB0FmeRdnfdZae+wXES0qZUkI
TX/VFmuNb/E+EAFF96xFo+uuvsJOSJWX0mbl4VInDTJZXVGOhDFcr4Oe4fwWk1ARHzvUistR8jWO
PCgnw2G4ZN+j3FucNzLaQl0ElhKu47EuDfahqfVmdPw/Yio1qHQlhSN6SEsd+3nnsGjv3C9AkW17
WIKI7360vggW6kcfbN6Gve73y3m+R8NkEy82fUVgyU/OSRjobT/We9HV1SEtjRXUG39v5MC71Ai0
GKaoXSfaCV3mBSrdZJPhncokBuUxqWCTD2B1udPYalivg8uq8Fbss4tkt4ncXj2X29CH+19H2/i9
N7k/DDNmRQhumiV+185XjTLel7M1OvnTycbhKZPnRuQerV+Jku9gpjuh0TNV3eL+mk/yRSkwXE1Q
F2MZt4a3P5YghRAe4Z0ZNSUFGGyxd6uED6X00FyW2th7jto6fGhPK6SqEaVZLgmoZOblz2QYoyZD
KxGAP/FDsQHurrvmSMP/21mC3Rzj6ovAZmeG7CfdJPjEV8l+9ikEdrVPvLrFh77DKwLfoxScTTWM
wvYIvqoxO6w9f+k3TDKj4+f/A+VIqZYAzr3fJgkGMEysn+9jMAp3bADDkN5gKy3f20oZ4gWmoYEy
p2JB+rBo5L2j3EZkCD6Z0SZg021U7xTHXX6j7dBOYdVP0Fkco46CsSVYPHDMNnn4tBjaI7pnn6XV
vpCr185I99hMjpiJHT8tCBxsHVRWeIIZW3yTFulM5hE4j7jAvob1QuAaD6vb8Pt/XNhWQVUfNgmL
kYRwR0CRS2V9HuBId3SRekRqubsehK7a/2AFC1jK/uBGg3YBnj5F0FOMY5d+pSUFzJIqsPFQakLC
8K2/EHiK7dfqGMc4qnxBwgWfhc8bcG4EihP5gCCvMb4tLrTEDGfADFXOYMi2uSD0Y6LFBCOU6Rz5
tehFP7mvQgxV+nwaK6lYMFPHdADqQeVW5hHsW4xb4LNKFk0yenA37+rNji/wBM3TAKNeW+NDaCg/
LVUAR1JB9goUTIMT18s9mqk6HV3nbGlxFFAjkuevnvY+XRX5nLlb1b7b+SoeNjxnv/m2TGP/VhKD
gE2gXZDpGAeSe1CdbizpxjeKut87efS/oK7SskkSpTMG0AaNpO3yri8SPS/QTeDoKEwRpwfR/YfT
+paK+vZc58vUqykA1eYeL9Cz51o1ONhpNbVP6A9A6fm1nnH8rz32NOklcnDP/cyA/qCs09dJiRG2
MDuV7P0wGFH4dv9k0wOJm9iS+FeN4zQMdwewkuaPwyXsHCIul7p+bBnsbQRh426HCywqZYArz2E6
itSQNRrf92Lf1bFyRAWVqojRYw1LZOf4bwAI3j96EGwNHdjT94iG4LEJlbq6bVEJBBd2hRpcDVnD
G4iwYtsJ9p2hoFYWNQFMHi5tY7AtKMIIltAmAvcXojiRaEQ9SHnhH4suHHNUzT+DyXG8Ob0+Z8ld
U7LrRSZtD+/gU9SizM7NzGZtQlKzzuWcRk6WSzgN4Obxfgez/LFgYIPYUdLrgP4UWSV8eSHJlVdT
zmYpXMvV4Ut6pbDjfkkTHBjX5iQ6h+Xj7gnMJCEjiRsvOc9szy1Ba5TEupzCqt+CwNNwpAvVz74G
J8lIKn2p3NgYS1IASHI7PmkeJalFKFxBIXyAp5LTHDvMODDflMronWO/lc9O6jMLiGblmYP8BVSb
7VWuKYw54q5+EUob71Uhu7HHmaJxze39Y4MkNEBwJ4RPzAqtALEvUGsxcuCx2BX1FFYrdM/wc8jR
obwqmzYiEn0iNjdcwZA+r4Oatak1O6L3SDRHH0emouF3RFBfAa5lmDhj/4mfl7xjqw==
`pragma protect end_protected
