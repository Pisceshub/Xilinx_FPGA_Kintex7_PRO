`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
BCC9rc/UvLO+60OKG37h+5K6XVw9+xBlmGSPNNtCyHiGBNAs7uE+P7kAaWn27GhAeEpR/kFMWCax
az/GVqBT8w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KqqDQUWeBjbeC5Do4n6RoTO+nx+zDp05oc3Bq7j9aHdTCyJc3x0fyRiN85/GGjrUv39QuhEX8Yfc
PQieFCLLhIDiLcaO3g03QeMtoC4gucQf/+wx8FMN+etUNIAKvGSpHcDF3sE+QU2wR0z9UkcquWwd
T7s+2xbq6nw9IgjIn20=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ArQFRYMFjfIqnM01+3BErkf89TR7vHqh8+aVuOpf4ehtdLgHJ/5eVLEiyKB8J8p19WP3coK1LCXX
zKhiKuxxeGtbGwfm+yWYlBx9ENRZgRCMJMCvUsDVN2so7XdAPwkjqSnh0W76/Lhaf+d+pvRWlgkW
9DQk2DdXzM4eoYWj8692SXfxs2GVr/LFsjE70VNgWii3g4b6hbt8arRzcBGb7WdSP01/Vrfupwes
wvc5UsRUnFw41z3BPXfnJG4S7TLMUaKkpXt4XkwlgjRwtf/TFvPay2nUHGQKbMhpn3k11OWjCVq/
je5H9c1eGYvQsLZXkrE0A7BXPj2zxOkaxG0eew==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D+ZRBE6u1yF80QejORI2YlK5RectTc5Hc3ZGgcNzOnHuwsKdRLXxgO2EwzuQORFrUAcI2O1GShfJ
cDaxaqcC2RUD7RA3O2LsbI/gqaNLWKfE2cPM5kyY4LL3UpWPM0Uo5ak/GypCYQ+UOf0Kv83mOrCw
gTGIytvAqr7oSLY9s9w5ayy04DJKSe0dAiinfq3BJ0yg/LnSWrLQBOBrA4Wdb3lM1weRawy6ucLs
RISAq5pL8KX5nYwI6yisEb3R/a68Gt9JyNzCGetfTfKa/ZmZFgr4Mj4aSY4hNGRM3OGia7fX8MI2
J9WLaNV+MP1mjqAewxP7QuQOtPQpJ7jXaieBRg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ntat/Y12i+xTz2OshnCjcnc8y9zrqQygo70X+7SJQZtc4rY0Zflni9gN8Z4mJ875xuUjX+lsIH9Q
3xBNfK+u4PKka3FGIKhp3P9okYAJ4aQHDoQHPys7ay3p9o+QjpDu+LoKsYOvKcQvSTT5h4JB/ADm
8cRL+CJAT0lnMoC1oD+FzJaGD6rbUe/m+ozDAZO3EXBxQhmIERbrgUps+YqPcCfIPBOirPKyo36x
gPacfOHCAyEnDGqsYlZ8/OKD+fUUWGYGW1h+tcsLksdUksFOzpwjaG/aylVqeGnpGGdju9YCZsxR
FTDPxHHSYbWz1IdEVen5mJ4AEFHyNM1FWcDu+w==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iooVi2sFmNJOwue8KHSUPRW3tf4tB3uu74gs8Z6LDvu2knYgcu9jq++JPYpGEqao7R4n5XlVPf2c
k4alUHvp6Q50up5xf2+TM6YAlKOh56q9Kx06TJnkavZHpzcVUxjTO8lhG7ZWXd4Gx6jTrcXay9Lh
hZnVvqIrYIf7F2M9BVU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TKJ0HbePLQGnDE6xQ2nS66ju3E7NpHUMIS0eN5TmIrTiavo1ur6LEw91l2unykROGHhJ6ADO8P3+
+vp5WK18tY3bqWh/q6bhiVRnEA2oMtztFhG2JpSy3iPMMzKWi7QDcZAMQdJjnf/G2+bGK0FCj+pn
IcyQWYXOLQCp2MP5UnYVxp/1/Rseo1YZ2mplACxSxS0C9v44JZ0uWfMD6EGmpBALrJusrcpykUXD
E/ZZoTwRUL3BWG4AsvhqsJUYITtSPAjRUg6DenJjWOgD37PK6P1nngWyf9Jjbs53XYO39akVpu/l
Uewa4cLxL6R5/kYVDFXX0OuYcl7BxOYxaBLIeQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7792)
`pragma protect data_block
eAOL/opCDzBH1z0QvPCIvO3t5YHaZnTDBeHrraC4no8/yN9Bq7ZNopu2QoqF0GfPaidzA1LDG9im
vCROkVXjqdGbyzqGi2E+kabhwuhyzWeNGaXeXnw9iCPccPclNjJAwiRS7WPApbZTI+Ge9wQgNya5
e2R6qkzqnh2cB8HLJ0ZKnt3PPtWE5dIdP1qsSRXOyCUI0dKFQLOAo5r38806PKEbMi2lVJ8AbdGn
QZdJKKDutf0UarHwbg+FAUT3AkRkevWY19lBcG7PQrfRP5X5mSzewVbhcdhxi+3t/VNKCSUh0bnw
PQOfYaEyCnfl2mBIxo7J6tnTAU3/2nRPOCP1e4fj6ve/IMKFV7ZhwRhXzgum2LjNQAap77fqVkbw
XCRnJsKxjGAFIOqVFvo7NoZXcWOaHlSB3gprhlmE1BPMPNnQKH5+OxaZJG7VeA6WgrriIvNKg8Us
3i0NLbw/cHgExF+vejKZegfy4ug0hRpED4b4YtSod4NvDHt+gUqmiZOoS0dJ9RnLcQVF80YjED9N
lnbNOGui722TLuoXUmdP758K5bKqUu3x7kgvJHackU7I46MWrrdTwHTooYDoP1GaO+CIPZV1ZK+K
S67svxDTcDLz9UiuOvrT7PjWS/w5DkleUkXanlDJlyh+BSTuIbZPof3ETSDdvpEf4hPX55oBxM6a
dpM2zDfWhT+lOaZoelPE0pfxiJqlsxyj9m3DZKuXI9dpya6K3sDPSchbhsNqpHiJlp1a2wAl7rfI
8LALl1gtSl17sukWQKsgXVr32um7HpyanW4qX3uKKG6EIymzF4cP5PsNOMexDg9OwT1I1+s4AQNp
WK5fJZBJsKVXbvMeAcW5czU4MULKHtBs0BQYsYSWSWLuZS/WHohWNZVIAuwekQOAxkuSsonpUNaV
pinFGs3K4rRxIW5GVooSeYKMhRKdiWSpcjOUsUouCA0wD1EFybE/4LuQF4cdiHKKd1ngv3iN+GYd
qC7A8kT+vNrT/7tQI3vASWRHg6x5b4Km69mmDHd+yuzJ7+FFOZJW2l3QmUbpYiPnPw7v/8K7MC5/
OhAjStByr8K69NCqrvYN7s39O9trOkRxQCqp/dYd/Yo+nLMXX6AgieMeg0KpAkzRDEaQhyD2P3ij
xjQlk9KYCkuqK5b5Tv0KDvFFt8eVZ4q819TnSvWEQz4yKENP2OaRZwzwvoUGl/w5JZsi9Ury2o69
HzxVu2EYBC+KwU6dTcujS2uHyKVr2oEeiyZhgrPn29Hor6LVRIbG5Vc/x7DV07VZfQIoTdf1C6WH
fE2AmjlQk2+Q8zyDmyYm62geahRwU8O1t9lx2OdBCOqGYC7FEiZGAy+NH3340n2znuBFiyYrXjuW
SNWTbULkJkzunzZrG8YGOmKBV4ySImyvkgkOEFLaYv3p1mOSF/aIvxNOcRU+ggffvVXP2oj4/sDx
2rCXcnkHTIXGY2CxzUg3ZW2HAkoLw4WBkB+nmkl7cyE4ufn9m+HDh7UrTJY6rdR4PvDkxfmHZBaS
gMXOANFAdLUUxhbh9r98o1PElaoW1O6xQmbNqSrE7bbG+cCbPQAW0ui4Yn6kxzr9aH1lH5OaaVaZ
910Ye1JFec/MqBipDe0oHAQeVAnnnPZheKnXn0GSRe/kHxCqUJDMoovXoq7ufVBWowALJhAkSUWd
KyoZeuKXEQMvOdBMuRQPDKTWbtnoP55zdGqjX+iXjwDvdY0qbwFOdZeeX+CuzS/awiHDuJY017sY
OkJhc//bi+v3fXS3YLkp4KFUEv77hSOGPL3RYAreWBWwazl9WLWhDwh6ErjGaIDnqp6YzLS9xUCb
Cwe3uESyP5H35w14WeFxsCaywI3o4H+UxDmrPHWEVbEdAu/t2D4ykYGGXleJ3emW3QnVoNZgubp7
BHhJLvyvT9qjoHBCUtjDHP9f5MHVYSJynjetrWfGJqludSV+EinHvSJuvyK5++tN+e/xqxdf4qBZ
hItgmzWyarWVkW83pOOu5Dd7kRd+HIZAKFCIYqPr7W75Pt9cL6SX4gQZH/bF+JTafd5hx0sAPmL6
A2AIiPYtajaugWj4QXmDKhgzPcrrTSpNPEax8ne+FJ1I5XfH4jEGv7AeNAVk+UGwuHg4EDh7peVn
JPSk5PvCw7as8zTu4nAb2pnTWvGlMTB5X+js1ckN3S/B0JTxuai7RAh/+33Bnf6rUXD/3eDJqDkY
9tz1PGeMxeC5tBMQRxpPM4Z6h/yawJv/uLu2d1Tg8vhe6Wq+W7ZJ9EHmMdhwAqYeck1J6D9sEc98
yAVGtc43vBb8dw7QeMN5cktPPgb0tj1LQlOb4u8JAAUCPHBN/RfJ+PEBh00SEAiJjrsuP9KvN25n
Yx+U2+cUj0nFartoYY6h3gNFlSH8MYdfDhMnK1+AbnsF8E8Cx+/ILCnt7bniyS4KzWM43awNOW4R
b/g0yvr00UX8oUG5NKP551hoqJ1Ix6+uZOsrnLhLLNXPPJtprhv1df3u7DoloyDNh84ZZMxmzWjo
4DmWVDeIC1DQKKCZ/V5hsQkC6d+W8n9xa4VFmkqFOk+bzpvG22WUMG5hzaSNEL0pmaQJArss6PLt
wuB8e/rvN3R1oEtLEuqvrahk5VwULulPgZcDF++6nY8dYWo+d9CwwpH0HVUELkkACbR6erHTJUD3
VzCqFjvshk9bpsBvhl64XI/3LgGnvHzE534iz5xwUlsVzoezVhdea7PeNMEys+o2HHPQtf47UUQD
UURx6c3G8A0nHnNtwd/rTjp69d2GkbiuW9K4WHH+dumoYBwI+KbydJKXOQBzNnb8ZgHEC5rmEFD/
fET2s5Q31qRqa9uCBk0LnTXorJI/AIX4YeVfhH+e7FvmwpJxdsCki0XcEucyV5YxtsEEtbd+t4G8
cOzCJpZm9FZCp+SjzNj6PY8N5IQ3hx34u2z1JYdDgn1uxPvcffysmT1hseh7ZrQaZKWtfquXcdzI
m7j8b9fKmX5F5pqeVAx/JZjs8cCKMPsU8bnHSGtyzbuDzdR1bKGP0IoTs98MUNHtIHLVjc87yRVX
foMHnEPnVeqcw/PEyavxIjXQFAFmQwxSIEaVgogax8TiVG5SkiGBvR5s37SfuDZpIicnuiMZcoK4
s05+tPLR2IUbxkUGIr6Hqw1QRactA/YsmjWw023qeTeejh5Vsw0+HziRB3XC2U7VfgWrB4rPMm86
8NpZMy7l3EclLBuiJsKx1Xfnfn47Ml5HIKkVw3UwibbPQ58HqoJuCxzBoelLQ4q+Azt4E5x7xiex
RbQd6rRB+zGNGLD03lBlK6mRg2mABP1FWCaea9Nj+sRIHQ1zPm3C17BvRjYR8r8e5pQgCYZ6HAu+
NGGUVmj6CHAz7J9sTt4wXSNFaQf+dm9yBFTv2kmpk7saVkLHLHoolCM1/lmlHHIGog9exTZxmYxz
mfT4kUIklcS0sO9Gi5Ekm48E9BN3dRJtS/f/+Vz/TJmlNv5wIWylNcCwkpZ7NFJDakO7CasHlTsv
oxWRC58bW5Jdr/BVpkOO+5Mo65bkQkkXAFg6GJ7Q9hRqpZtvhnNT10t0t5IQg8FaYtMXKGikD3C0
xCuzd9zRwRtLXMbQGMhstJRxEt73bm3WGdjgsHRE/UXX3eUg8/pihEjyKzRn7duVif2YfkyIq3qK
qjyaCk8uhh7jzhyOOI2KFv6SYQLUdxfw93xP91sSM92EzjNguxdl9JnNXFje65gSN9f/igonithe
mczAMKrkcunQpviKqWkIjVC4QpRh3X09KFifkEpSH32BvmbyzxdACvU1VJvnYJ7ffywmL965YmER
V0Dgxpj1uQf/9/po4ik/K+R8ANRe7QbTHgG+Bs6jBVk1MUY/JKAdblIMylHUVYNr+lHnggp1GklW
ugJG+kqEW7QnMj+z1007lOyiKh7XbkZPX5L9U4+g5ProWK0hzzlBmTgv2HUIXOjAFGv/emx3G6TK
2AZ522Bqlr22ntOQgLpXlOifQCG4rHoXdkEYqy0f/NxupIpjXGfiwc9xtmu2/MRdPgRNPGeIyWiF
z7zKoqcGUHo6UJ2cOpWmQQoUp3VZjMyshNIGZpVfZ9dPjqRhgLPhB/G7iPeoyy3FKIUyGHpuu+5g
MgCEATED/rfNMicd78ZE0Fyk5oWQYUVPqz7UuFRkT+oom9UmSdcB3ZYaYAH0cHnYtSQinMHXw/yT
TAlhn1NPhWpxvPjgEjcBfFUXqjjHBs+7BFH6LUWt4SsKEiY8qHRJbvX1F/jlqArvO+653/+VeP/C
G1XPc/s1pAW5ooEN6zvJ58WCqJY8UrT8yULqAUQLRiRQRFxiHFzCclagSfLLoOZc3Jifqs3FG4Vx
PhKezEIfwwRHDy2e1GzhngmhRyrtetR/FfxL7ubrSWtP9sg0+McnpWMAivEVxDlAUnDRQ94Nk95b
o8I/go/L9s+vlAn6IM1zv6cR9LquqPNQv3Yc3VIeeD75H3RQa0ZaxzyQrnH1ygILwzwnp3z++1A1
4A/RXHi47HbHzl1w0Zx7tJG3y6vZeWsuxiONOr6yYsKC1z/lDD30CRn2x8pZBIxvBhrM0T87XWpi
s7rxvzAokS30Wor1ocR556RnNL0oCxoBkpoCzWWsx7krWUENrtkrDbXkhxo4EbujHW7oZnMcZ78j
7xGZyVuEPxZdpyq/RGVC7WcRxrKQM89Ocm1y7jWx2clJ4tKwuJRvStb7c5ahNV2kf/wlDbLFLqDe
O+I1agPp0c9uDg3GLUGTbQZzR4y5QaEo+qrJfGBJjhi0zfh9SXtQoxHbkkQ+rpTai058b6XWM0zb
dIYrOylN+xjoa0s4RkLEX4CsNtZEhgZO/xFDUacO3n/gjObpa0C5aVgUg3cED6qbS15p8GW3s02P
67Z37WhD5q6647JA9Xa5CL3ucDtxh0yErzJOZLhr4m/ttuBTAQJhQxW/i3EJFGXG8Tt//loQNLG+
KK7rRouDaZnkASo6i1sY785htz4BwjAsf8tts4c/uRNDmaGZx+X2ds8Jtd+U3QTPrU9XH30qNil7
RXsx2GOvUEMDQIyj2l/av/jD+y0Y8ok1Idx8sJfgG5HkjGPJKpg99QYoGE6SuG1akgUUWLNOmhjJ
Gi2+x6+CPi/BHGmdjGhyT5BTMDEz8C1if/3numU73SC//l2YkAzBiyKEk+RwAWSLRn8reKht1IUC
kqXaE0wDCbgb1CMnCL9gsLoW2BRZvRzNQiVZmssYGgM+6oQwa6Y9V5VMvTyjEmMxDQtns/FM7cKf
awYamDE0urRTgOMBLkBvlUwL3kQOQ7qrifKJo0O9HMeEpSBPiUdUJyqjaJZl77kWBEQ7/PMo+/bL
JpnPUyvbcjseqV/BZaUx6uEmW62gCA9SnhVDvj3T+Zu7qH/C0oE8u9WkFw3x1XQaFK7Xptnx7hai
zWkROxCjmYJskJc4UldQDMXX+Q/CEXIckITg4ozBrHhAwIqta/hiKR1mKAZZzRcHZbjYVf9oenuM
n+/2kRyRmet+Sd8qfdq6h52OfJtUTU74EJftQEYXuE+Ig+1UCPLHNvA/rgPa5cKm/Cd8vsxTmvHl
WDeAoZJdksKOfdmSxzdrBywK1eBDuDyj3xvUWDhsetjd0vFy7EESD5GCvL6aoXA8Vi+nB+PWhD+J
YG9XOiwjr/shBVEjnlkfVNlx8yS72CsjYAN1dOFBmAV/7CsCtyP8dCXguOaK/pnK7QUIXPk9MRH5
wLdUi1Jzr9wEC5iCTfaOCy4EnJx7ME8gaaxPCXIXv2qjGiLfXo9bIdWj8N/VWB91ne/bicIqfz01
CnOX+0VEw79H07eKJLZXN3/nECx68yNExmqoQS/knvpqF/DghOOWQFNJ+56hlz8asM7wQRfuW0It
0H3qAguCanbGrLfNyhG35mDaCXA+CfRqdcDRgIS5Fz3Qh1bgs3vlJwTlo8TuCXaSBurwHwTIqKrQ
Twm7s8UiaTnMdqCrQG4T/k3+6oLIh9S0Et3QvFzz3txHHk9/kw2dMp5pDoi0BKPIWtanoFgSo2im
vrPfYKVKHGK+rPZK90LOqq5noEPFxma926kyuBxyAr0Lg+XlAaW48+MDzMNdxMvY8apWrgSb4IvC
Aa6saaDggrKeqZ1Sv2caWZ2pFAF1bE57eQqt8j6e1OmiuqwvecuqxmrWqh30V5MYXx8ZW5QE0uF3
XcWiJcA9oODtSZY//nfRR1QZQEs8IJktI62qW5WRXk7cil4FgOPh5mdTzbLhqvWbmQIonVdGUSex
37Tc+X14X4dRlz3MS1sQ19m4j0/ivqJpCkZa8QfZUYETRxR6h7yt9c3pUd7UsHSsdo9tIcTFFWUQ
L9H5bs6/OOtYcsHoF/8zrU6xlnzxmAas4CINB0gUXlG8gdU4AsSG8AD2ZwrqND6WZisvDYnMIAGs
T0FshdF5QfkY4lBu7FX0memuwT14RT6cs/NRhmHjNp0k1068j3wm0jwlJS7a3oHu61WIG5RsAz2r
QizjoHcOoPo6sQhj0FxIKr5pI7RKwDBQmWWcSMT4VrZkOmg1EWmF2UotUhR5nMN/+rMzo9PJo4BF
5ds5KLzH5xjcPoUiRs/NSKuEFYCTAsm+gtum5orIgc6aBqAmT8Hhu4DlM0hWeT83Vu+mwe64mD4n
v9+jH42eA96nMEGC+10pd71USTiLW/7eNNogzzXXK/eF5wfw5uBPdJmRQ2Db9Pj0cGqem5CRyf/i
T936dOImn+Mt4nIxMB9w8jdk/Bp8pyPi5r06Eoh4869poLYLvFbBPYZ+pwQZQ+gpS4B5qkuH0Wh3
eX5vrOXoA45PZGbUH/f5hyfRWAQ/t7o07OlZpRCmFyqpWxWlGungIlRntfegPJP1CgYPR3k/w3Q5
K35BSl9Z19fFN1sGvMT6DCNTkrzYq8WYwvHCtMDbLKzjabZFMHCpMNCuH7laKIcKVcrjtja287ux
A/OcAQSTnHIqZoM0wv0BBQTBuGBLZvzvEV51qFRvbZTYafLv4yvpVHmnKnKZUD6YqXu8qkAAotI0
ysO01Qv0iSJVKTzFvQYSbGhN2NR/KCBpdSxTSFNeYI0EQvOl3fiSZZ072vQZNAMtLWmnFCUdx3DV
2Vba2OX1TZ6wsLbC+o8joDapUgKzZm/AUmw/csWHJbZvMseQg8yVmFsW92BHC/ya2O7jnT6A53UM
K4+i43NY/4U8aUJqbUDa9XmOwIm3gzjO3bbEzE6C+tYAcCEG0r1WOjYhGRXDGOzlN94ZF3Im0TvB
s0Ael1DVTRMQlXwlIGPDRHOylt6kW4Wj8ALTDTlZvoACn/RDfDw1YIKJw4TU9KjDnV7WlSJqA4ES
ce/ensCrcmhWJqzH1uEhZzBkkEeCTOReQIetU30UTVk+hB51MY6uIi+9COxdeVJq8bwXdRRfUIkp
HjjJCPKpoNKh6Si+vExCGYVu2yui4vytODu6qjudljFSFRKBwzU3KpAieYAk87aUR/2i2x9jBry4
s0McmoCfTjI5tfy58zEqq3mJhKbmC7ZClF1XuGvMtV60Are3MMwoEccD+kvirI+dni9wbNorDpwh
JotYlBWs5nUpERc34+JEuL0KCTvwntT7OZF38sT3jxfykW3x0VB4/QsPbmm69V/5vdGu5KACJV9K
91qrnMxcozmU4/YkY2tQEJi5FzpbqCQ+0H6oUAyR/q9njCZswyXcYZBqn/X/Dk8+D4JtoiLWdALT
lGyXkCnzDnE9Ym4rqrIK06cSoo85VFap92JhTVzGaFcTzOsN4ff3H95cL9+KuHuU3caixdbZhsZb
bE8evbxtxEHrEJwdeXJR7SGzpc6RuZRSXklH1lCKxj/IK6PMDxorKpUsfkWFZdOPYuRU6FlhFiCG
o8IHRKkCO4lPof3eJyx4wCDsxc5bu9zqjZ3n8Wdelb3O0pHuhamhnNyZJsIJyFSex1qa6f1EQ3se
MdxFVZmjdpFbssxAs9Xt7ib6dkh/ZX+d3pPg1SgjnMY6oFkaqfj8Wm0jlZMAjXn0YfLn71FN0Lo/
W+llQeeHgePJcTPxtTQR4FnDh/zR08XRtfa+QZP4eVCHhcVSVRhf4nysEeo6+dzmU36Hh4vcGE6b
MPoNInkl4mFCv9D93KV+xeBhVz7Hb/5tOB9wEYjc+w8BWZuy9RzMz9/crgR36dg9TZuTVdEy1ycB
8oGfLSX6DyRgqJ48Fh68oOd4PrZlAQWP2oO3jnaCZ1CGFDExe5Wr8ZiKiUWCbKSApqHeUWMyMrTj
s2jVkThWTNcb4zGz1kFcELab62XzggQH9baacaW9QRu3FgU8pdcw9OAr54Fthd1UIvVdn1IS4SGa
8KXU/NPdp5TptnOVgvgSbTqjKo66cfJ2EEBr5PMb23dx1bi0hyD3v6169ygHsOUmtBWCAEKSub3d
yNwLLfO7DdHEiy5jGGAyNRv5DKXOz92T6om763N3zyjH94Xs6YWjIxhvcb9RXlmvg/5we9PGQBi4
LnP6WPU/L0oAyL5zPNxGaEcmUCPrFU4wKX8uhbyKEfcHlS9lffzEp8YUW5hmIG9JTmp56Oqydjur
CO+HsJyk91X7mxAHVSGS8aNeJlChr4FXZPLQG9DnHRcL1rYQKqBOP60jf/upN2LcL4rTPWdPvbnn
YTY1NsPZYocLht07yyZNfZTSM12xK9iW5G8VmeSc60meMIyQRg0IUxVYnHMFYAGXDGGXYEDXA6RO
qMCxYId/Lxns4DHs3keET2X0oaAKVzo6jsXhuHx9SMouQXfjajgY8oTrS3UVn0GHbfJz977zrRW5
LNFU4t6Inc9flH6NHpXEymF8bYkGdlr65Tnhd5179F3B1dD2IxZnXKR4+8OadVT03OAKoMc69hz2
AINFrlZ8bSDq7DngFh3pckA5vaFh4WZZLm+ywsId4E9vA7y0SSPI5H86NRfi6iXg5w48W7qU2zLu
ORf80H14EL8m6b+TJlwoxozsi1NqSfD+du5s+OZhOj+pdW5neI+H5XXwQArILL+m/LMrD/0aUJxL
l9mZ5C2Gx5syXz0ahXsGnAo14GxBZkh4rOgdBERXGLmp1E6+GXHT0/EPSGnP0M4SguZgkbTKaJ9x
tNDJYKR2IvFSa13dy0IHPhzuj6ZXIRHil7+vbwrBEnaaLP8kgmqnPyZiOwEgb1+Q8PzGJ2weTtNp
ZA5Q+31KeXGrjRfBJQOukDV6rQFEcQWNTVttpXSAZVRNX8+Nmz6Bo4/VFWzfKPmAvmyl+gmiDHS8
ohwWzCLF0ceQLXZK6hEsUjn22LTC8XmefQ9Zgu9a+yaNDAgvWUH4YlBXc5J0fDEvEJsVYmByfKiw
WOxh6b/vzyv12yXwd/V/ad+KAaRzRSz+d4TBcZkfceB2uj0T6G4HQGqAiWpmcWLp/YjPzFVbfcjZ
wQm78/RO6l5a6tC6CfeKda1jTBWIWwF0t5dsBdChVC6A1B6hLxm6HaQVgRvWzKFMYJQg/ytx3BrG
6RDbXgmSyEqVcIOcpKZ+HbKT0cxnd8Esk2M3LwjO7fzaneID8w6QGQZZto64IjDefv5aXNNKnS83
PxsjGZakKtw3aMLwvuc0uVTXJPG9NIlPt3JWjZOkt9MjJGki3vrzRUM+FHE7VCwTIm+1N1BsRLcs
zbKAqNjSh2kDrluJfY39dIl3IbaViFq9Bp9wynNCw9OXlB/5R4MKzJJCjPlBrY5l3EhAJ5LTAetq
rgkDcCIJ7YpKdLPbe0hd3nTjJdxyfodkz4YevA2ua5MbzbNziqT9rr3uNR8jKoI18OYO1x0lxlX8
gyxKI1llQTUjujSRmQoEO8UMPm2TCUdd8lCIxCq3PXqRttvER5iO+eV5T/LX4UelQCETqDdCTW4h
08ev1PDlwiLWZ3eJkhaSDGMDYcKZfAoXXau6jT54Ol4Zoq/Yf+qbUEOKj/pLoP/wG2hRR6xF8MS9
mU6H7QWZqcdEfM+agJDinxktTkzJ3ISm7Ys/pOOEnbPZ1mYu/K/bjLQm3FJ9ev7LIXCJVDUKV4wv
2tORNR7adP0kCjArGS2Xv8ugmMmMWtLo133rS1PYh/9Q9gv7j8vgZa184PdKwDMK0r50HCRn0eyn
dd5krXJyqPdJcVVPNL7dQMUrF02kDBk8DbaqihvSvhrqDm3xI3LnraPeUYDFw790++RWHKnwSoem
vu8k+kVY/kKljBBhvzk7rNRkgYbKNigZmUbaVq2atjZtKz60B+FFOWuN1x5eqQLaae0XzX9ED6zE
RwybmnJDEy2fJ0TdWhCrgqsEggfPcgWLFACdNXDBr+TBZCo12gl48Lzd6ITdyFP8oTE0+Y9rNETz
BVKsaz0oUrHkeBF7TCR10kOvvN1GEUt3zxhsUO/bDVNhYZ6ZCBDoRKXHm2OTjDJ0ec7e8TeFQ8Yp
f0pmu0a88g1R365ZK7WyLGT6P/QJ5O8E/5me8X2EYu0FJF7LcORRrA==
`pragma protect end_protected
