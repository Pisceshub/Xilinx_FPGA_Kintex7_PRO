`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17696)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEF+6B9v0ZnnQiHwZSLKOS/Hj9Np+Be6FU2Zld2edfkGmxSQfD5buG2px
mUFh6G14SJnevXdlrOgyXKRQ+vA6MieCCI6lx2qaNtLBKZyrrBgVn6QL2cMA9S6vn4SUDJNpR2jt
7DAnBQJDRxMURuZe4gSaLExqjyBbsoXSIxkbXhTjLuo0jvC1UTh4Y0Odc5vygWkEJYsJs8zvm/Ik
MX59FjNUCs+DZ2qb44J01va521p2zHcQ49uwISuYFg5IdnwXjgg0LMwgwhtacmGpDc5tU26lbEWb
xlm6jBRE3YPFtwj7cmrmilewVNDWcJxR9dsInPHGIweXQ8UPUWUC7mxV1jTCcV77fzrLCa1+uttz
7qSH58VWHLwBGs9IaD5RTKbVo/TWs9i1xMHscxvMhS+sHGoSKqYK7orQ6TRY0QvSVrI9IBkSIFh7
AcTmDU5dwTaJkpLObrZfRZB7923101GIlo2bqcr9iGx+A6KcVHuhUL7Xud4LA48hG51P6CBosngO
iyeGxvNtm9AH+KTdVnXvHMEPFKeQh82g7W6EQGJrm/9Tp5q1+0NnPX+s7UeeRaQLiQmkeMEm1H0a
ey3b1z5YqTGQhoib5bjCfmE4oN+w53awG3nExRjXNjN+RNG3rBn4jS5wzz+SYgyAVHcVZHK5KmGT
VkNCT/aEHK4eTtVx/Z+T8K1hPR9FF3yZej1gkrsiulgqQ1RjXpcsfpynzbYMVfLavOlrZj3CLFFp
WWqKvMP1U1vjKEC6ilNw469vB1ZE1cfEqNIuYgR/hnJLBtLGMfX4i2HVw0y1TdOOB+AbWYYngMPw
qVVY7ljOtjCnm3p0sGc6g7fBt9j147KACaKhZc5hYZlxJHcrAbRvXQiYxStbjm1Q8kXKaC8G14E7
9qcQ2Bcpmq0TqKkYXaN1V17OhCv5qvyN6kncfeu+jO8Yw+cUshPeimLoU2XOXxonBeCi/8koeUiq
0mP97UC605Mqb2sjMHFkc/fjMW4PMzSXRNqe9Bt4mzWDDJXdJBXMs2JTQPfK8OufEUnwUSokq/1w
00AzGyoLG3IBd1OcfkvL+VF39cWudBiJO5k5b8d1u2dTqWKpZtR/tX9Ox7QIyCGGNI+jeypcsqj4
aS86vf4q9PllmKr/fjhVScCUHkxTQ4E3qPwwZEYyQo9oBOUAe18/uh1Z8OkakB414Yd2OgwzNE8Q
KNDk2GXSi5EQWlWbJa3i5BVg8hNWbKYA9aVw7jzzet9Fmcol8Q6SjDl5oeMlZBJ5Wfz9NFroRrIo
ltlAmOSTftCUxSmzO8s70fdz20L/aBaG/gHqVi+NV8OUHpONfe+liBUEXA5g7OySFYy5xoDsuTlO
K3up5LRfUKEKPujt1uTIo9TsXrpwlswXAH6PRnN2oGCy/plwUUPeMigr/tAUjGd17UUqehyHQ/kG
1RlE/enEPVWPd63ADc55wZAOxVaJ2mlvIeVPCZbyeHk21vWG8tcE9K8x/2RWrTTO/+uL4AcfcWEA
cdVUiOxcSh5SK3/71u5bbAEMifTqJlhvpC8SLgx8J6mIA9+7x33D2MrCaRimKzgbqj/gFPBnVFbH
f1bbNdeouiX0JTvD6o9TZFy4Z8lVvriaCkVH8bqp4n6lSmgqm3OiMcWc8S4bu2y79g4zfzte6BaA
cpGHJCpC13/yTfrNMJYvxEr+FCHD4X4bmT4bKfD//W+KemxtM3PryI5pabcVODnHk7mY3TXCVd9L
HHFFNQOJMOh78VQc2P8CZAyNJdhyI4vHESQNhey10IrL016OjHaxpuQxoco4mSv7KNwt7PUOS5HM
BVdzxQ3vKUuFx4R+qMrhhewwd8fQF9IXdz81Vo2EnhqZ4vOQ9sm8rwLD+JYbzS1xC0YrYEQl2+Un
w11bLRbBsxSkU4TT5275Wm19vExwIxV+mBZeVp0O+kzGLNWn3HhOrDyEVrw3uRxTAqmIbr5JiMHB
OduYEpC3bbaNW7/E4DCwJ9YK5jEUp42SUNCdI9yHTBbECR5Fnilfj7n9hT/9KamlDPqLGb3Zl0su
knO0ffnSRXUdQ8LyWXpI28+dQFhpFJtVDGEkhamlERBepmRwvgy7WIiBIr/BsihLX83epRKtsj4u
9pqhABFJzI9HXHBYhWLNEa11H8maF7He/YVr9aDiVd+1obDpYZ8MTboRcgPvzfKBFuTnFRmfYNdM
D1AWt0FOdcL+giXJIKNsR/8LkH/RDgpMTN4+UwkaPLRJfauHhsY1RBTWulEeIYM/KcqrPSqWe962
QhSbQrvKerEuzWcidxAThhy5b2p8LxEJ2OwAVfeVPUFxlMXYtid4S1nTTt771ukDf1Hdos/RsNND
ATUFwQqyeEXEfpK4984Yd2HedbPljB/mUsBsNidmp1NcjOFi6WPhP6yGJKS9oRU+72KONu6f8tMr
A/vCa2aqCCddrFpSKJJ8PWyKjhBkvFVEcbyaBrF2UbGnMrwVHRNUn/FMssU7TipzU8pTkdQXIF62
t2vx1MdzozltXlSr1f53Kqc3p6iDz8OxnkNrpf6BH659ooccMaApDdZ5JQ8v6w8SPup0nE1kJBjG
YyaicR3TlkxX+TFtGTdNZumjHJFUbgRs56BBMb8J+h+fRgcd531PH2Ezk9djhlJHQeaejzChPDDS
hkmLwWAknoj4/Z4PROu0X+rBNVRwKOCWolOafUviIAsP6efXHdMOu+2AxGoG0Ra5bnHCLXwxgmuS
L5InA2C8WttUJLqfBSIYjmXk7UqvUZkf/LnE9POobAggFxw/dODu6F849geh4A1MbQ3RRNU6V38j
5u7Cqh3rj5jTlfsxSq5MAs71jTVrQwKq907DGbAE321xC6e8rIXEVgrNKt6REu8vjYKmnR0yW3dz
w4tDdpVOG8oUjmekbF05XrDcZUePfx8ET4ZTDYr8U7kYpx9135Zb/umskBcz+mOYBYA2w48oROUw
/av/rf91dN5k+iStQ3ntBK0qfwL38YFSdhgydNOLVvt7bYB9pGpVpmSIyGYRwfcIqaWxrC2HDH6G
b6iILzJ51FXAKHjwv7RfoRvtJR24kOOB5rCoblAVm4pKbzZVKIB9QKLvhiX1VBtnj0moNrfFAi58
7HgUUv3+0fSczAP/jnFJZlFd+yc6Dto5i1YPAPbhZDQrrKV6GHMqFsRUs8vYvwyVhnsqEulGCq7x
AH60CCjNilCKQ3/0pKi3EbpZQVMyTinRQ00QtqyR7PlyM8XA5oU/1p585+UIQIzOucVavHG+N9PE
GFXIlispPTsYqtLAY0xH/+nWMB+c4grVRZ8glIJsAihW2t1SrzqnqzfkYk8QEp3eLvgB4l8RBQOR
DNZaI1iFASp8PCAHQtOanlrvejpPQjx5UMr8fVXwzOw/5l+QInDNYw2IJw1HF/unhO7yxm14LT+C
MaUDlksA+3xLVhqvJ4iXj4u04eVGwKIdYplPHRipwYkGDL8G1D+AlwkVZlpiAiFV++M4P1mbdIf+
CPsFVSWFLV9PPzxNnsZDcDbPqsZaaSOymZYwBk7fvePcOxK373A6ySNjoxOAqTaJ1N8MQ/muy05d
JS5MJ893nVG6qAG8IyPA64XVAxi6PIOsMUEQeLxGMHqmEna4vaIyBMl+e3dNj0R6ELywguZDoGjE
g228nZNN7YIiI11J667plnyGEuSN0+zbZxeGzSjLuNkqvfjnRDDLsHcudyI63NyHjwt8RWI8t6cR
bBG2aEhiB50bSpP4hhmmEscxNaroswgXVFIK9lnD90YLzWXI89I1JYCWwQw+BagHTALPmDwUacR6
66fESFBLiAOce4ngI19fGJTFDK22hzNKrwvctK7HeJasFfYURBcnddz8GG/LTjnELK6suQOdAzR7
7Cr9cq4vTS6i1ccA2pQ1emIAao0+5lRf9mTKt9hZczXboPyiAiKFVjvVeJNaG4nGRtZMvRCKvbqp
ZCK/vHDLk77gd2p2FPSUNTcbTfeg+SxmLwqcRdvUHhvYH1LOITtKm5AqyM/xmkz7ea9BCjdAGl7L
h90sykSK/Q5JJ1nYpFpC10AxIODn5OXt8jGtf7ovjtrj4JPVUGWrjGjEMvCcyP0KeJOXdnf8v2Vr
2a/xtFIqehtg+5r++VEE3Avm83sUs4xgL/gQ/CHN9YZgWDu17dWfBfyW0WyIua0Ea3cuJAs9Mj+g
yFqBsseKqFp2Bfars3ETYGSL/5+0yvxel5RYf44+lKqn7RG0FffiI0Nl50PRvih++pjJtE1GqgVB
SL5aIzBvdqZhRVfWOa3wR49QPvKP6vB7/HUbzUwifVcEFJQc9H0TlsOuSn87HuiaYj4RBklFbrIu
pCiTU1cAELQwq87xDjxdTkeatZbOKGlcYvYYba9gvVw1xsuzKdv0NL22jEtclOAfmgbXJ8ad7mkM
HZpLpdls3AbnBilZCHexAWWMgQDlECf5XViVAe9ewhZ18WMPYbHOP0cSoruC0SVzlP8NpSeS1n36
ukC4CmiXUK3Ox7H741xS7PJibLDBV41P4aFkPqb6G/N0LSjE02MGpH5D/1yHoVX4MKAyBJ0QFUIN
osk74GpJQSHr4YkcjjnwW/kmrCSnWp2P2I0DdPLQT6TDVRTIxaqpS6kphX3jgbEFx+HsFXLAFp8U
KHrlddZSByiJqkspvgtb6KdjF3Ieow2ZL1iOG4N0q8zStCKOdKznuO2lq5N1K+GdwSuNlI2Dmc7t
gvpUxts4yYLiMGbXHyt7vE5NKZT4jax59WauVUM8qeaE6BRtSEQvZbN1TjWbM94d9/qF+A4Uw8s4
jaCqQYn0DSl/+DJmik8nYOiG+o/lyIivgDA6zDtL3W1u+pXLXfDrIzeCLN0cFdawkCro2FJpbLqZ
NDla1aQaitDQ7cWqDmLYI9LjhG9DWwV5fNj/bI8B+8+DUduLmIeerMaR/hs2+nP+EpPjKRzPxjqd
TTjiVYQDcg/F1uP5NiH0bJOgQQSaBzyHBf0oAiUNn0eLSpUuat2YqXnNIqLENSuK3Gk09gzf35cC
Fqsqiflnsut+ktgVfb5MBHhyXmHgXMgPfmAN0VNoaJD8uEuN9fzFNVbwbtgezCvgHt9jVSnpsKdo
HMOIsdzZ0ZnSBCUN9E697IbaMcp56N7ZYcarJac3g1afqvP46T5ov9jwF0SG23l0TnzHZd81Z+YU
+ZGct+1rSrHt24fAofk9I13husTFRqK8HIrTtPd0eG93iE4dti5L3yeduvzAqpIk/XjmIlE4ZRnu
N+sQwy5vIoQjEy099S/R0uq9JfyI8I4O73spG2lu6zqAyWLiXwcNj4U82kxiX84BrqB/aqPR9pEO
3ZruyeLdvQ5qklKPbTRuJOkRTYscryHMBhY5RMMnOkdf2cl9OPAKTdFlvOlTtAbzOkNVV9iD4y6x
vFpkHXA01zp3BvsmjwC5BT0Sd8FrM0sM1N68GG7q5xQHPhY/1p+ceA5SCDWPcztZlgsGJIV79dDn
NXz1qrPiqsoib7aYS2lfX2bBGybn3CL4/LqMW9rK02s8FsiFTxk8h42eGhYcdYYTPB+qbUD3Wb5M
VFMP5P1Ou8/sGdm7Y5DFF2DnE7dBAkTTq9/91aupKOxAxG3vf+kOgxwTpUfK8nT1jfWQEOPW5dod
Efqmk/1FeSUSaR0asOyZn3/BZtlL/Lz2f9yvHmZoLM+Bw9SbejfNN3K3f0nK+E/x1ES8DcEYOm+a
INomlp39zbasMgUUYvP70ckAhjUrHOVF14c2hPUmkVZtdWPf/yMQTU4fA1rxK6CfsVkyU4LxgOP1
VibRMrO/n2yuWwt4W8aP0BWRCPjbH1p8UFPHAqu8jValCWMIpYjS5FN/v2lKgDAd2+T/OvRG14i7
dJZAAvinwNnpD7bnO1Jl7TPAVflecNMAIfZuZlCyCR+oero0y5nXHvwRudWQif3QROygWWdoHWtX
UULNel67CEHxNIshoIxhRKGBnl7/+o7BiH/+JgGQ4D2brpD3djNAuHscb+fM7awaKM7L/sbpSx5P
AB78gv9qBMixwWF5tHLmUoiiU9iXpG8RpLuDVs7nqAmA32GIczJ9wAE01HT2OjpX0UQL+IZBBSlU
ayMkFvSwDLgysLyyzEJ2YELKoDGGkq1gkf6cQDlOPlgVHHtF+tC0H3je5Azkx9259rWmKqEbAVM5
3U1j4D1eIKZ4MFEHTadKfFswW9VtdzxtfWarnAgSU8/V7E3VkYzLKEW0WpicrRv5d50kqE+GiEbH
Wp1vLy+okDqZPAT9efKeAhc0kltTm1SWl2dyvBJIEcbFF+DA0C5IAlp0rsV9XmaeBEGm9vg993WV
zy+IACwDyW2CcRWcEFLv/c6W0g7OTVXuiGcAjyK+9h4ibqlmDb0Q7U9QDABzdxQ5EIZi5BJhDzRl
Ou5fHKXc7HhCbgoQM8YEnO07PZ2UA8nX7w/cs4/CUoxSZ71VDyBJnfyiRzTSQVQGicQnTs5Uabk8
m5K3x3Fid+2DDFoWqwd7gt8d06Rl82IBxWaGt+mfbrZwG+Fu8cX5Eb+rmswebOU1G4LVLLRiDi/V
r+STuk/tWfEfPBV7u9D0WA/bXY+P2/UR8lOubsAlBIaZM9fjbCx+CdLl6Sr48znK2T3YARrbvnTx
QgQy52ea++uOX4djxIOIZWZTpgZebym+61PtkfhOGX3puLhsJ86qXmVB/J/iaHwKcg//d4PeYol1
HLQU+hUlcRVo41f/uEh+uX9RksSdGUlnwhLe6h9S/1ogUiJOBByo3Q+paOYeLPPeu7K+ltJBGasH
9pL+FWtEgmfaoeIGJDv9WqdPeqgalsWQqzvPgsV++L04jzOxrf2NNsXHHesYa1oJip1kMdplEl9o
+0LF0722i9ie2I868GcSOwxaoR8vTj9iitx+/3UJ3qie8mGi/w195KcSBJJtTq1wumWuZ2Mqcn64
km7ZHoi4XiGA5ov/1A3XbLyQywDHQje21IO8iVm6aoSe4dbHCGwbsU7zzDE4jjnOfN31G4YaqPJT
fW077naZCRxUCfdogMqhtbQ3+fT2kyMlT7FbqrmigNROHmabhUHXJkQ2XDS/AuflFuRRWJBYFlXU
iO7lOJfmCcCt9seKCW9rQ0xA488bLHAQVuVa+lK26YPTanKJ5HWQvCf5BYDGcM5C/hJWT9iaMILv
jp/lJedZdCf4cO9ZNl6WwVlHxB0+kHKOXgktqfRnk1zEh5Th0bXnHNIl2nxKFxAU3o8cUk6v7ycH
NM871qQmV5dAl8DO2R5qdVztZqWHf5per0ar6NDa/Rw4NENUIce8PP/UJWk7zhL4UDYqZM8Kd8HU
Q2SU93tJQWXqIzzZDI/koFHZM1Oz4bYwk2LIXQJWsIEPEWyLykQgPFIJHiuBrYveMTS77m8VRpoM
AX9cete8ARQWR8gn1/0zAqlNKJIMvWJqKuOzNY0pdhgtH9HETqvoKCW+1pm29id/qhza/7Ek4ktp
OpdYocstpyjpPdcGOyDSISYI/3HKlXfXof36ZiuqT6ckrQaaANn6VVrX3IYMDaCj9NHScxwEsAI8
EbzBmQjfIPBbE2YNFCFqzWJn/McJ/EDWeexkJnrzjxZ6LHg0I1gbx7SdQYGjULJHUNC4qHQ0A8/r
+sAogiJg5QqsE7EovFwAVomKAH63muxDWEW3ytJ52EP0SsM/45ILTmnvjc+1LbsrbAywWhYzhQCE
d5vDRrSKE27vZdSq08KkiQg8cvfQVZ3lO57ZAhtoJhd1wk2glBsqnA+0TH1/uVonpGSWHlO2hCyN
oxbyaEQFEHFbq7JH9FcfxkGaATySoEA2TLmusmNx3y0Ji9MJBNMe3PndeSfNXH9DJfiW6Qd0Vvfk
stGMGhIPj4h4rsGXQOMpLljNanCQYAsHYXgMKp/9ZNxuoWr4vkjxBwyQJn+umDO5/Ut6QNc1I1We
AWjcNLsGxIstSVC9ynisVUImCYpL/pc6wncdHdljyZZP3bIgP5T2TX4wC4+45IuiC0+k5s34uq7n
mJTarru3yFlSbktn6Vla2Rde9ONPW7dJnYW6qSDL0b9WrP4/nLSbuz1xY5NE+imunNnov782QJlI
TM1GRc2JaORlCCDGn+va4GgD8Mr3t9Vbp6ubLsHIFk0kYVFZQfZMZg2nOZQNtGeMblHWwFSB4TF3
KNdi3lMMP+0pzspbJbdOt5UFKkXFLAQYadbfMU/SuNr1KiAXWu+U7T/oSDng4D6TMGKqRCGQwV7y
LhtTQcE9sB5bX0S6UdQcMgy894+bQ+MlW7Y0IGFyf74A9b8sExQpLVYmsizL8Y7+BBh/ncOj60sJ
SwWV8VmpEj5Y0T7GnWRctuFKowmv65Ecbg5X/TtCq1iiNk0uSZOdFjkbj8116lyvJl7Sigcww3g3
D7QIm5LwAxiTwkoEfJgiaWy7nUxo2P/Muwh6TBm/VFMOs1VOd1cYwo3dHsYKtR1XnrNVjHrKHsUd
MU4FH0RnX9hCHlQAY8M6U41bQSzC0qIsCS45BctE/BeYXowbrdyWoekVc0AkeLeajOrur/4ggJvy
v3P1iheSWgx3Lyu7fbQZy+EO69pSYsSbu091q9COfKoMQcoGUckqv6bNU5GqVIRMGKppomeW3Plt
FrLFKB1QIuG46rEsirrZGNi27kocYXMnHevLDhZutEp37OQV+310E5WNjW9mSDj6BiDLl4TsJcOw
naDNC4RJzWI0rv3rQth4CtMRjFRhOWxJuRo9CWRwH8FoN0tlO0nddfZNlWZp4qAgRhL/yfv9qoqV
vn4ytXrMXFAZu27WTjf9RpMMIorClRXFsNw7IiNbi2proH97sTg55mKSY57lmS/fK0mhhZW4PM3v
XMKYdSfQ7t1SxQyFyo/eZ5E3p1mKCgX6HwAMUnsRxAuiqvAc2/c6bZdZLIdVjF8ubMFVmjTQmdos
gaTs11bb95BdaN0rBNfoBt8gVF2cY2sXM3ukAQtkvcdS7V159mJCdyFJimw13bZIdkuAmQKzkEMq
oyTLoUes8PpI6TfI9eOfphSwOautWQM4hjn32gdUlGuFuqjxwTNpsV+aK383gUIi3e4z/M50hjcw
keedzLo88BYCRuvj+/rvxa2CDsJeWVFZ7RaFahWQQvz/psKKO/gksl/Gh3EJsVgoLcMOduLzgxfg
dGQTBpedpsRBwdDI59vimFd3O7MKNiG/QyyDwiAYBU6Qi09A6bxGDZOORUj/SUC1myso+kVz0zGr
36sYZxvVmHa62nOukGRTG9jOccAffYZ40ZB5MEsrBa0DANCpuuxcPhsJFBVAFHotxO1lFlfv09Nm
RbLz2sTlxj4CeybprEbB+GjjtyoFdJdk5xhzHgkooY/pSpSlL8hgjADhiXmxmR5DcgO+2PEX66k8
ghn8Pz4qLcYOVBNx1VTAN/bgZY5k4jRWZk3K1+d2spj7do1Fp21pcUrivYKvRG2Ql8ROh4px6lfk
MzIFl6WdylquC9AI9V/EKIXX3o9Iw2y9OzoTeh/KZPnDPZ3XkkB3YKh3S5Z2CUVLJpw8SX23D9Ep
WHewGrtnF60EdQpbWi3wHZf02ZORePckPc0xwCUHCaYEu+eZPcalJ506qFsEUA9EWbGJ0fr86ikA
hjHCabvXHr7cnU0IdqCmIuOynfiNZEKouPVKsyDEGqrgNz6zeL/FQR5qiZ6AsMZC4pGiYLuoV43B
BIIVt+fl6ZZXX1rTqzenXUE2RUyRHXVXK9ZQUF+u1KxPGw+wqlgjV6SyQAzrmjtd7z6B0Z6f8s7L
PdJQpRnHC0rY8DT8KR+jH+A1GQ/noLwbTQ1s0UR4Ta2XrvR3N245ftSbB981X+Q+TQeJw7POXBLj
JyFqxwR0ITQP66dCCQuAMT7UZZK/z1gPtINnK8AnUmInZCtuYz0ZzFUrKt33qZtjpKtxTNnqGdHf
0ZUSkGRkVFtHDHpD6qbglDsFQZV1hgqlvcqzAuT7hEoui53Jfb6RHyPKPH3WtX1QBWwjHQx/h3cX
8zx2ZNTyryUruBDl7aywgTUhYXb5a03fJ8CLJbqCuYFMdncCcig+n22G5SZ6/b9idhIOZSwSIrBO
vpe+SfQYl2p1f2UCxmkEDdb24AuU5W2Cg0yInGA/xGs+Yz7smUXze7c2UUPc5F2mIbyln8HBTfeT
nh56+V1w+vK7zI0F0a21+szvEUUNa9HWiX9Kd34lHEuelg2/mcupNfGFLJ0gzBJtB5JYJflQqKXt
3DHB8zInRAoLMIKMV24aGKKI/wNvjYqjnN+oW49m2YrVXrJMh7Uqu34csYkWsl1Wofe2RTmkzkrS
wtAT5UiDvlUckXQvwKYs+uSJd2SnakzsN6Q4rUyTZyx7i6QVQl4T2WcPEnlDjKJ/YS4Wtc3i5m7O
/z7TP5FRmTjGTFaiQECTGSCTkWLpfEGpWUfdAjzIVi5C6EOR5MG57Bv6R3fGJ3FQKescVD64eO5c
gS226JFPIGkwRhWllMq+FSxfkK6gBWePY0KyGVpntGn4H1bkHKAb6/jtKLbV0kJpraAatH3B3/RZ
oP8IOX/9O098JaLCwQkpaFoKZBvK2dInCYO2SVgkc+VqZJKbsLylrHfaZ9RY1+o75ya30Syh/RsP
L280N9lGvST+RI5dPQF6haF5ZduHw2v/YVuMsuirlOvUlBHut76Z7N7z3ZLJRa9VskuYx36OtWB+
JKp/9v+2PH5hezI2fZ+xE1nq92I2ex9OGx84kbzAqj/fsq4nyyhbN8aTFF3an4QVaIYwpNX4kCnj
dLZI6CWMEc6njekb1zpPty3AXFhhi+4aXUQreHDFjeqDFPmHd4mvh1pLiABPVJTXdDUKvbpyAw7r
Ef7oP9F2QqNNdTe3TIOvWpGOSNxXcBuug6zOtJpFo6eeUybD8OIzigUxl3Ej89sLDA1+qBx+L6by
vihz4PIoFxAdqC666wVnjUGqyjsQE8vV9N+mzv+tE/vBUCVZgB0Cm7mS8o9g+uX8Gv3Tvd2oNhW7
lQxsYtd/FZHPYDM3fri+ergiB1VrAFWXv92wx+sW+QKIJ4RdiThZKYtHlBc+OJeu/7yNBGWpdlhZ
ECUPjXspDpNtcsARzB3Bx6PfJkwPTNufxUy6tZ2zBNHIcgt0m5cJcVvbq1bh3e+ygs7j1isC3exZ
G/F0XE0HMRFZNWDZgSXr163lrIjtNFdaR+SVsbE2cm42CCaLcFHP5A6dY22gr6NW8vjcbdI7o4TB
u0BGPfghhy7cp7tFx93rdvacdoeN6XgK3ggHeLlARYviJG1ij8OOectRihD2oXNtQhlVY3AnvbIL
1lh7xWX201H6TZWfhIyj6yW42e2UCTdHiFPWh5xI29h37WR7TSYLuYUdWZWrxdfpTiLs6qKHt6Pm
5TCPTeyyegRBbzyd6XReQCfN/S4ao5okFT57+NSjDdvQNoAZuFjG8db/MEsiWjZXz7rJx+QF9Qch
EqqSVpBBNM0OuMx2PafndFE20r210PzhHnKewtHQEXnUU6RZM2yEGXRXYeqvSSI0xyiQEQXO/peK
uPJ3Wiwxml6li+yn0MAC6u7L3xGmejIekz7NfNUubs49TLdn2+81uZf+6HLj/lGcfjVhfndU1L8z
cZSCdmaCAID3nw/WP3UACqS6ss5t8fmka4bBrVX2xwOzQCvcJb6q0wyaZRuKkxsr8kTHy7U2DLfj
S9Y+aeDaoxcNac/KHpR541KFCwMyi374/RpeJny+21FE9GVciJX3y4JY463CIghE4bQ5rGvDf73q
ElX8U00uw7Ms3ha6IelfNRBlMvYCEW0Eiysu5h3SgkBWEzM94MyWEdJ3YUE/Ceq/umCuYJF+4mPx
UV42F0yuj7Cby5zDBZZFgxVitMKm7zE+zpG9RuYLKOe2QN3RwIAlPNVNMjiWdyxPKdJPfHe7Qeks
i34aNQyIcrYCE7JUX5m3hVFXeGrGW8hcuzA1f/M1bpYhvPPf80sZHV0gCjJ5KZ4Ta5yW8zS99rIe
3fMFd594lcpG5YBMv1+KNN1VlMPc//Z+tXWuB+yd3A0zBc6figNj3pdmPpZ25sw0RdWJ3LeaONLX
czX0OOLgWgHZtp63CZ966FuvcBrCWbT2yKUlOJ43lsJ7sWiR7JofgjY5y/Axn9PKTPTDVfYP1OhM
XlipNG8G0cHdpe102ye4KNwQxbSgcfsQKaiBtraAABPa+bbzcjGIBCi+w+1G4cyFnZBEO/DDtUUm
tVhGtkuPq00RftWo6+l8Pco2XIonLhqZvVmwzd6mz4bsaGqDyEM4bB22o5tUgOWtGh3g1ASXU5Fx
R6SuuB0Ygxqo8Qrk+iNJslOvRafyEpMcM5+VYcp2kLlIIjbOXWJq/r/btlEqLjxinHAyFVOGuNBy
p24KaWKFTRHzoF/ZeQkjamFdzRb7WI34hIBMU2ILWdnbeqatRU5ogWHclJld+OGgmsWn3zTS/pU1
Qkh+ZfxLP4FAvDBQ9j2LaicrNMx6iLVr3L9++a+FxBEOhFM1r9dWJtc8+ia5xN07a72WvvNTCbW7
YKUWPMHfjdTlpYA8V22Uslz6shEjFM1m1THTb3OnaMvBjnR+EnU43Pe0QhaGInL3ZzH2CuW/uY7y
qJvepBvayIT/5137+wx8ChPShKCcKOHBjCDNZMfhtHa6c4mYXd0oQ6W+2hxF/CtypsyOExLbhaGN
vUOjKIfbsuXct1NGl3cFnvM275aYvGqtTQatR02S3Ndb4/ZHReBDBOzlsL5nwG7l/W2+amUO70/i
QttNO5GSFsuWeOWl9XieQUi28MTPCom9n2ne75pwSXMSG31Zu9tntF2ov5myCGUCMKQZ33Odov22
iNw8+JHgtuW+lJzYjr1IxkZmlaxcrk8iCuqOvq9oA71YhmZgDJbBEMuyMUuwV4CZ34yxbsWu0dKr
Go609TAt1WqQBR9WLL6LLxSq+WUpERxxrOiyYE6IgjCiFAIUhUXUoZ3NqnkHkwOJnOkNqR9K2aHd
y/g+e3y8yGATJ9hu5eiVY1kPVWOqWYsYOp/wjRtAhzt9msfSVg7QWvJ3/+BS8cwrkaAvqbnhUEiM
bqVDKInotqRd3zLtDL0E4cX5npmlv6MXkdT+8NaZ8scgHhv10mz4FN4eFxOD/EAEf1EFIdMe7OSs
cgThnijK06DW72aZ8mfNHduYT4C6ATs3cCn62TR8x2XoJ0nSpj//l4RnnnLzJYOxql60MG++Lqvf
oC9MNFBCFrRsNY2CFKmBGlVqeSCUg+PPeMifuh4EVwaG7D9ut5I5QZO5s9HNfHywQ0bJPAz/qCig
JoKrVf6ibjOVsewUxNR+WMNHoqGhL2KsFeRId9ZAszRFRXH1Q+YkuaJ0huNuid3TeZ+mun8RImAl
dMLkJf4Xqv26b1q93d6QfsFslZOxH4a5SSodjPOL4Bda+PXSJFlrEhmn0w/HQK8ZnogiS2RFM8XS
Vb97Sqx8OcS4MTfZGW6eVMtW/kY8C1j98gvHlDq1ic3njq9VzsdQSaZNIVAzIjgF02r2dfSD6cho
FCtElZyfWl8H10CO+I0Qqh+Olgc1KmlFD/liYjjuT+w1U6CXmep51cbtpkBwKZwXo9YUJrTjGv++
4/xNbDO+1rFaJ3P46VZ2vHY55WEPwEIv7zZ1Neh+NKgzWgX5NAcXCZXYhfqAASZRsUmzovWfAXqD
we3FwjIp8QCLWHswWJgU4XtbBqSnSdxhyiG+Vs5w2VRzOtgPcpiMUbeStqRGKQCXQeaK7fEhWMvJ
OSMNmrzal+DFcwtZHEwdXyOzt1qkllhWNi+gS+8BmN1VFr73SzOIe5HFEzf56WhtA9OBmEiwt8za
Chvi2XTA9a6WemoUMMrF4jA9vDykSKs9LaQ70WZIGz621I2nWfmuhAnT+fbc5uOpuW/SIrmoGczL
7JFOFEzUIAw5LEOTUHg3q5OqhCD3BMkkZD75N3ACQa9PQ8itLVQQntmrd7H+PtcjYMB1MrBhu88j
xMG1my4rFJW+Tp40cDqsGlCD0W0LgTW42m4aA8uu4Pr0IHc6fgBOzEJMCmuzarGj8Teo63A3asem
zW+DMAB1cq69vlZiljsNppD8fYvIVVooxSBcaDiVuyneZv4ZjZsyP0D1z0Ze5OKXdGbrxUv5olW6
Bydc2RrGFnNxNxIwncJEd9rj1raLAccKEGEllQItG/Ccufll/0bSSQwYQ4tql8bA+3zmTV1tz2nX
J3DAbFz//TI8vV8splbae4ckFOMUt7hGvlb7LtyGHBMl/KIizcQ5Bq9h1TpUpLfotPvMxP+WIS2o
Llp6XzmiEMTZTur/6dII1M3S4W2SYZvim7t9oNE8IOjwf34OWDBRy5eWf+1xOP4wSpDula5/aptX
nhKZ7+8VlJxsczX4PMvXNWrWgwqxBQRd3md8pARSTTxknOC0uNT66p3W4diAZpVr5FrR5bLnOIlp
GEnY6HXB0p+buoMToP2Y79HBxJsIJHLNr2oibCdR3a87sXd+L7dhjEB654u2JzXAdwtcdtaOnpc/
D/bAo1JNh0dSbXqNMKcCkJ3bUxT9+yT4/MMNPol2TEVaAn5PPeA3KhT723iRND9JiX4LS5waprDd
PJSpjFoE3jtbwouwxtM32AclhMY41CR32FJnT4HgxaalW2Zp38X/NFhd65pyugzj5absMpmWlf0B
ioap/yZVtlO+TieK8IoeSXkAfqtG4jRI2uyQQOP8Ako8iDvQDXk0AwLBx3V7npWH1d+QVU17VANM
vd4n7uaTGL5dVG+BAVGTGQ7OCG/vGJQGM/bsSuU0oe3ilIVkITqpxyl6fD4jFGFkGO6qD+an6z96
PaEn+jMEvMD4JbsUvGnlE0fYPhGamCy9t+xPlMI03QDFc0V91Q5L5LJgNpTDJYbIUUR7ey1SzSnl
pbaaUvBuwO8ZXuAeFvXZjKa3FDDxbNDoXtSSxIju3CCehAE3orkql+pl/D7YB/nw5OFrSX3qCGWd
JFSsrapL7mfLIXZlFEyctgc2PjhgHy0NQa0iLB9tfX7/SFwGgbSZ7B8Pvs34KJd4YuHp/IL0S+89
aIhTwtAr305CnKHpibfO9BOGH2nfdvcQ0sn3bpeQQhclRSV1tysD/O0lUjZp4jha3dqzq41f7gai
RM2Z1pbU9GSMAzwFAzuOmqYm53Z7WsR7efs/MAep5FfXpjaNjSR9H0IB3/xzc0mIKFQ6cfbq3VGQ
utMEQD5AT5TijnkRdeLBUoGLd9lfzYgGqnr4A/qCwKfIgM2GY09aJa5AbL3R4fqIibZzc+uO8JfM
FH+1K5YNvVwbiVA7d42qLIj6iyJPyusiN2dnyESbjcUWBRGga08ucCGPDLLoZxvF54r9grBdQdsV
YbX6VqcIqUFBNvitwD1Rka6aF0D58bJoF110Hn8MUYXeq1vWLtMrmSIo0B5SK2mQlwTrlmydc0yg
J6L+JOwx6Pek0quQrSzTB28XljeVSvsEd8mU3yUSJUGUz36FTbvZozRWSxOw5QCkL2swzqr+az/h
buS4E3iWQosZ25WFlooKtgTgxyz4O+/qO76jAZgwtliQt5Q4C0CuYW4kHRFvhmHq8End8uClWQqC
ejLYbBagkIFbGqzvOwsOGCmeu11JtFltj8If9p7aymba36fWGMtNTr/4bmp4DyPpnjlCuLb5q4A9
K3IXlKl53eOU1be8xMaO4r9cy2lTHj6WyFya6BlW74dFOQ5uE0YkpihIi7pMY5RfdOVg7Jh/sGc5
+xPZDGvf0KtU1mqD+MDVpM9FMK+LJo3FRGxf2S7kbH67cuWl+1Mj2MvvsyboBWwO67iGo0sIv5xS
+2oBqTd7SMvICL4asmpksF3rsgK6mxLyiFJ5gtREeVRpm3CEYMFCb8XGQvXTpxIeprwuqzj52Sw+
PiPGvduPm7s9nMP347hCM68rACSy0dJysM0qLwIKIiSGxjtxXVe7k5TE2HG9cYN179Wac1BVlX2L
a2wXdAC26kTDOMojVGYIQBecQIV066/gzp6UGhV6IVh473/yh4ulBeJci4FXWTKOHHINvX91prKL
j0q4QQTnK3UlUrz+Qa/wdTc9eK5bWnARTTZHKCn03RIujl7D95ruOV4cXEdHprycFn999ldjbpQ7
9N9sRnmT2V2+DHm4sIHYvAos6x07xR1Jzo97bueqFoF4YFUyXyaS6EPTFE2Xy1wN3uCd+1S/Mdl7
RnF69Dr3aeanXyZtyGBJAEXBuzrMm88InL9c+8eFXdBrt9IpmLERTKN8e/MNGFpvNFKEK0lG5opg
an12eaESh3jPCDf6ALvbvbo3Et+78EPFtpr2NXfPCaePhrIjG9+BGw7DtHaQKf1FCRNqsg21XfD2
1TOHTXDPmWi0DXlFl9wvK5JU8bj7k2V/7cxSeMRY+ppA5FMC4Y5SGaSL7xnYKgcdodneSXOA+Z64
rMBcN71dUZ8svApRDTOY0m5WAOWlMBCunNMRqBkLXY9HQokPmWs4uFvDKSNDarzYL8DMm4xDQYAq
kJejOzl+W67US+wYq+GKFDnUVKcjHNOE09qg5Js3FaxzC8QuMXc6y7W1miIwiSNirvLy7ToXv9nA
C0nC92NZ0xjqd9xx1eE3a4Nbxre+CN4+Ay5HEqOaoN0iNw0OphYQhkmE/u1v2txBWx/WMCPd/hUZ
T3/7BqlTkqhaD/guiOT7NgBZ6ry1pS+JHmxf8gGqhPbeBl/XWSA+6UXDqQeaUSCt/V3KMDwDg8lr
IumMBYPw5lXMsNXMU0sM2nU5Nc0KTdmAZP0tau/c+lLrP43Lj5TskIGBce9li+ciVR9S3Or72Ljw
XDbJaUayCGhPJHT1LMILw6dBwAeT7Wzr80ea/fkqbAdCa99fK1pLXwQiZmqA2ae6dqv3vvP75tYZ
PYIgz3PqDFvoDenUCD+Mqfak3Az0YS8YEHPxbPNfLltwEn9iV99YcGX8RuJKg4DwK1clrOes6E/2
A6uhr/Z9Tp+iZBtc68E2TVW7FKKtNxZnNwyBc7G43d/y+MmCl9861qgdBhqj5G1clqaWiXFuLMyO
24cXYAEKvqdmb5/BZVmQl9vCeTd+fvdrS5LSDz3WlrDK30l39/zQvHdzyJ8aQ1sdPEW55VUG4Xse
odxBUYBh4DHhFIQ9nzvqfMHgxbCMyyknz9c933VwR+FufuoKWUJ5UBbrUcQiHdLNbDdDyA9jEHEB
6SEd546I1o0+e0iw9uwj8eDxo73kHHRu1DrYLS5Y0uCojZ2oTz7NIREgVV7ogDHXtSImYbGUpysV
ngYBHKgLNSqxBX+Kmi8789PLe4/GNboMm98UOwNmGiGog8XYy8XIsan4QUGwKWCdJasSG5602oTq
NhC31LeggJ9zUS/Aluf9leSsI6dF/sMoLPJ6LNI5uh5A8YyO4Lq/YHo+O+AT7jAQyJp0b3l/OxVe
iSKUz41Ytlfsk4g4SgX8DBtfRU359u/vWUs/Firm4ft3AITxgyLCC/vjxvGteRcLiB52Mozn9M/d
4BT/1RNCQk0GnXXVpJIR2mAM1H4AulUFep0Q1A3mvdnPK2yfq/ixMyUKtoXHM58sk8jp4gevxUPY
+DUQZ5ZlukFrst9km8KPxUj8wq5rwlpdTzO8XQ+Q6IB7hDEP2b82xLLruDEf5w9tbCLoIE6D4c9S
7iqAf+E6+S24CVTALOL1oWbTTZirjThioL1clmzqfp2bQa2D0RngUM59imXUJH6i3bGKV4jac4Fk
FKnOyj46uNaAQXmKRX+Tr0R6k5mGh8nHQK8HkyFrXrE12SnXyTj7BCfQioaxifNQGhmrxE4AXnwY
1VSIFejMM4DtJywtduyheyL1m7LMN5wsSGmvDWZolrIaKaZ/Chmu3AySui6hRbumJUJb8Fuil87w
ecRGC+S1cYRhxEQmZfANiNtjFQ8q3whb5P9xIOl0CgmDXJLHbJq6HIWXNDm2vMdhXRpk4tIziZ3r
lONRcBr3krHDcOU0QOFu/rifM3ky0tle2bXV2NIciGmYLRigMxcxbu6/cLR9nU2YUkpbY12+XhrF
H/7NZ8O0AbHQn6esuSD4wlk5bpnw9/xkbVg54E6+LgS2nHJblK1aeNJWTmnBrTXrUkSwivTrcRLt
+zc7Ir4bP6lVrSnlOwEssLFA1E4PNcKfm0UwJXIdGND2qaVc6rE81XQxqkdewllbLkTdMd5BIZW1
X87Bo8/3/LXl31hY+ee0CqrfvkEH9I7uctmEySzhuJ0182rq5zUlu9ROjDVNx/1SVoBMPgTwir31
CYFeCDP5RX+DOp4yHxSxxuIVHZ7eUXLBy+FneExVMDrp8yjJMejz0YYCqh6XYbp51iL/F88TX2IV
OZ4T34Pv3pvFgWNAX/miKW/teU4FnshMaobxS2PaDmlZWku9IaIyZQC/uNoD12v05v8Qnhcxgb4K
Yht00496CZciusdMG138O0zlV7C/O2tF1mauUjSunhuGli9XRAe/QJpGnwS/ZrQ/ii1J+ku7TdAa
1pAKxBqOiFm0zCvuQju4IORNB1tyzOdYohfaY/xuTFsHCjEQUUR3CSk30h8KCvpsYXqlEUNWlIod
3rsQ2Xc+WY02vFkuNsP/0KyxM/J3Kf2v6RDAsG3XOTIhTQ0n9x6r1qKU8TYHk42X5Bt+MfB90IbE
sgjOQBvU6SiVpdOiwD8Hr0F7Xt9vzQkp/2XXWEgd48b1QtyeW7f5ufq9xqJuarnlTl5449FiyriD
04h34WjlF2yJ4EA9dtDCbpRXdeLugpl+xUebQ0ELAUdP8PYtztT+COAMl9GTMHYYVFAs2K53mWet
zoNVLtQa90Kx+Kbp0GRIRC8uIU+j2CzyA/yko1MSq9m1t82pb0m7cbsFrOtLbrMAOqnb8mwnnurX
NaMGpqx3zTXmNClvqxjn7B6ea4YDy5Bquzwgrp3CplGK9ojXGJoWTlD+ycfhEz8P30tx0V1njMLF
OC3PT5YEBA80pDOkPpx1V+2WO5xgesT4DcNMzcgCUqREGljbAS/Ic0SX5YXXq2nFachD3GE+/KbT
WpI1GehOisZs6FCl+16YrjwIyEFSqg+Wdo6GQzSXgmsJBNvWexof/CtmO+/yT21VHagWpYUYlv3I
hLPgs1tkJioP27Oh313CWFaSq6HQzveIJl4yGFzyZTiWwA9DUamIuLA2DPwOm09Oep6vv7nExzF6
vnS8dw8TTU6eSpN88z6y+hca6d50fV7cZVdrAxzpaXj7bWPy67aGc+9OFZsEjPMmEAnL6pGrlz/C
H4g3uaorAHD60N4DmUiyzR6ermypR43fi7BJgikfEADeq6Q6eTqH0H95+XPZBU8keDJ8+IxvXhff
7+cyjmEWSnLSFXCkj2WjxGPTYxTUFUFnn/oqA/D6KnNgs+u/9ClxsAWaDyOmNKL/maMEOTcx85ik
FidaKWjazejpAs+hGI8pD4Bat7s1oOFBOBUTjKaIjW0a2neGI5xXAn463513wdTByGIDO/Axehko
vTh0+iEkUFq38KOhZ+vKq1nmcpJnkW3PmqduJCR1wsli58YQcnx2RPPYi+7qqGm3NTvTtGmLyKOi
Ht+gjCax2XpV6xuGaS56XHXUbGQNH97Fj7broq8flIAosPWVTS5PMQ9Rr1Uv8874TB+klyJF+q94
0XJgHOJqiKgALYeQcotQbzw/J1gP1pT6lSN+3QBZqTpQ75zAk0nXkVN46gzc72tZlr8jkmxGpYWg
xKdTt8yXR2egyHUEW2ZAfiL2q5XL3R0eAAKSkkgrzILJsu4kkyBnek+GKBErYsgqiLhXlElnbmjf
gF0uo/DMVqA8tUY0zMW1RRxz7ebPRVcC7VlbOBRaBJCNEVLRWIEw+deXN0yVexP3QoXG/89X6waX
/9hy9OP5UZwURJ9yRaRrFK8ruxYg91Aso0C+cDB88oiEJfvCHwLY/OglXaeqk7xkOJgH6BCsxTl7
7sUOcKAQ83GIc0ViR3FpK5O5SDBQED62+SdgdfJNqa+YRqcKpzN0yDy/HhsTVU7kwXkt9QNsnovq
eagZ9NotUUiL7kl18EA/l95M4/3qWDMQrvse0dOztqwqzcD3L4vj+bKhkYfQZHbKVRaS7w1bdTon
mhDilw14QtCZBTRTjYA9AvtH2g0HKMKrzGH1tBbLkwVSkXJP7XaIQ3v87OKtyyVIY780TTHAuetU
fRA7bFjDduXBzDL9yf6xj74WQ7JsI23ePXPxiZPUfQvOkM/7Odsuc7r+4ULpTYI57BpezfRKrV9n
bsfnZv1W0r5i6TCSoBKDyqvNC8o7PQsssfmemaor57QkNF89r9AlnS95f17XNVrGRJBnl/Z7w9mW
AJGbCRR1ZhMRhMlaFo4D8vlpwNwEBCiNlesVLedYOtn9FekHytCLkHpwb7UY5SbQ4p3fGqsQwDnj
svFYD5mYYONWW6pipu7OTP738vrJKpiN0CrnX1jlcV31cv1nrdMnfntMMiNEos9aE7xNGDythFjk
mKzCf0oQ3yJr4+hO+Ibi7ZrudQTTpohXS1pTdHI26fIWgN2XTyNtd6pMcWa6rCLhwUUcesmDq9sy
zxVR2WY5aYQwrYauMcpz2isFcaEgBewhEsVuC+4GkMRxYcTm7XZ1v9GqffJY2Md/WsBhHbjs333s
s7kdoY8MBSCeOMQXz/Fv7vZd0SL/3MlIZ78Q60oIQv+BUL8GAsFafTGaaxvPuOkhgqffIgttir4s
iB7Y8wGOLt7Z6YiGW3ecaGHZqUqOt791O1xPnfHLgp1HoewEMX/ZBKW0elPrHKJEFtFj6PqpfyrP
uWx765w8pKYqzCwsW7D82DVaxO6mWSEaVoeKR5lBbLN0d7zkLPE6xwQpn/Oi/LlYjnwgJK/HL67p
MwWaCtlqD8uerF5kF+1YKcULnrSbxqMmkRw9BCKHcbb9xbsMNYmzGeNVYKtwaScFcf3cxCibT5PX
ZSkS0OZnvvhM2cfaODgJRnVhBQhGBaPwv40nGXV3RZ3UFshbC5cEKQCIusBPuz8FAZ9o3r3pWZB2
4bXF/RvP8nxIyvH9FZt/Wd6MHlpoc9P5I+vVZp/3zmi1eD+/8OwUFtSaHPelm7nzHjH0qPT6cvkm
ETyBaxPA8gcy1yiZnP46FBrFIyTBb40LV4CG8fodyECKKS3ibuI2vwxIxPmg1ukZCJRC0tkDBC+H
HYg6WP9oU2zNR5I+f+tEu7NEApGYbj7BuQpierGEo4eUk96kHMi3tyPTohtbjgQEE1yqQ4sosfwY
2wZTbYkXXd7hQ+3BIG+xKC6uuK2uT+ib65lMvn9Vus10oQwsVQI72pKwuGy4IWvbauwWVQJ3S1Z1
itsyw1WarykbNtx19u+sILpZ1C8ymplbZk3syRbfqmqm3FzuEoNOgnQchqG6m8GzKPcvc3oEwZ+b
K0Aq4aoR4V3hLqRDJWZQeS+Vcpt7+hnRX1NEmNK2PetaBk51/bjiXJxasaKew0hsRzobkeA6PrtI
Dm8VpS1YfBjICLpz6nHOx+W03xmInjcSX4Sx03+mYnxMtaVkxtFZxQtrlY28v+au8LvCCh22flnS
CAZAy0Cju5m9knkYGUOx1XpLqt3J/57zEEQM0cRgVSFd9dnjMgHJ5nyHMgMhX9Gt8u3LogwpO7O7
9rHZGLmoOlrQnKguSc9cinoaMO30/E4z+Sm3ycKdpvi6GLZatetrM7ZR1tPgNzkxaSxd4cblbVW2
Zu+tf7VH9MIlkEOLSqtFGVCoBUUM5hGDqwP4a+jZrxkFlqU+HxS6aIm2DISaPQGGfGqLfmpKuQQq
bmsiOR9DzGDsVpSW5nRJQ4LrfJg5fbUZ3LN77PkfJ/qbtThXklN2ROaYUJ66Eg1n2nCKdBJiW/v8
7wFpWgs8Gl/WIMNiP5zLbh+5aD3A2RAFipsrm34IhkK2rr3eQek369ajllDCAnCTts/9FrHpGFQd
OGq6l9Ei4kG42B6hcX3P022c8Vg5EVdtVEYsTjrf5DWggpYw7+bP3HWNVr+9xu/A6ua1Mdus1Acg
j0irxFdmGGxvsyJlW1wFj6ULfdzBRjcETTv3TBPCC6pgjJ/ijQSiAhUPYta7JsUAPqM2+1/Q155F
EUi1Pz/DqhN5D7Lp0oBagIjzJA4i6HSd2mnq84pYHQvs64equ50KRRUKmEc2MSkdVQemnyL4JKCM
0YxbrVDkrvRDgBs5nqrLqrnyGtpB0NuErFYGymlJlnGRYzfpJXWH8icbP/6P65Wtn5MZdsN8a3Xi
c1q8ryu0qmsB+O+g9hi96DPG7nFRDJVoYP/H6jOhjU6dUH0gWO+hlOKvMX1vdoqVLv6j46UEoSYN
rTybZniOgmyjO5E1sTHHxY7j3p1+7EtyWEwegHY0b1L0cS3XmHJ47G/eGgRK216w/gynBiLNa8ya
ZzH/fkqcs0EgHC1SGR2BXRzs2fCitzYabk5EjCaRSkmaUv8CsktPaMBDT6yOt6zquWSHCZmD5hx6
coWXD6eg9lDerMcW5q+fy2IhwakDXlQwB7rH19NGuzQw+wbbHbXEKG1kKJbO56kiR4ivQtuP0kPv
X5x3RSMpIHZfTdVt1mS4VrDsUYhl4al1gyJEfVtfvNphxCDgVA7slRwI+HIu5p5kuUAjeNbF9ipx
pge7KtrX4ieesHn1aJvB/kWCt2AvwN2r//eXCp10bOJcYjnCAXRE5DxjcLWEd+7Ue3GPOyZsZNu0
CV8yjnVm+m3Lw6Q2Uk9ozg6vTpmPoABtgbgP7PgAAQhk2G+km8wJlQyfgOqqAWm06BjdykcJoiIN
4phMUAyyq6zqsF5de11az+MLEwDW/bnN6ubcQI06/poKcTQDRWE9PdqtzQ45UxXcaJTeBeitQG7f
LTHFByM6yiblX/DC2EjABKpFeeCxDjcwLVg+UQjZhoagVMDNsreSir36Soesw7VerKRnOG+3OMh6
XS71ytLAw9Rt9s4hulJ7pkH3SQvwAZzmQ1bQnN/DyQR/DkHYqvG/orMOiv+1FynmNFoMnrwuS3iG
/tfdAtkO092OZbMP94wCXvCgG30xv/Ac4gR8X3a5UlnK+2qGhteKIuqDe6BD2oW131vDOeoe8r6S
zln6d+Vbiypd43HEgI61onbtrK9YQKWu2Kbbbq5OrsSsMoTz3HsGo2fqufTdChS17pkfY0YJnPwT
ob40nln69bRpzus/ksAw80iANBJk+Ub89IrU7nZ5RJgDwUYpp/uG79G+oyIyJLNZismDxsd3U3pQ
KGlfOHvYZE2awkR9+SL9o4SX+lg9cQhTHXcSYMzuiCqFOBEtqE+bv75gHGnIinkknGKrxmPHfLiV
mejxRcsvsCehLfczVp7PGnONVfxaKEw+m1yDcTytYpv0v6iSqDRItxjfQvAavFEmoDA+Y/Xu7RUQ
LwOO0XVakXDiaK8jFK+QYyQKyECP9dwRZVGXZTRiSlODkNMUDMm/aqpA2kW1U5s/TpSWAwdrgE1X
EeGAbyk2HVeKYYF++X/F3Az5HbbQCTboKSslujOq0OKcpA4SlfE4JetoZ+OrEjP8AahNXrFy4qIe
/58MX2UDOmeAX1shFee+uH/RKkK+2Yln4LEJVBZnJLdEUOy90k/QoRPOILV/3TZf+zw4AEXDM5tW
J62Xf4HN9mj4+mcPVU/6xIrEMfzndzYeEstitux6u+nThMVqojXBj9WCfiwvAZgHbDh5Ug5oluaD
Vu/mxfmd3lLb5JO1YNBo1dxLWdqTwQepTU8=
`pragma protect end_protected
