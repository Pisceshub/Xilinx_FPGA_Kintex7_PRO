`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10176)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEFAeIFdJsw8nqrbeqLVZGFxhSk4F0cwY5Ne1F272o0cQmxeiMIrKUrsq
kNtg5ftPPpo2wVV0RLB8+ELuu+ISPu8EzSxxRDIgD2CfspEhJ7aUgvwTWyWT3WJTEsyCErD/A8oj
u5DVj+0lzp4tKCXbOpxUCew52xjZcM9QwrRKd/qkXvTeQsOWZHcVtiXjE6PKIXDmCwD+kZ05jXBh
VYbae6ymkAsWx5cesbWIAYB6QayGjw6efiO6VbVDTfS6hFpev5FUmum0pFcqi9NlHMcyUQO73vKu
o04hhKAE/k42lLtkh0sykePoQPnnNBMVRVQDkwDWpbk36CKRJt/GB3HrZuas82nspyLyqIra4TC+
q240T+39vf51VNVi7AAIGBtTfQ976NgOFrU5xhKnBznuj9l1YlW3eYZr+Z90DEG7HzvB3Iqe60Qa
f3gkSGuAiHbcsZ9XGOipZAC44BbLNLHegPJofx4j4GS3QdK/8PQCMHpjs4lW3elNRY+sZterLSmT
PF8lHEp3x10qORpuVYxYMjTErfJ9pLLOJt3zFDMAq/on4lNKkrSX9RxBRyuJ0QRIqUCacqNEiB7E
sklhKyd8Rnw31kdoOErroUx2lZCPBQOR34Iy1I08+KnfKtUKe32XC23fNclWKmTMJ025tYRBnRwx
w/et9ejo+HS+iMUZmeCSkuKA5+8bOJRaitWDZ/ghtjwF8jvKfLcxVOY/i709n/XkqnttS8djY7QN
fTjffhUDKoFGB7O25JijWvHr7es+cp6uJEVmPQQqpu7yVWn4IDaksPk7mcC1AZMF5YfqMRWqOjpg
B+YO4JRmyD01HkZVCkY1HS8xqLXE9zXg47vWeYkEHZHLYc/wwks88b2U429FQbWcujMaxpzQNymD
5EYsKRWcd5xRtj1/MyDouHkFJV8HInGvqnzl1OuEHmgg+R5MzGQPV0FpAc6ZwhIizHhN88tEW5B/
mijVo+cV7z7utp1aBxVf3pVlvNfhKvewtFCuhFvv7kEglAHck3K9fneyNF7YkoVUPZ9Ofk1pZtjF
NmCKcU7hSfI+GNByoV/Id5AMOGEOIpo9LUFgfeDZtkVRl1w/+ILPNeP1VaHxHGYWZWR6mmTJwYXd
RfGMdnYpZ1CR0CAMdVWqwuUr2jYPeoaNGExrgQGQsbBZL/YJRS9Rg8kKHTW4Ux0e59+JV2zTy6YC
XK6BJ8DtVUhXzSg8KeWz7CV9urWgDagOLIBbfBKo91SlGnhvPWDguI0nrrBZP5MVk8yM1k989lFN
7bYQy9MS5seuVR4ZgddyYhLrF8NVinOtxYmyjP7QBeeZyOa7r1FQI76HMkW99wJk5A2tAznKuLJb
YZRTSziR79ZJ4odtMgOpmaYsoG7GOkkK5zzNA6SyPZshkxrEbuz+10yYmjwQhH+QyHC/gR62XYYh
juPRxqDIwxg4K1kqCqI2SQj8YFDUh5V6Q00WxTcco7GFQQdW0IJnKlj5nD5wIgozEvhX9k7uO75r
tkaT31N+ftnefbCIegNyBhkEIkCeDX/p6t7TRICmeBNjEemMkbzsG1UpioFM0WvPxs5zj6C1yJF9
oA9trSvrps0yO7+8TkC+LPeSDmXAPCzSNeI5wa01Rriv89lV0R7Nb6Se1Gai8z1jidvenW6OZtwj
zg1Y8adJSpm7WckCerSBpcraYvu/aT/2548MaT1fF32w2oalf8WWkji/BGbfCbuE8zEEY56pnfA0
jWvn5fqkq0YIAwP9iJxVsBJE2sUmhDPHSHoBB8g3ORAba7MhbN+EoDzp9o3R47Jm4kKt3OaAhuJX
k5m4pfRhzoRBxxBtryMsYreR+yF1SdJRbbtTRCWhC3oIZYTmrXrFke6d77EkdAl6lUPVSDmXhVYZ
TlGwqdsdeKHhySqz5Olr16HyNQ57y04q/ie8A/VIgzQBh7O3xw6E40/URxOEYAhQYf8j0V9R7LGL
jOgK25OZ26hYMEgD6A5IMVmn161dmDSJITo5pZMhBWua0R4ng4Z/m+ZLWmj5VCNdodB2RMa9A3aL
5QJrTZMg8qAeNWiy75LDoRvg+hGz0CFc+a2d/tUObNjTdqjXmFUv7AUoKQegJTvLG1bYy+CeKl7h
p7D+u3Yfk3+mNIgtmDLon7aSSqXn/5k2CvOuz4UTLaiykbuWvwhEAloCKHzD0/+Uc/3P1vpGYVXh
G+MWQCIrgeSiN5B9+spZMlVfUj8S1KhBRbjNppmr0QncUxNXnWWy6UydObS6t61+vUrdHOXFmBDM
kbdKIsInBmlk5EfHTnAGdST59yFd/wCSzPcAyxArMC65ysctYj5ctbj//M7cH5/MknXkiUAeOOcq
O3Oaxs7PszLcVMwL02swjfSzVAeW+yZqe5HUnUk1+6AQiJ4R/ak38ODJolha1V6oJEpvhnC/qSF5
e7gulQOIillmffRavBvWRrcZtkLObvBTz+MWxSKOiHF8grfeZ0+6ab63Ll5BkP2Zvi3rd4yAYSD2
VPh7QpNmEF6ANhSnNugKpn+8FAds4WuyVi+xi5p0I5QC5kTYDtKKlZ4rK7wacTglqSJOQDdIVuO2
cdNfZwcDJHqj2YLNnxzTXLfbJ00sawzkpYxzlnmqpfSqH8ll7zyr8Ej8fWvYC82cYf0SZHeBCpx/
m/Rzyg0b7g16HPr7bqHMJnJO50FM44K9YoFvtFk+bWlFyxO/vQapLEB4OLc/OHqLxISXZP0nJKwB
uEngw5h8SCyNVX2BZxTnVGcL1Ej0/5MZm3uzQ/orEQS451bAMYonzkNkPOtsOeW6eJ9jmkb/m7Ox
HhokG+8JYHoYqAo8BPsGoMrO+LF0dOJz5SM4zGZZpoY4TKqUG2OfTlbUOmFaXRHuPl9Yj6/OJPxt
TJw9OBEDXCrimHZi3rM7rCjmz0bDOwcaGuh+yXExnYyOTrOuAPRr764LXxXZQFUFxGUUvbz2XZS8
y9K3jfjj9nmju3DVp0ukMH9edicRGAtWo3CZzpQ7FDfPAwvus3CQjb1PwhPxmhzCMgcURgJ5FSDJ
duYENZFU+K8IGAbBjXBM9a8ECuvTwaFrVpRtyHazHDGVmRAgmDEg5IDGeb38n8SXK8CkmhTOAuXS
rGj+bdpfsEN3g/cZ5iCeJR1DxNWaMsmmD0AoJx/MWZ2wdNRizTcgbKFRcXzk1Lv3U4FDlP0jcpGJ
Zhq2CZNMnJQfeJGr156PtXPIbtnVvxV2FWSsIqaHXijKtBHv9kOlaI9z4Gf/3P/9fJZPT0wvO/xh
RfduPzYWnGV2+OWW6O+fnNKE7+2HTWGGY5rC0D+2KDRk+zg0jGCjRmHooEEWHiIFW18aHbcYeGBo
rPphD+c8lJLmayq1XK8bP+bjIu/GhBj80OZW2MVLp38MDPXl4s+CmOPr22DO5s8zqXAQXZYBBtsX
PBrN76rjFAwDQQzZB6loqy8GlrsP2cJ7g/57WQRk2dRtgtQqIuL0K3souKp2vR5UKpEluyRilovH
OuzWK5e9wTlo/Xpc/vuSKw3xifPzNxVEWDoD1ezXuu0YflXcxVGTuvaSJ1CuaYMXN4CIQKOAH1X9
VxoAKmPdwrRz1uVNhrwdNBg9rnQwZoCihy/oQtM98P6nka4AqgfU7+gcZdUCEygU3dLuiEMUlnnI
FhF4f0cnFgbF9FXaQeUK4W3wd2kZrMEQ5pP+6OpIZRCEsQVtUTSwtewImADclIdkFypms1BXZIaW
IfFUSNC+SbWK11/Sea2O3AFVIhMWD79Q4eFPR+S4cKIZxHUVAaNsNwK7qvrtOckoMrYzBIaJy8fe
Vta8qP9JFSDaClKNkP+wvBMzPGY499uERyJZtF9bhanr84RxCes5LMX724oYENnvBSgqqFTf3zgI
vp54lTaEhOkOCnbuv6IBwEisW79bsDhdvsAYs+aub0wermiGj7u69RANbvBaIIxzTOr/yg9IFNVx
Cnn7Xx3NARqLVFW2frQCNpP3F8I2ld2Erygz9mXCkXrSiWyey2w+wI0JyP/Yjj3XreYMQ0tohvvf
1w2fRPg0DGce5FzSQ8GLocPZkM9K96IsfKl/3+cCQh/IZ1Zg8UL6TKwRXDpIdZkoHM+KRL+WEMFQ
2welOc+4uCWMLuX2VwHDhyFfJritYr8Q7JiVx4rBR9Ana47aDWAay2qZMF9CclCIkXYHE6kwKhiy
btW4NGy55z+H9RpiE1qijY9WIr1KiaNUHmJMQNOPkXFu/nrNGrwhLbdpypQQbdj+nQmKM90jmcKq
DqZhsWIHw+9p6JEjfLpUbMOHdwA3zfw3ztGSCr87vBeNNjyVtI1snpfXXiNhsJ0F7Kv8LlOlF691
HTWvjKQwHWOfoZ39RDVvEpOLUB28nzwu8T58vHCLI5qu+N/E917JXJvFaxgbTghXmwH0omhtkueW
B7L57yFeQYyt7g2qQRPE4Dtt7A0yRFYGWAE51WAgltW2a6OeRayOYQALWkWQ/PYcORJ6Pg/TyeTj
5f6pQvfqKNqFMEDjiuVUFda8jVusT3aij0NIcOPKFcBNcyXwAGggxMsF3hkgxO+EdiIw77qm1NOh
3uZkrDwAZ2V23pP0fP7JUg6muPI6v6dYrMm4/SHdDkE9towLxUbhic3GZuO8L6Bz+srYvyvT/5G5
5RuCq0VIGoICzESy3R/4n5sPpQCe38C1c7P1PA2P8X2kcVPgx6UvVRWggMQRyZEKUxLEf9x5dM9m
FSJza6UbvMLFCwWJvSm/mJ9lIU5LcSseScVvu00xxT9zR9jWXvl866cfhHh034fPvgUCX/rr82zW
OtiDN+LVPnOJ7PQ+POSKDNNfgPF+sLzphZob5pxqeZySBZzmJZHuHipgsIoZbyxoZsVHA1F+dFpJ
3EVznVWvSm/Kh8h/NVl6zAMUT4b4DMYadM8HzloaeL+BXSpad9KBYdQT2jdpxKcDKi1q98gf2ZMW
dCJ8QgPBCvJmJLhsGgqUqS09CfT+/m6eRmdNHK82qZdtbTsUVHzHXLUnzX8sbuW5lXhDjHjww2tg
xBvS80NoDJt/EvNncK3sv8kX6lceCSO22BbvK0oCHZEpWXTxfn5aEJyI8KMHRGXHpyRQMT4G8DsQ
kWSFz4DW1oTgh935HuafvrXM5BglKO1ChwdNNoJhgafT+F5zWSKcNXsPq+3++x5d6wpGjS5jS95t
KonXDecBYB2guZ3GJMbL0xFxXhgm4zF/SdV+1Z73HA0ZR5fFtLk3Gvdxv8IFlD8rXbPRaqHpWzkZ
1QT0l0tWmK9dEk/xGFOtouC/pdP0Uk7+CkpnZsTZK8CG2dnjOwPhKUCh/3oQ6SvXSgH9+IK6TvvP
/gCNFEKIBcPqYSP07O7I108KgQBwTY+zWUdxDS1joe70wUaPzXtIV8gzS3OS9PJiY3YzyzmN/xhE
5XePRkSgjpqjdEMWBT9VEHrlcTzYN/NZuvEYGJN7Hsj7t1ZhA8FsaF9WEwKpIY5VBzZmf9yA7TqB
G6xwLEUecBMEp+4L6oO/H76L7mPyq1jTvhs00uJexXPvpgPfsyI0FhIR8gc6Tt+aa+C/BYamvHdk
sTc6KYDAjVj1Gi/vyin4QBsDPTWqtPmCrCHVKrZnNHRqUPgT4j59mCgCumfytmJ9OS+aiVY73i9+
4gw/j3Z/0zLqRIHPimProULuhKGeqZhXXo4QucdtSuGeHmBfktAyuEmGggqkLRA2czagztGD8S1p
YbccSKfci9msrhNdMD3qyTAR/ITZTtsfG7mWxOhgaso+7NZ51hB0zPkM1ZEwakgqRVU6M2/wi8qT
dvWjhHqdc0z3Y9U5AWCz4/GDIgCEoYhxgpxUnp/Xy83fwqf4zyAoOnD5H5hZuyRxdspIVtpqI6P4
LVTISD0kmZ0/MfexExrZOGVsf1ys+pniDPt++z45c4JikyDBVT3JbCQyYTidE+jZWN0oMk/b6Rco
75b8WAHSEo8LDQ9uRZV9FpwBeiF0hK3Xsy+21qjR/Tt1wQzZzz42Bs+XoxfQS2m8HVvIIM5DY3Ij
DybMBIdOX81tjjcYVi605zkqmSduQfxU+vuuQ+n2Gsfav+e0OUN6Xkva2SVOzxNRFckC7IUDKvK9
0Lrm6p8uqGxaOzrblgOIAXOAO0q2FdueMPKBKTuiLEYXCDhCik+wrETrF9OQvXBR1UULN/tC927R
djMpWjMh1x0zwrHSTMdDX59JZVafwwA+ffE0nCQ4TQ0wdlgqzsnjNvxAL0nzkMw9YcjJmb+cmEx1
Clyfsw8202gthVCzPcvRGrMZr/VPfOl9vw5qOQsAQawlgkXAul5LmebZVS9RTRDDRXtIXjzXPNAX
xRyq0dz/CF3QHFU23LPDldSy8kbDCCpVC6J8u8N8EoOeUH6h7h/8p8Gmz//ZvF7FsXC+AjX1n7nB
4PNnKmhhZRzDef1pNadYAWOwfAnkxQzWrDsruRnWoSZ5uOf+ZrmbrhUkz8nOILwLcA+Fcs+q2NfB
JrNLVUsvQMvoa9dIEaRJghZ9KfGrtb4mLCiTstdjNW0GYXwmpOfx2hPFBo0l/lVmPfwcHptKChZ6
n8pO2psTNalCnOLBS80zByDPsC+ICPzD9+Iqa0qiBpTmnJjgO2uE6ALVTcgyLwx9FvnFQX9MnV3J
FhX5HlMWK08mIAOgSTFbNqm9uU1JJXTOPYudsutnWELrNScUzhBeqJ9G/ZKBKdlQqEiSF5hKZjUx
aePAK+lMzVD5b6II1UljBKQfi4rEVSX6sUDeTM9dJbD25WXU24essVFiWdfqyyIWOKJzUi8seJ/j
ejuXV2YnM3HaTU8G3GzATP95rahmyiIgoWwC4OvPazdppvElthJtQzz+CNxKXW4OhI7EuzAj6v4C
U2TuJ6EdOkRPTYOXDgH9ZZea6g4oHyEut89l4j9J4PJcjGp6jWAg5Yy5kdrngJBAgo0dk6Up/6+s
n271J2tanon+Rl1yAtiVQIOG/zlDSbBrY+VHj/7Bkn0e8nf+PgWjZwqyYiNI83DbTwE6ekIzvPEq
SGATtl1ouNqUT5SyosCnQNcw05zQXLSfemFO4xY07yErhmAWkXoX1AMAoiYwMANRSbBWjW8BRV6l
P3aD0fUunRI9WtdjqvT4OwFzV2/PUrPfJ984f1dM71WDXcI+T+VyZPtz4q5tGlQbFlrg7dghG16v
BmjSZMaS/YVduiKcD0WdF274khK67ekRfIMRhGaosIMumChAdUqDPW17wkHwGhWXlEbpa4LJrO12
32qIyn25Zj0Rg+1Na4oqOFwwZHBNbe0nf6TG0eSCQ1aoI2K9IDS9k8qqGM5ojcNG0HZLWEdITiOr
QijY6X6quhDrBdjSHLVz3+1LLrTc0Gm/hGP0xcMTyionIhiiwLrYZQzBuake5k61p3BAnXKeawly
cqwhP5kgz4B+T7Ir9o1AqNw5wclXeMOaLJhHx0cEv0OtfdyognZtcDaikDwGqvslQXiDYe5np+7X
3l3IqKTyqVug8BmyMcg6gUxymXHM6mtFR9HvvGUMSLSAEj9NgqpSUukpT/ZvXkkasFvpnSZFXTFu
Enx8hmpZoJRleY4zd17xQMPsOy8SQQxAnQkrx2u/Bv+zh9pdTLvTMzSLRxa0J3BYFAkTa5Qrz/ip
3iLROveXmLBd7QH2RYTak91t6MF0FLJrUZRjSPCnqJ1WfNhnqMVPsfB1j5DSWr8cPJv5rVRiCSZG
KhNjvDnqJtM5/H7FoLV9Nn0Hen1EOBKQjcFYgyLTKOYm3JHB7Te+PolaSORAcp/k+KQHx7vJcquA
AdTh8aFXGfS/VqOBlCsQlEK1lvmDR/j+ggerrM9dsaNLSS9Q9FXsg6wSdY5J6H9g64et3NFd0x8U
if5ll287KjtaZd4CWWVKkw2FzIsqTXYPuVJJD6KgQrv9yMLHr9oWSW1bmMGBVCegcSnVQW1ldAye
CAeGAshD7HHsqm4XoGst3lLQSsRcRhEm9i4TRfqtiPcDAffQiigjtbC5t1m1uHOQtv4r3AbT/ec5
IfC7pRK+65QXK+oHV72q4ouboXpfBXxfsvu6vOCr/WblEnAsK+IdSUorg84O0Wz/tc3UJeqzqZ1Z
LBoCtFJT6FWweUR1h8l3V4e2OcnJEsddzHwv0aQG3OU5q//FLnX8LdryeYl1gdz1zyH01cPI0UNK
TkynTrpR+cHYV3dJfn43QPYmpp0Ymu+uevxJP/+U4qkkrtupVxpDcSsP3pdX4OqnBFDXPKVJ6BxF
V5NtVAXbqi8f6qXfAORHeitVFRLzHGfiJpqmSjc0Uhqzy1T3m88166O7sdAg7eVxyUdQMnqdj+Ir
p9jayqpdV/hKnGZEudAZ5orb31TQuuuFIu3YzuCgtPM8vkJjZY6pGPnG+GPMxt02YspHJGga/+cu
GwKPdy6ico/B6rFFxxZzgkaiL8x3gcLcLrYIM0SMXII/4uWuhWquwS1ZYUuA05jnOiUA51I6AoCV
9cGoPmvztfDWfrnrdnkZmJXD7TXgeJzF3RpjLrwAbELKdg7xHdqCbsLbrvNVq4Dz5MTFK/Pw4g/z
JloG3YPpeOC8NVNcI0G490UTDCwkMXwjoKTm17ss7e+g32ZouYSI0MAW2P920lV/G1+/iXKpig2j
tAO1Cjq00tP0z13AE6iDZCnhmc8AroYgxAH7GEGjQ3ctQAXFH/yW2h8lYy7RylUB69YjruJ6PX+L
idiI5OtayyTXTqbtnnG6nwxDZhM1FHMkVKsjTorDIZWKCpeZm6RPfPwfyeik8MPQVl9rrZASQ2rV
8ZS7hISISCxXgWVHiyFRloM/FGxf9CHYCsLyW4OqKRJLL68lBWpo9eu0NJ1Nf8w4WL56sVhL8y0P
7YQJBKDto6jAdD0BxG3/TNTuUJcexEnTGKw/aeGrB+JJa9BS89mhrvCWLOHBGDFtpbxM4Y6raLmB
AmO2uDfAUjM/P+uYz+qXWQyLRHQvKNZSfAIoKzXYWtNzg40zA2euTfjQdda0hMAWqYFstye/NRXJ
JKEKLu+wF/cCeunCkq0x0tJrZ9NSRad80mgqyOjU1gs5vFnVGRR3WnG82GojRAD2OjO6/07uE1Xj
WwKJCKMY+ZA3zn3hBgsbLui61qZDXwjzHs0UyvfuaFD0Q4Phf4n7o71QdzNRGtqhEzfFDI8oml70
ztbIjjbnN6n7ad+MZVWgwbCgT7SuFcAOHSg9lUaksWz0sFCylQW84tv6MtTzWgNS0ph9Pi8fw0Gj
aJRkoTU/VWA+xn7RZCIQXQhdFZGuk204yFcnXj//u9vG5f+eSs+teK039aEQkPI1XC490HGB0c8u
g/+tgENZlyK5OxqDrPtn2sUhUU2/m3OR6NOCv1z+Tn7xfzhzE2nEwl49nOtWzKmOW3vxG3WNny8J
Tai3Rx2gf9YAIVhuBSDOVQIhGX/uBmQsquuJbnNfie7SxVACOwTGUQCVTfTYAVwZfHF1K5OH5AL2
Vp7MH0bIuggzsJMEekkdj/D4OGko11+1VBTi4+MeNL+3KlEqLFvxcjuap2u2XJ2ihD9q87DrJdAB
fXp9Pf6FUFoDDgDsL4oQD1rzvxU81buxEdI1LrJdeMS3jr1jsxNyTTdXdBmQbtZmYsg0NqyeVrv2
Yj2hbWSk9IEaMtr9JUz9XEGLnAD1VBYaRH7qFpRNQvxO0ylmWy6UDrVHgqVs8zqycf1UtseD88ab
0FPWn5cGmuAmEWMb3+xMstS/6KGtiMJaPH5AOQ+V4PcUtK8Ji/WDfyikqulg97RkcQLnqwfEUDsh
0hLXG5WEq21ynHb+7gj0PtBTosMxp9R2c1jMXYeg1ZEL2sDsgauwtowwy15lBX7JlYLGXtmjZOUz
S3GWdfWyprSui9y4dE0HNOne7TTPRU6dzoXUsN0zH6lwPIA7JDwMqa64/A0rLGpgkNSRIMq+8Tpe
lwKDQ0+Z6a39eM/0f1p9A79/Rwq77CkFm9jLVZb+wKVkJZ7c9OcZyacbsia4EAulKm/Yt9cOOnSv
Y6r5o85v6CYKH7ZhOhcGPvk/XrsRXAD1p0qpagB+aD7dwFaT/C15D5RZn/QsiEzhlzDYJySJggdp
3uAvPcPlI+0PsztIdU9pW+8g2QAoXH0uMVuoN+svmuB8j506xH56Y2xlTbi+QALHJir6oz2rWx3x
Eco7eabTrU9vsxpEM67gPL6X+XcQ6EjSon+jv8OnQOUmPKhhO3aVS1h4UuRl/xFR5DpDPc03fMQL
tfvT9sez6rpw0LB8EJOUddbS3rXeGkuwpAoQJl+Mn7RRNoz3Z0u81w7SoyN/fKJehflti3E33N0z
kGcl+6ZAHEJX17Hl2ZYDeDc8xxTJoPDTf/H1GwXK1fCCwSXrOUPSy9eux5Ggh3Z9Ys8hgq7DrGId
+JjIAcI4QGJUvrSeTc1aUCp/P1sWF4O/BepMdKfM3HlInZZdV/Z2VfNxT8i6KReRqJlf+T8VKzYL
RNzLSdCVZb+PURXB1gI6RD8fq1hiMmuzMnoNSDNIaiMRKKUU52576SHymiKG8IA2U6kKuV2ypFJS
8LIFbdHpGsvNCbOLMm0iZPldqqXl7jLPLIi03JjDJz7ozYNj56qTeJX+C+YXtCHfTTOwl6x1kbMW
TvCQoLvshMtsLBsayvNFgpL37CH64ndzIP22iEnTB2t9oQxEpcHIQq4O+DaRmZVizsPwGHB2VS0t
MgSQv1IUdRpxsRpjD224KzD0N8L76a5M1GAjQczpmhWH20NRWy1RGP5lfC5gXPdO/chV92/8nCXK
4cb7FKn28+6hlppKsqTDn44H/P5crO482gHIiNaIBWTyRa03dNsNaMCpO4zonVIqKqL94zE5kx0y
XWYJdPzlHbPd9glmG3DDtK5QPNZf7VSjQ6c2cEi+LYYRFJokPSkJF9voPuFTirEdAl4vMGeo8wnP
+8Nm6CtEjwz/4f0pnyD8YBzUCNQnsV4ycPKqesWzJfNp8uyFaR8CIz0lNpvJsGtpSexl/lZAo9vW
Vy4hFdIs2QyZwPubF6h9b0OGsk+iEXFHObtGUhkjmUkuICfTCU70fJUvkjSkILm+IMWyOpkjHkfJ
l++OneYjbD7W/A2VDCvPAU1w8qhSYpPYu40aGIfGA0mVe5dch4WUdEkuw92pXl5URrHNw33GkcoE
HSJZUEatmKFN6kSy3NP3jcZn5RIV0Y12UXnae9jESuVZJ600dCSo2ZIufJvsd7yJBXd27IalmhKi
wAxHXkYZ96iin68A/6v64q8CMXmUJkPMm7MZEruy4pXdweuMrTjNOeu+nN0b91pA6wHE93FLhDFb
lXPOfWexeboSzoFwm3LJDRueXFB2hNZvA7ZB1b5py4Er39jdWTQ8S6QInkKUKgh62EcvX/t05Grg
8t3+TuI/sKEEO+pV/mxtLYwiwaitQSo2WJGI1D9k6a9bVr6/kNwaBN3ySaztHlJcXu2R+M/6uTMK
LZp/FrkrdU4kstxZAcA54U9cg18Tcr89gzXY1RsAOEtNbscMrqq1zT8qIXntIvyR5HgVt2EGW/AI
9GIrQZ8L6i9RvORZpBrHchuP5SvGG7eNldoE4mhu23tUNN1f5B6Gk2Yi8TkRCq17VynjkZdwNBb9
eSoNrOwvjEFSdfjiQdKEUjSw16z+73m4PA/0E2gBS1aMFangNzyou/nXqHKIRX+1Ut1YBCiijkgJ
pbes+Kyh2b/SLCqmoxWCZzefy8iapZrsiyOEgYW6n6QgEtvimV0Guhe4YEH6klvnN3vyL20dM8fJ
+OXAhm4fLYV03MYgbu3iNtJOCT+NCeOftwJCL7k5f/6ybRP1Kd1DrBdGZE9isEX+ELkgu1ZDmoMC
GHeB/azz4nrX4YS6plr1yDjrWilKqMpgLBJTPPnEbVTLmtzeQ1kpT0iqrBDpzF7wKzrnVOLUDgtT
qlmtI8hc259MnpGBXm366KxS8RhhCmrb4FoWNUp6RV9C2INUuGFvRe5MmGdT2pnzblfKRowKrPa0
6Y3Gzva6eHxnXhEajXRrbjOIQagYpttgdZ7uv+e1WSyNCwquCyCbJYNFEDu7UXbJzdKyszqz6arQ
BH/4YOl2MO8megvfUr6uenL2jylnuiyo/isN/STa6LDlY7NKWwtDefpHDiKbSFUYkLs7vTp2UaVN
XGw5x9npMDqATAvhqDii5X0UXmrK7G2uL7slsBDNfqKygzBtaebat86pAd0K9fywPLnvq/9lXwnh
3S7iw6u9w2aTSyva4dnPKFyvw0xdUbBu8UVa1tlXdRALQRhVLpaeAF0Khco7/HpgrblhtqlBS4Xb
dM+cTJm+ZEOcWyry+dIsCKid6RxvTiVoVGQf2pJmTVB+1Unbu4wmbFk6nwVd7/hpoT+5lF6DeeMj
fSqW2Rn1501V4Wpb7tSDIhDvGH/8vdhQT93b2lhVbjyu02q6Xp+WFb6ipfhk5eYhRAKXNiZtp5/N
if7Vysef5BT8/vcu2rxxQAKRSHnjDaj3q0W+DKLKvmYFuO1tq80O22dT7p0rs8oH7//t9GhVQo9B
HhPhYwCD6HxJcs3xlcpsiLF6cs1H1861GORm8m4cjALLmwYav37Sjywf39n+jtvwF4kyOptycbfH
UOg9dNnjWViCBiUtbXa5sB3tSFIBwoFAg1+gIJoNXZM80RjmQ4KsHNDw3nTbeT38BZm9KdcAMSrz
ecaVynSseR9oyiV83hAep4sUSqtrubmlVIn2zvrmpsEy5aqCq5IVuTYdpHfuJDE9Ic1dMgbmxT2Y
FXlc+hXmZsharLcZAqJxfWbmiEyzRGUH71RfYA425MFFmKPs+CfIf7Ksh3T8d9QG21VKPSwiaYh6
wMbaZEeoZM4/rmZptPUqxFnJAMCfqNq7U2s0QLLbmPe7kBlgTUOoZg3/WwX7wmxvP6t4Va199LSA
njdH7RI3sGWikngiGAkrzq9bwjCC2APV4JxeKHrXvGPBPicqAGZQWYp8IG6NLXew7WDC1T3exJf+
H6vVxjQXfEurrShdaz9GvuUrbGZxpjTu5jQXXt2lCTq3sTbVJDNbfVyS6E3+cxDgZ2IAunrLmdt3
mDPR8YaCpMz3ybDxVXj+m3EiyMux9YdwdPrpAZrR4R5pnwxfAEkDcJlbaGYG3z4ICS9wn1HkbVNp
2LJzpVDAghGVQVzuhkXYDumKpcw0vWq3K/gVQkpMOdPeRTSWMdc5K/OBGk/98c22ytx2v2J7zsYN
SbOhrdP1FJJ3+S7F4kdq2N61mAMbat2H5J9n8hmTlw8QbBA3X0cZwF2EBBqKvBIT5oCS8/zUcOH1
L6/xXoM9jY3Q2XxXPPabi8TLgFRUt/rR/LuhM0nxMJQZTF9Tr9oyFgN8YlUVsGnPE7X7yd706DLp
qVez8ws87nRwFM4seR/Fk6HDHblA3WwAU/eZpfUGOpTSoliaW/zg88NK0pluDget7iu8bFQsT8/9
0ocxSMku9nVRSz2DTWOdLiJPzfRxZ5YB+U56VjsBA412b94XwcvnsPp8pbCgRIAq5EqRHaEIejrL
0dCFUK1UKodWWWUI8kutxz+0EEOYstk0vKOsmsTHtf5B/fT3WszFWWsOO926RIDp1/ExndOPNKea
r40jgo2BQvfR4dTx7QGF72fFMyh1QgbHqq2Oz0kb
`pragma protect end_protected
