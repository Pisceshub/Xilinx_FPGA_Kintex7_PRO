`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19696)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEPMUq4kJG+en0TxirJPL68jVylL9snUGg9S6VQ8CY9jfvrO6CNLVw8sM
mK/bdo4e8Je+HNJtXawm/RtH4YwwP6t1/uL7hUgK036Ykvwo+EbVYQWOFyVX8D//+xqVjVRc3504
+z+2LlvyKRX8ypLFeG75/+gkiqbbH05AZfkVfkf5RgL4e8BE5w4wGR6cRSCzCVBqcGMeRn+CYlrS
0M1fZ/hQI10DV1sJZHMpMW5uDJcmb9H49REH7dzZ7wmsUPAKiN+c5CnZePif/XGehTsIPG2ZmS9c
uvYu91vdnXWCq8dP/HRs2e8LCcxflODoHIencofUmAkx7M2wcejI3wwXkqt49wZl16n6P4xmcypL
gm+9NwDBNWD9xRU0MCf6sa53DvUSzV+3NoV4isC0JcRKfQkXAZj9d/VAqJX2caaHO+j+4wrqXbmN
JdgFyCpDidFasgswOos7uY9xH84LpZgp4q9BXNIf8ctYQG5x2HSTZ6OYNVWT2ZHj3ANEur/hu2Mv
aC4HdTDP4Yg16XxbfBtYDvENKt+Mb/mkhsBK4EA/IdZxnblbQ8gWqIljj0qQSaTVZSnuKpDuFTf8
8J727l+W3isK9wxeDwIV35hKkh2wUlup8Yys/yjpyje87rKJhL8Ph1u7LiP/tS14vkImZL7Xma2n
AXqkHauY2goIq0ujJ8949ktxzbYupxpUcLvGtFividTTklgLUb4PekAJs3v8Rsx5ZNuu13B3dJDl
s5CJEuCI2pWb/OdKRzRxIVq9l+9sWyD/DWFeg/NpoxyXGYqyQYtbWTKdCdGmgKkTo7yC+edHUK+A
m8IRArlWBJjLtRutnddTErOwskXxeSYu9LtbWAj+JnxHi54cAYYz238cn8nv7dAPqFgT1Vj6v/pG
eeCDGTzwmvi0WIUDMA015RrbG+qy/obpMEhBDNU3B5WhNBQVs0S+YO+jbY4ZY7oyEKmMkItfeAeb
Qiqn3aNAG8jaefZUc5/Tr+fJkuMJk7T8oaNQayh1pzCAcUxs0IwGKAA+OFrK4MQD94qFEBg0dyZh
HpJqJDFHu1ZUZ1x8s88XgiwR/RAiD0TjobJH8D3J9IbmZKWI23736A6tyV5BEgB4t0OrYsEMxR/r
xqhYeOosdP0UlF1SXucKzT9YEf7MHzXWVRObBlYnimuIL3wxr73gPj4LzcqBsw+pVTkKnTMmlJUD
a+wxmhhNCrwUL1aiskIIBYd9iVdSVSknEAe91Ib7/joE03Tauo+KCCx7kOIiF6Yo5d5eKE5Ojn0s
4vgflcoVDdGAzvM4Y+zYKEPKkh3ux6TcHMI8pEM80MlFXqNlmcN9h3f2mBKnv9RdNqXWXA0ogFJB
qKAsX+o6YzTClC1qH3fH0Yr5Nkxiw7TH2a75xEf17J4zUmL7tLh1hEBRYEzVlSozx9fjXfWv50vq
5uuPMBD0oh/MCmIco3io+Oyp/UZSGP7HzzVajKUb2+AbgXJE/To2iKdo2gGbjd9I3pYaJDzJV3Rj
iJwzzxLoxaSAi76UKLxrFW7c+gGi89XeQ4nookVXYasBMJ+7FFmt+8Mkz0MWg4PPlCxtj702dI9y
KPc900b/DyLcaRhn27pcEn/ZPc7LFoDoZVlpGxhUDyuhx63k5ed7teGHUugPILk07vjj/ES/6Koy
/ts7JEqYhZKBrPUeXJIBqOWQ0Sxam/ofXzE2qVBjr8kjVbYtp442m5j0cEl0yajJkedHflnQLF2S
iCdE6HlhAaJcE6Plyhqr//AAtNXG0DEfxyRfbWEMwP42Orh5zmhTOMp+Ej+XgXQqtnW/UAP21Bz/
xi+r1jHwTri1LW3U1D+a5xEDoCuq2skAn2A5Sm4fkcBHSzXxU5pkrWlTQ/AShZFEnCjK7qBD6+GP
oPex6haTJgoSTPDkPQQh1AFotEEwAUvVf+TFinW69dlDLzvw7Ao+5E95oCWJodKqshBQiMvkvBZm
W+bsbSuuedlp152GmRX5zVP2rKFubAYI3qvpx7Mf18S4nGOquk/GBMHMsaDBqCvbKNJdW76oxy2p
RrWod2w6ptlGg9KeRAS+VZXWdJxrPuPAyIGBMJQ4cQRfKrqqx6oAOBTzbA64Rwjrobo4HnNlOzcO
c37spzgagZAeP+wT4OWecIs7u3PCS/9FojNfsuHmU8mmASWi4NQeTI6gSYkg5fFNjCTSLrZcR2j/
16CpK3Xl10nhFnUy33gJkMZHHIXF9enZkOSrCG+IbUC4ImvkSOFHBNpcy1fTrTgzEZPC5HoRN3Jm
ZZ55UrdiYHWUyh3Ne/BXBlFOgvDDyVokm4S2G20sVd+DSvXh+h0qhzneoc/n/Ewu5/tqChpKhTNQ
q56FYTyxlY8rpX1qmL3Ze3J5159zJ7X6HKeU0nCuCzrDapxarz84QarrGfh7u9toIfDLKIczqJhz
oLPsaWZJrRdQfnABb3RW8L32T00jAkOS1PYXyk07l8Fm4EsRrz5B4RyKzTDQ/fcdueWQByFM8Oae
n9iEeb9rSdCe2Udz50nQ138n5Lyj2GcmYFANTVGH1WVpKkq41xPtLHVvWUfgkZN2Vix/jLrSP+82
MfOCDbxCcXBMvgBLQz/dqeGwwf8tjfM+vv4mb3rmJaflTIwC09vYVmUynG9bbj62Zj9NMNdIzY7j
gzEXJMxVM2jDP2m1c5R40Dsj2TjvrW6B4HZCHdtDzUA2AiLWp84NC0bcT1x/lyFCO2RNnmy+fvAk
mQuqwqPQ93G29zPS3ROEc21dQ3ToPlwJvimeKy5sMsO/tq4bndxJZfl8howXs4sGm8TdS1ikzwrs
ZgJ4Cw7a2wTm9KlrxZ7SsVforDDatTWcci0iIPAd6hNMtmddaAsG1kN4vkhsXJJh/+xjrmDmJyxY
P1s/cTxOfoMTtY2yXztCC7q+fzlkJNWI233oojx4LY5aPuqOO5jkeWXGHT6vxn3dpsbOXIEWTNfy
EWi6qOSH0R4qoO9rVjq954VnzLIU2pNerQyBw/rIHwrnl0aUHdVZNuBw0MDXoYKVmVrxonLhX1PB
ZJ9lUyVyDBTtlCho9RXTAgy43cobPEP0W9HmPly7FG8XwVheQr/B1Jq6PpM7FcaOemYXdmNlPS1Q
vOezgcXIRVsnxxPM5W3mJka5ONTQaAWrTuB9TeuZM70Z5+jgslGdKQbIJgjvO0TmhX9HxN+0D0cu
B7M0SzYrz9mE0TNvzVszDzyOcKtcr3AhkKDHBAzImvCGm5XOb9tybI/6eZcoXL0IB22YTvRmh2iM
yf2XBLh9dd6hrK1qfWNWQWnOw8p4cQIKj0xfV75ckdPa0redJRXJzfP82eRcfADatsk22d80ReQm
q/ksGr/yYGAiLSmzprjbtnYjWRxlP7/jdHWpFESzNT9uHKXbGaB0pdI3BTouL8TkgnfSEty8sLfu
50lHhyJuV2h6/Uk103Hpdv/V4xvdMpB6T+Dh/3JZL25Yu5gPNB6TJOYVQpeA3bPjudtnJQ1CWdIR
Co8T6M0U7MqSYs4iwAKDl/GNYthvS740aOYkUo5mavlP5WFjui5UJc2V1D+iLFfSPS9L0OBvfAfT
smB+wIUSnPgXH/jK2warJyp3lrk96SDgnTaJvqhOs9n+HPlf1ozLyPdB7J0gPnru29pL+50fS6yP
IF2QfX8kghwz3cvEVcX0b8b3ppNMCrpdh+Z8n+aWglchxs4X4QTn/mJRmIQ0Xd3//CvJH4sTa07t
smx8rPW0ppcMWCMXSeoUW5LD2SrCzR45GmH+jnTle8UcDjENW+0FWLy/QyYDISs4Ad8m8fBM1uqo
A2tb//kJ5Hswwr7TlmMYgv7nAs6Q9Hu9dO1oFK20rmnerwfik1DZ6lpatujxurIfpUOqdFIWQ1u6
uYmDrJNqm7iN+PvoluYYctpmmrTMEbLohUug7C8eiEL6EUEm/uswz+uN/Nzp/zDK0J5Gfj1UBlfO
wZxMzT00Dx4ehTb15oLvjKI9GzMtA6MIaKVt0AwwKpML/7ZSyioD2tHOFXX3krLoZxAxJ5SnTtuH
SQMEOBGxe0YFXh0nn7l5LzMRtu+4g0G4GhQ2/S0q9tWk3TtnDe8Ozxpke3yuGwRtkjbDcldtG4aV
gC1gviAdzTfc1f9/aHGbWQkCvj6v5qyQtQtg8ZPMC2T0jn7TTmH4fZWfGGOefV0qiJ4r5U3lsl5M
bmUyAb8MueIU56omwSlfjfh48KX0cdKJyVleycfw62ddx2ZxNU0DFR1dl+D1OMeKdXMjum99ipoX
kgS3m5jhqb3oF8X7VS7fcb1G0fAVuOo6JpBflMbMf2v0mlGwks8gZlXWy0X/1w6xlzDznl00T7EH
nArHhLDGCgA13K6HujkCKE6t8iCFdbmIcysPFJKYuhpeMEwQFpktCu6irrq/z5WtW3hU6vlJxvlo
UlaQItwL/TI44wNanrfmeuwKmfMJazccoHxnBa0DsjP/GvIuqKXByz/sRez32u/TgbwxEkmIjiuC
WUFFALpK6eOMfdtwej+9YAt7S1MazxwWvrJFeWs1OiQAedSTlth8YgeqWWI/x6O8cJNEcAOo3/HX
LqkOFQ1ZY6+i1sEvGdCbjgO5cGTkCQ4+IDyXQa7MUXUD3srUAgIbxy98V0MBLMWzs42YFB8/dpBr
Vik9kPINhdoxDSi175cUcC+xJnLLYF5kX73snAxGF2P5XQzFl7P7eKxyM9+bhdEhh4z/2UlR/eoQ
qLgMU9ZQpfVnt7sFsZ8ol5CIEGn+MGBuBHeLTNkP3ylXW4B4Ik29vfVc6kIK+/w08azkgvwdcMbb
dmhYPI5Ozn8Zx65y8C3aMzVdVKsG+xLpWFn4/JGAMVWsiaCtqw1cful29n7u7WvO3Le8HyQ01bKq
ZaoHNUsJ6zVFUXLQ60wZFTAfqy040Vo0izZDF7p3v+zJTKCP05LzqZll0sIyp7zcCsBpmU9CU4uD
3IdAcwH6sMp6Vmc5QchfU7kCwa9nvcTQ4uAzYw47FCMYEStemfr/eAbltDy5rgqlv8ZQfsGJBfkn
p5AsEa2/rYVPcLRUUFFaWJdygPZ6Oa+urygPoJxgqZbvh/sic2rzgon7BfXs47fSf5XOxljZX6Mt
73748fTsZb1fvzqgGnt4+9JxkRjHLs1EECpt3v982ISvCA6qjsHbJlR66AXCMFlus9HkFB0DH9MY
+ly8xrqg1OGi7INF8x6pDZXx4RGZ7tv9YosOJSTdhaNS7Mu93IIpNcPHaI7nt/yq5fWrsCpoZzxl
Fp7RFrnFHNhRI/qmNNYVU8XXqAOtUihc/PRZGJ28L7D3Fg/VHAmEy+lVTHMd+YgsAHkpJ/Y05cDJ
mZV3PhDuL6NCbIVuL5SrhBp4u0tjWJZBeCUQVboCLX79LtiIw7opHNyOJtqCbH/fX5EQTbRIFczz
7KXkb9FgiPo14QrKAYDPZ8gk2JqpSesMl0Yj0hFG3aOgj9Lfq0FF0nM7eDRs48Ys4gxHlcHSX9G8
ccGFSYqd230KpJJw571IkzOMU61y9lnJlG1ItJUD/G+Jg9+9NdDkrKzdR1ihEuF1EejI8UOOp4wQ
jZ0JNxpPl9gvo7wLQmzclOo3SwqRTl2bVqz8+fR3tGJ+XHq4nf1PkGeHYeiEb1MtLWrURMmxA9IX
woJClnqaMw9Jyi8E9RrW+aN1tNFSxTbzEb+oj2eWNlRcHuOuOjttP5MuGGrdsoSeDLgkQ2GQznPA
GzE7Edl87y5XcOjjkMPsxw8qlj1Thk7eW7SkDqYmPRkvIUk5qtHT3PZNoot0Tou5lXxJjkl7XY+u
OP3UM6Tw4hI1Xxp3XsiNiHTNIrZNf2bE58Jo8WtkykerfaPuaTYeNcL2g/MGofxG05D9EnB9YEcT
7kzMqVgl48F5LkTfiIDXLtR2vigp099SZP+nWLjx5jhRmYOtCj69EM2ZjVAdaWnsgkCZOcaFZNr+
+WLXEExc4uyo48NXKx09md6upnczcosauo/h4jJAhRY/1x4s4MJtdbqOals1yO4Qtelo8px1icJ+
Q43rGc7CPEUYY0yC2bYsZJ6obvg+FU8W6eRsiz0KAsw8DdU3L24aGjXSldCyXihoJ0bz4Pf0nRIu
Ztqxh/93iX0gCyWc2vbM5CWcyzonDw8zE2dEEwO7Q+0e/JB87q+cOYUbwX3em2TXrGMnxiaBpaSJ
yPs1DtjR9rmZPJSdrNTZPbuySn51kc11o6v1HaWMG42ovgCSmYL724775SXVVBzS2v240kjHS9bx
68Pzy6oNF6th+B+NXla4lZV6qOQSGDJHPALzMsrDY0aaiwVch4rJ1nY+FnGASHyTk7J//VcbCK79
6hh82Tue0jqR/KZBR3UP2PbduVxI9iAVyI+6RMU/uuF6x0RiIJC7BBZsxUVKH06HA3RXc++Y+ft4
IEGF284bO/h+5fOIlEJkkthyKNdSsko3JqqPCB6J8gJR5Ngn0sOTaeqzD0lPrsTT8gqOrtzvlGAX
ZGaPkcbGlUUKJlzNzoXmhJiEYsdfL2X240D0vazrM9kxzpuR6zuZ9gGXGZ1fpUvdW9NO7iZtjtaP
l/oDpptDxJp9eZCYz1qN6UBpHxmUipQnjZqVVtnv3N0WzOTBTphnqu/LINEjEF5AnZATpsq+xZBH
OoawZ4/M7eLQ6F5SMBruOLZaGDwVrrlOwx4soLvPcs0BqxCXo3/he5XuC3KvooRZdIZg4rN2TdNs
OhSFCc4dJ0avpnGmJtriRukKh8W0DyLCfWWQwFt/LA3UK7GJ7mIpNhoRdQL+1x0m9I+41fLpIyfB
eWLdASPLhwJLy/3Dn/CA8NVhdUfSG/jUQ2NUbrv3bxazYF1d6lKz0RuzlyesT4CZvj0KW8ZqWgwY
RxZdFMS7t8+JcUwemkycsu9tInaDswUxxHl9iYZ3SEWNFg0/lGlagb3XWNUz4J40tWWYYb/Yn+mA
bAxKZVYYotgrO9/9mfk2O0RQOJCC7BOqgAwjaUZijr1/kuRr/CZbMhPkngtCIwU4NdCgXq8xUc+8
IA9ahL47CfC4fNS9ExvN6NXXO3zpAInKX0qOO36Eoz305WTPiuhCj+yvZS6hOcSMFFT+2eCvvMf6
NpwcCNQCa4XasUiPnI340swUTgBrNAaMs6eJWy6Oyk8hW4sNIspeXQZ3CspoiyI3qDdcReJtTXWs
wFN+QyjYjvwYUXALpg+/7IlQq9V37JoyVA2opM2VAat0tP9x1yPJciq6skNlkIE1U8eLbLGHBdp1
iaxXYPp6woG5p/oQHFN5+EHOYqURQJHxijPBHX5BsiEqfqX0gdF9CHe70AUfIl/UtbffwfiOoRtO
EkUZ1DQx0yqzmAEExwhthNieVGZgpDkQ3JHrYE0+zv7mF31bACcLR0qur6KyZyn5Jo/mokAFk2fF
DVhxImCoduP1kDwm8sPtJgQ16/LZ+U5ogLpz7zzhCVd/dfey5oMK9MMf6QlDe5sqzzynDSPlxc0l
ht9oIiC50mbwnI3xmmrZbto1Ii7JmmoxMWC1qyUnTVyGXzeUjzjiJ4dFKgUop1/N4locLfmiL3G2
B8dE/bTrK0ffd9eO5Rvu8TOwftUbmbQkfHRdeI/r++6Efzwo0qzsqXoLzOqKKSJqE/1sJxX+96ly
Yn8xdaCZvk4G4mQnECs4ilFkoQnEArihO8xxGki8Ac2gwahN094jLy7R+fU8qsrvYTvVIhgEPHQP
Ndtz3+T+wpL0AkxBtQOAklpgt/u7fSJMjm/i3ifEBX8feODHYzgCduj0U3PlWATTZS2BsD8Hg2ZL
UIhENSCVWOQcfEdXUyxOop7pzls9brevC0WShpVGF9aLhqww2Ngzz7+scCEf8MGaf9jo5c1LlBgw
J08WguqdBnZGkSPC+gud9GWfBrOkojCenHHf92Vh6ILJXT+DxNboRem47w/KqXjYPSueuXC4GP9Y
ix+II0PJLbiwZlXrlmvcqL7hGGACtd+mLOenOPnH4SRbt7Ypeoqk8iND6ul54vpcw6hP+rmerr7s
RzwJs4Ol4BlzsZuxl9uRI4WNsw9mcleHEf7js4h3VyI/jMNt7eYz+wuSL6heZ4y+dfLA//f3styW
GsfoHCDn9VGUE+lPwFPUrSotbgnjQ0kLdPqcf8yYA/uX2mtoQpYW8Z+W2UmlDMkdvzyfi1veCq66
BoUzrQsWmfYQNn76A4C1Hbm8HkOMuVk5dnJQhWsubLdzm07pnRaU0+7O7OXoLH6GZ4+xp299xphO
yeqOxOlboH3PM765m9FiawMvOH/EPXMvtTa2wjcDZadrokCPynHLPheUJlAhQmZXfe6HQNKbr+fD
RFIxBNf9MnURj/oKomkUWUVrSHtAitLQyVWjN7amvzIOjBa1feFUN9PGm1FPNbBDF+jQATIMYz1O
sPWXKmry8rq/WclM7QhaGt1eYmzIqLjfRwGCVMKrKYIw795aWQsajU9csOlEOo3V19biamqTkf1X
2FAOvmz7pEoQf0YwW9YTg8DKEjt86aPUHWsv05/0F2HsYwpOq0CN15Gsq37V7SnSe8gwhwwtY/nT
75HCx3jIrDP1HX1BHuE3DwRHiF5v+gTrN7MZZJLc1Lf2QUs0E9TuT31kh5KoLzQPqryo4gRIfljt
T3w78Ibwmn7faJX6lZlwiRwRIAEPIpuo4FyhrBJawuG86eVWFLe3apI2eNKoNLmABxfrj/YdqSaj
aiArIPu75TKJMiA3R5QPWLCcP7G77jtIPw1numEvXArpcaK6G0bw7vrDPZWBy5rMBNRC57ckxw/H
W9TrVRnG426NKSEmNhB/RkYRa4BVdi5BlBc+6Ihgclgxip+TWf39XmYGXbHT5QzkAB9IoH2PdLGP
MSoFU/nL7TI7cSKRqmsB5jfYELUd31CPi+NeTpUa1vv3dsqjj/6pAr75mJM7GXiBBMlb0cY16t0K
ewIYNU5FcQpiOZhPHBDS69ZgqrxOSR2Zb3gC9IgjSZx4VRau8RCNU6+mlSZNAtBYSxOAadjUdTDm
raQFgCsGs/kvkeMtdSADqmvI83aNab0U8um9ECm9o4ZK7JniXCc/uNvg1VhWmRAtt+eq0md+ZHqj
nc4PexhMtDdbtPMKftUBC7F8spcrqsXPsadJGynj2ngaPj7WfHv4mzjYPXr7MToO17mNh3AIo/ue
xAzxnkXGF1qU0uhfP6UyZSMkgu4gKyTPxRvkzF6AzN5B4sH7rvrPIUj43S7W69cIqd+YB3bIT+/q
UeIiwkvyF+cobbvtBdrL4Iss3TG7zXokKN2faYmze4G9QGBbG2jEzLeizcNHNp4ZoNQ9Xg3/rs5I
IRpegePzyG/T6lCISgivQpGNfF2DizKHtIW33fgJdPf1Kh2OTdWutdg4aLNfM6nlVmkg1imG/b1b
7eCFLV4wZ7gUOJolKEjv+84CM5gimsvYwq0vpSU8dvV2jnMnY73VGxiTykP2ntDtdt3+x3xLBITp
feMJBiV1E3HY/eztVNq3jgUGHUYn15fIsWEauGEWvxWTZlyMMuAvWV7OTEHt3vQub/kfN6R6jbS7
ypN8vcbl94IBXCW/0eTJkQS9/boUVBM2rxNAmWLHJF4GKYErsVHcoX/Zip5RsppORkeEihmvTTgh
IwlijNIi9iF/FcoQg7ZX9r4cVySG+HmRhoUqox5ibYR0faluMtGfbDh5BgglGyeiQ9QPxckLyk3X
0ANuuqtF7jzszbkZy1MoCMWlfv0xQEsPjyn/J2qevxo8vjbCGHn+UH836HduezMYWpvgKNrXw8Mw
4k7pqjDCwFtmgatwjpu5dG4iswIFRwKalyHoTTEFARjpHGYq02xiDRj7R9rCmLv+Y9IRdA62gRKq
JW0bsPv845NLGpQQsTtHU60Jr1XYtiSc5m0pZqGEtnnQ2xCQ5hptjBosCUNGcM8DGh7MnwRiQQLd
WoMeKKl8wkPhalUOs/5Ycik9lChBG2ikMxksA7K+rPj3/kJkcybWhBreEtJWpLfMd/AO4FouWMXD
boUpHaame4o7UpwEWJd4cjfLP5D3XSkBYmOhPj04ZrLHnC4oCtb5LRwhWsdsyer3z0go7I4Jrgh+
pWuoLy+kfSqC3Jlt4R068wNtapQqKO0j/pmN+wxl2rNPgZ5r7+AbnPUxfxGquw//72n25Nfb78tj
x462Wg+s03gtW7B2NQOA7QXgmIsB7BXcg9kKtKR234diigIlYvMY9r3/XQZcYmz2PcPKv+TrOAFU
6tc1McwX+VYH0WH2CtcPZ4HUTHSUqJFBsXMMSHid63G5yA1G9jEED+u6jh9+8Y5wvmu83pH7VXpn
hXu8liqU4BafoAJQvxQe6POd/Wko3ufSHOjEnz6hun57/KZG0LMNkwfKpl1mqctnJAwT0MF3S6tz
Hi7uguCPYpm/S57MhJuJ9kVieE+H5MSyBn7pB9ZGyhTh5ckuxQtLm3MX+NoB7hrTsVSKU+Bfyvtj
HQQFPt5dFlaPXnlOElMS9GYB1VYNB8MbBAH54VtmMUDapvjskNmxCOC5DwiD4JcngtZseSS5Rx9z
3mrWldBNNzd30HbFg7fCgzFPSKVshlpcshWzhc+bsydqSVOgPCSmfVOt+1pInWNdVyLnJGsyBchR
x+MWfCOTAQxf2OvSp6UZVQk0NLs3lZbLjesURorFhxcW9JujxEhf3fKbptsbKp/236mwrvIh7dUe
1COJhHWkZv/q++U2NZLwI7XcSozCE4JvWW5yVtYbcm3mTnhbS9EZz8zng/3Rrqj/uGutWI/fmf8k
K4zpgbj9DOgrPGq5cxGXPAo45GuHITJ7nDju95887elkccKwPfubCXVYL38RDQfchhzFmFOCOB6M
SczgFksQJ7aaApOKZY8WEjhoKkBaEDDHqb5Jk6Kl6V9HGx+yC7S86x8Jn7NctOOcVLepytmLALmX
CpNQCJqf8WDfk0M4QZbDA0uZvojkQCqibSa0uXyRtUAB3sfAMYIzZ/klrKF+iuVr25VJm/MwSu/s
unPcGYtDREmau+DhmfVlbuEzN5GibOyCw1yomOHfymoqUpet8AAZjorKrACqMSj2j11BdBLAxv8R
dI4vqOfNEGvtcFBOigx9y6jEysHbkAMJZ7cjMoycXcQhi5sWFGwSrhdbxMPFt8A8oq49pgOIO5bO
SWQivn9m7h1pCQyLdCK1ZtUHY2JTp6RocFlsyBTyNmkhpB8TOPjayxFIBWqraEvXGXY+F0AbYD9W
VLRM3xnZxYXylwENT8cGBcH/GY1L7jVqQuPo1zUjdJsi8YHwYdlrQHbZgLBZyuOdEJvgbaedol1I
Ykb2oEzsR3yQhu54eraLlIf/cpdKD9WNUEisOkJSfAEcxIqpzm5iyoM/ZhuystqivC+SE9TIlZTL
8S3HiRKkDSepT+yNJbmSlFWwcFtSQ7awoOlSpB+3eYAyaWxs/T4ZHSAUksFMtYRdBfGp/8Z+jZqo
8PRDMXhJWFO9ScChjyJZtlSFa/qCTvJHgoYCS3tTri30Wv4USQuGQEKySXv141uTQWPHEwFfPrdo
cviFrC/tUo0aLrP5sJeuCcuOwaHYvko95zJlL4UfB9kJfrDhfi6eUPRg6AhSe7qiN++7WKHhDDBS
yXpY5VXhOgyl2ZBedUP27HPizKe/GT807VO2zOkzZ0yyUbKr3XB+ZsCYTbn7YpMqlPXCpJn3NDkE
zhe9WXGXKt26B6fWnKmb8ajcwL/dkRNI8+4ARyhcp/XGLWZCvPGEMXuozlzEPtPDLHEJ0SzUaLiY
ILLBcjww07gEPzoor+QYq0vNujU7YcI+kpjZEj+13tTKW9/UwcNRcA0dNT1mjIxG9ufZ9bCsHf49
151wOtoWwHqqVT6lu0z2geVMQ6D5F1z1E/Bu2OVbJwMgvjiklk6TJUokJmSlFmjtNx3nQnsJWfhi
id7cY4tG9mOsKKgf+mvlDERPLP+Jvy55bn2ywv01o6P7tsrxpMCiBkLWQbcG3IQaKqGLr3Zs3VL9
zdkla6ra1IcbcAZCQVFlOhK9ciSgNcIo1US/ion2eiXtaoQhqnD4N6SzOMFVO0uwboUud6oxtWWx
vVY2G6pR+auK9GCfV+Lkydd944c/4S1lGB3XtD+45HkVmWeEcj8j0ZNou/3Icjh0a4Avee1N/hXd
Y5sgXUHVrztGpTeCSFjjBusv5TaiZ477eEL4RxktJNXfU3m5MiN2zd//Je5nyYrRxQ28Ut7n19Ji
vh8xNr5yAFiEeUlbJy0CVfGxa83Rn0ub7r5nUrV4muPILw5CoIPpu/zbSLWfJYf9aPpYjO8t/hBu
udZeVblNhBPqMts7IOg35sjHUCXdDjkELookENmoEdBTSCdO9YK4AllwomaM9QidNvr10iMRSpqB
0rix8KEXiE0VjfY9tYINt7u0LimOTrn/0F2RKxTugzDnFhOubXewSzVZ1+KQHvOAli/qpCcB5+2X
ElOS6wXoTzzZJTIybxhHefbcwRzLCryRVmDpMB4bn20kXYUEsVTrHhaAzhOctzVcf136MgkxOHB5
gchc8RXJhLTMCl/VM2g18GY6WhovbKtEGCxBv7YUwtHj86+c8+QyQis49AQIglYJm4W4u2ynOm4B
xLXaDD/0oG2YcTfhs2Xw+u65//RXhwXdwOnYLTA9We3OOzePyOzRivMMnsy6T6+qufvFoY6x2DmZ
3Va734vAYOf/VJxZmjCR5mQg7uaZ3G+Wkim5w+C6t94UVxFQbUEzu6xQH9pInDu/6ZWQKHaBv8Fy
jsfOlkTJENEJyESRlIDiMeqb0RlbLhQudlxegLb6lY/hIbKB0PClkjfVSy2s/FSxnC5FFyXp+TVt
y2tf4AgSi2PZPqMs18HOabzeUtJl6w8ko9tKcLL88e6csHKLBIPn+XdxfVyVMoq9jmRXNmwVYXuj
4Jf5y8lYEe44uejDp4rhi2EDpmks2/0pndGqAtRsbcpB+jQw0mxoAukjQpxVzbA24lTHlyOoO8GV
upkMU2Ntw0zdndP0yNkFdN/ZmtZje2+dzW1IQkdLA0Zs10L5Acjq1FwuJR1G8gXDJR7kqpTqsxL6
up7Zctmb55BAw3fTcKynOceGDzPdR/J/c8oMD9eV4GlSld3wiuRtEMxGap7wRBDjLaika9jDpSRx
5fLZ73Jh9A2LtGDxHjtTIA6MOTfZu+buFVaRgkXaaT1Hjy6/bPloB0UqFEGobHsoL5Bzd7uyxys6
U2ztNKc8PiCcPuHGaqE+TxJmh65MsGLt+2GQFE55ailu7GsjgfdeatQU3Rq+cwCmVx9Snd6fJEQY
P4ev/OqJxyX6wlJor7JezO0qUoefPaDb0BcK3GurRlmiq0ibLxAMpO7U5IWpxUvhi7BDTSA+M7aV
xKBMtf6YHWO0VibqzUwDpeMRrRSAbRnzR+FrgD+bg0UWQDWkb4BZ2vpR6VulHoQ4+JF8L9Nnq/ik
1tRtaEtTY97I9YWikcOAqX5+jAsbVqNnWLVUQaoJxvbrwmi2cZoe3NoS6GHV602uIfNC8NRN/uDs
Omb4QzT8e8id/7u6J1RpQ8E4EgItJoRd4IjY3LmUKUsBAdfjBdrv2AQ4Xugh8yIoVLYt+wiRgZ7T
dGRgDsWIazk72fuDNXqgZXyxKcnXEnU1NrgF4GtxKep3kL1G3ZZ0P3wReV6I/ul7zq/Sib6HxxYf
N6F4Ccptp7D/bgj6Q4o3cbaondAUQ2pINR7NwCHD+Zl36oAP6p4Tp1bYhj50rk8mFBbxqubCAzxg
290bReYLUtZu5s4WYznwvssjP5Lk+IKTFyMI319IIYzl/ATB6s1yLKLFSlBqa20mips/X8V3O9a6
hSIoL+9wsnOAooQL4b4LsHv2WZq0teTVts8Xk6IXC2UnZXG9hOAYSxcLh72rTu78kXaKKNlIf1sh
EEb872dVO2Bl9upWqnqaVOrkxZVDaB5Hv0RqJLtZgV3alRuSpnwnjSJFQQO+SewvtIb41lzBxsow
KFnjiC8Q0ixs/NuBqfcD41WE0gzG3tWwNXA+HivkY17q2XSzmRLAFAAQ8juV/HYH98Wa8SinnjKQ
6R5eFClk6cJ4J5fCQwUUtM0+2Kxh66ws5/k4Bc61Vk6hF2GHK9wS1+YYVKAVn2Sc6rKm/iize590
PXtH8GBcZAcH9SvBt4a8EAsmblgser4KVgCfm00isw1viQ92EEHEKufOHbDffRvsUlGUCz5q94x/
cZ5zCYtZrGjS2FHw/or9KarucGaTLcrZ7LLxrZCjR+NJLteobpR02ZMg5XWuFgjzCoi3qVlSKXA8
5Clw+IWalKfIErJTRwDh2vlzENMB/EV/I5fcirpIKY6f+Ay5Kvn5C3cSN3vwYMQOLbspRV2wZdtm
rPIWOKmWyCRRbl3v7oO74zIzOhHZXjl1wNbBW5smiEB63KNMWDZIxJwWjYeUmd27w/sutFtuXHRx
TcK7R/1oR2UFZJFwrIE46Jdfo5eJIn3aD1rsWtO21BclkdqIG+ZPyJ8zdMEEV1lq4d2L2OskyuYL
RX6UefGDQKuLgbkUyDMNgTPcp/mZpbgGEzfL5inSfvW5h0evkQwhAB2+OoYqt+RhUbqrnmMMZ+bA
HmGn17/r8dUFMGFXUfdHJDNIo07VzrOecOc1fxAOTG41Jorlp89rrFBAqI7IaoJM16BVYPzNmT6k
1H6NCau61ehuUF5UpDb/RPEEMat2uLa1U7omDPpIPCxpTqcE1MO3R1fJzuhQw7IFUx0bTW+Knd3c
yhxF18u+Z7nQ/jxdtuf6i3SyO3N6uIwIQCJGuBZvQ3KkCVVHweylb1gTGZyYt/3H2lfISDOOweyl
nAsZBDKmKLUP2kpcwAZB+cfcwdsMA7o5Fjwv90y20cF1yz6uLADMIESaMEt6Ni9E0TELMZ4XrD2A
3boNqfbCfAvWRQJ38Jc/Gzwn6T7l+X3yqLq4dBpA8ZK687NSnsWEyqD5UeFG/oLi5Cfux01239x6
fZa46ZQUKWkrgUjsUQRwZxGeufCLc8N8W9j68S48TL7j09bZPMwPneqeKDfMBD39YiVh11TxSMOc
4a7RS1jMOY72NM/di18r7u7LCRKnWw4OGe6KERGXpKS/BDRtav+kdnVyD3oEjaA5LS0gRNKJawUA
fvx1FrLKFUPRwz2fkHIKDiaym71J1xW3ATBCwEHbyk69fzPYxfdF5yneaSixY/BYJPelMsVmhhNJ
iP4AMln3PrNPlxSB7JN2dYYHQ4ogFU+TQF5kTslSfRga0sOAMWbS720gIZHtNg2zUkZ/1rv3iDmn
3muameIYmKzWg4LEst/XcpZ565YubzS3ZI+br3MunX9R2XlqLB+ezzpjnndHWR4D2jX0ryZU/sWI
al7rNMNDNd6NGrz+Aa4IqAoYvi1D9rLL4BcZuk1AqkF9cA34IDtZl73QFmTT3cDzoPGGwECEaz2g
1MuD0tYMSj+mSSMmdjQ7p6rDNQSdruVo1RXEbUekitLyMvPzzIpolCDKSNzzeLHro9hqILfys+f4
k37wF3m82ibSe5Q2wnb7G4woPm+YClCkpPGUA47WgbvTnTbXQvgjIuFsF7MaQkVzdvpsmyveW1zt
IFhDuYAGEAnrq+sl/JtK/XnF6Q+9YdWTyAkelWLvJw5lRl3ghaJN6OKFdExU+l3/mhAzNG1SfQCv
QjYowumhF3cGfkkUguJHOPBVEFaP7clq8M6iGO0hTtJ5divUBgYuGY9WaAofyk8SBClfLZ56o8FO
wYHL6lrFnw+Onaazeo23zTaAnMb3wM7ifkEyK+iGj2t5tdGLZwVx3rHk0PKZv4oxmxeklvDNS9+M
WcRqkBq9mF8Ze9tTjeTr0wzvLl8RwzL0vYy/CYlL7LT/gtHsXHIhfLxe9qVQYqazVIo3SVc9LJfY
l9UJVLL3yfT3OaHBBIwcM8L1kIxCsxerNupD0Tsu4dKM8cMgJ/+jFp5UGyN76xILz1YzAsb1QmAX
LuRsxgUUIB4Xzl1XabN6duap54hYHFNQfBitGvmjyJqZvfzYF+PV1xYomplnG2+58flLo3SKGYFV
3hkO4JDPfL2KjogFfBv0BP/mwt0hV6JiWh2WoQsVRznNTAFLRD5JaIgqwnNuM43pIWPAEPXPV58d
cCOBmu7PlrX0v6wtHGg3MwykIViMTDSxWY/wLFsmLxKdnyxy/he8+9x69A/lP/fcl3L8QaamvPT4
uS8wDjbnt8BW2yqaEqc/2sJs88vtNSu8EXBJh2tVkzz13Qu70j0HcWZRQ91Kf3hRqo9G+ppCAve3
fE/gkakmk90fzPYyisB047W4yL/ub+TPYdy5/qTqPsiqnY2/VjgoyvyYF5ZgoLfh4C9v1YOGJogp
bVJSbIf0uYAH0LQyp6DPQInBMhztwPGnqkD2l/FEl6/2v1WmOKM0WngSyUvGTe3Lo+ZUX0dhFLVl
Pbn1ARmoD40z1LFBpG0jQAg2BAxw5hHdee0darXuIl0meTwXQvTtXXbDB+YkrhuvmySdsikntgRm
WYplxy27EXkMkKMp/UwLT+OM6puTZP2OMdTgbW/jyf9gwny+bCkVWDdSgBhavq6kG7X4/KxUNwMn
JdePmIl+GSEiBFOMwAaXfOFFCZVcDI9X03XvpRgYOHABn9CJNya7+UfFx1acG1NwAgYLeUEwGzC0
mA2gBtYUJr83ETpPGVY3IEQkqYohLh5TypBOpkOyW5xB1/0nTlejPpXl5DPCABu+jB8QToeAH2yL
Lhlabo8MMWMbJSafxrIHZWm4cb+v9HwIBOuKidn5n2Ju0Y17bOWMlvQHr2/EeNBEWShQ+xDfIC+s
+MUyDo/lO50Hffu7oVjqTnqtZ1T4uEKkYBnyp3PgPyXB6D8fZb93/djhZHDQQnsFigX3YhgLrs0F
HMzYOdpL6nNq9y0hreteMa6XrZPV7VNNVgqdZZtSENF2cK1iKtTEwsbrbCXSmAh4uO+MGmcn6Eum
iEFVMcu1VLHxIBRae9yt0c+JwX8v/ATcy6GxDbFUz0pehZDLbv9qS5R/nO5JFuGwV+BTKKlfldR7
IlD2UzRbO8VUtw1aLZzDEC/8tgzpUzNCeuNl4Lv8HK4eojKYHFHOYMvKKIQDhGx+PMODqHnWz894
4i5jlePw1v9JP7M/St1GawS2OZtdYWgkxcWEjZgl2V0BkQHdzCVpJNzBcb9+Tz+YXIYWO9sDJddO
XucyAdVE6tJ9v5ZHZ1oFYhLFy1FinaPO31+MSMa59QABK391MvlnyqksBUw4IdUBwuED0DWJ07N4
aNE/s0+84iWkCbSnWJX8kXZiGpqsZCcPvgs7S00vQZ7OdImDChwwjt8OM3dKOH4BNbaYAvCRWppI
dIS/VPQqcW2lj1/kNPT0Ivazx/7TjTKQBB1pAQukWxQFLro5VP9Ovu2p4kjZomLTrxMQIEz7MI8Y
etHyqa1wOrYj7qTkep+OGjwdmBloxlQKEYqc4UyeTgt5xwvQIfpCRp4z7lsD1Vm22R46C6sKSyNZ
gQ+8nwnvyBZrcp3j1Uy4L2f0iuWarYqgfCBLW4KzYMJbzyA0NnY/0FchrgfSNe/VVhhjbA20Usgz
u/YNyODwW1AVxcoilWw3auXdCvdnBLdckttRpYX/nIzueEd9AlJIdlo129ge+98Gr3VtGkImqo3v
Nkn/LJEHuFvpoO6EVa/Duq2MUhkwuHP8mU+8SD2AfdFf3jenCH/SFn2efCU9fQjGN/tuusgUARuM
3+3D5/83D+XouXjoyzDZooesTX+CXSuX/jmGnD6GVKwI+2cbV1YaGqlnC02VFPYWiImeMCfOpH8Y
Ix/AhFr4P9BQzGTV3/7mAv1paHwAV7kQ+CbCX/S1Zq2JtUaNYJJr34WJlpD7VcbHdbI1s4xWBr9t
zOr03szQewYXNIs2QBjJ8TMS8d5Fi8yqcIjUdKa4WAccrOCG6nfDSoznhJeE8Jm7AB4nkVugzmDp
cYNU7kRdWi/FRa8OFGzbp6qSG0HEFKTnYUy8Sf9SWGg6J33QuliRTHslRJ05FwAWfCYHoWcGe8II
WVgEnLi5O5Sq4sTfSEQxTXizu2anaqp0zyad2ok140sRKcAnONUMigJmkLny4bKpHfOIXwF3EhgV
6EkceXc7N0ClNcE+HC9qu+/x7IkyifankPjYWNHGH4pDU1yvOCg8cPjY20QdUGtJnsJR2MfeaEtJ
fYZOzIUT9jfvo9A0uSJEYSOOFFv29WpUPfK/r52vg7YL8K2VdIOfZ1wTQWHxSBWnR/Bs/V0uc4QH
20DvVgQ35i2FaA+uJ3nRSPRBh1vxiQoLFMWigyWFDrpWKlMKDsCADbT63pb9mU4PoBbPc2lb2SwP
TmmzxIONXN5zf30YPmkmSmlLWYABeWCNUDGsyWWncHgk5gj5B4c5RSMicmGUb3VF8byIZVeFdU+X
JuTFK8FVZcYB0U/YBTIoZo1qu37SHZ73I44wl/bp4zU8eZJIfkqHICTq54EFxnV6ud1LK21r87mp
QwyyruKbES8a1R/00FGD+QXu0u2vaH5Y3K9EQnbAjmGOmWpyTy0gT1H+7hvwmbtWnx4052FzAVW+
Z7PcY3nCJfvmlq4+3vqnhN0gCcIzxpSg9By/8V1W1avxSctailmoiyT6rtimcCrVMeSLGR4fh7bo
nlVhKuUsJs+u2ffDknkcI9eaJJSb4JXFMijLf7UNtWts20TQ/d4m6NqgyWGmYB2FjGZwmVSBZjqG
D1yKJxnM8ig40iYnIvddfvVICHSjUGJCvBgfeodViuHDdlyQxC0yb73mjHTJYEhJeLNOReOOEUMV
GSb2VNKC6r/A3C8R2rlF0CZhWy3deQq4mj7XTh+ccHEGc2Fnl879+Gi82O7K+HD635+sQoHQ3bmv
rWWWZ1Hkwg4bGihxugHejVTzR/kowRUcnh08Nzosltb/qcoAZVeIpYBoACRWjObtJe+ye5C5Hvg8
Jt/1Pac/S2vozegGHVH8lr6TfcJCrNOMYkH7clVf3xnpaGZ9pXPsyIASGxuO0M3eWj2ImJavkO6m
Qp/zHDqoAdDjVCqBtBKWFBDN4+IiR99wu3U2r3v2xT3CTCRPLrJxmnuPwfEySSL4WP1OzsGIGSy2
ByXqkC0Go/NyMkI6mcSX+o7Kvhlx/oU+NNkd5jjIcHEWUqXrpVR5QesKwmqawVZ7AjuIqxW90uUq
J5529snL1yfKvsIanLMNBFXqUBw8fNWl5QuHvSrK1Xs1MbwFjwuEHWk60oQ2Pr2uffF2KM7aypCY
T3j20FctNMfuWQqJaig9jQWdhu4urPrK+Cglj5i513ImMrQRAqIet832s2+MN+szAa9YzDKrhLkN
Q4xiggU11zGtgnXbuuQLl/EG49sBfHZPGltEL0rZvkUQv5rTgoG3MNNul+2uUhAPcdWDVSU1U53J
IQPhLIdBfNfUaGuYtUIMnzARbz6VGfdm9krxMlQHwa9bBjcdUvM/GyIQekHTAFsCT79xxg8rChku
4yLH3NX6cQ3tBM7CUydevEb5W8RFgAh/M+ZtCVjnVA4udfmGyksbKIZ+vtPCzUIdl35A1Uo7AD3+
1ksfdmJXwod0sehOI2WjXQHPojpbbiMGMfMZAkwdt4L1xzC1pFnxuL60ebLgIZgXXKg139eZwbd3
jPvt215uB7tlaD7++p625C6f7iUqVdNwjFuAvUpcm+Iyn+G1iW5NkMrEhWOkDZZMYBBvIazSIhYa
/6dyWOooZNxoRelrci/KaYE6YFe22MCmKMtbMK984MFxrtCRrDfn0LDCl4kjhNIYakKwMVY1GuuD
25YRLRcGaZ8/jEs0qKneOUg7DaqHLm/SrpqUKgU5D48+YHXTdQFHHuQIenauE7qbWtwwouWp1Gq6
3R9s8N2FU9DucD+gpENmp/EET+AevAvt7GdhDQQDf0GdmiV4MpHm/0OFoae4ZAeg3KUvWiTbKqc1
Tr/EIXEXLr1znYzW5KnTP1IYzxePoLUkT52Bhi7p2cXOxhrVoyQdVxxVmo4eCEZif5u3o4xjGsHJ
gDH6S3UEMORQw65CmjoKkF1sAzgpo6ObpjTUTaaIG9ZGmbygcQcpvw3m6U25PrUkD8o7JRvIUdeC
9YrwH2n55rc2W1rhir+LStzsK7gvqEILVu+XJIioId0VH+ezmvok/cyVsgzBglGtVOXTjHTPIMS6
/ucn+45Yy23EGQuFuXt6egGc0WkWmVJ/gDf354245sRtFlo+f67I403Os2lgubM1rYur3wXJ3I16
u++eG5Ec4QgD/JT7d4Bq4SnafpXEFO2XIz4RZsha6ril/epbW3idlzqNbROCIXEyPGGiuOUTr3LK
85U09SHY9BKDe/ad1d9Mddui+ChX93cji2zkWWgpUQG7Tm0lzSjTkb1p6eNqNtRXVTDAVeNNd9+i
Jss5IVk2lYCqKrPMmr1qX66Nf6aqfk0jhO/MWrOZ3Kp5GbuMQHyEaYp2+bMIvGsUgZxEZ2QsxMH7
aNlMDr2U8f1PXD02VB2ZClafZX0LVkiefesqdJGpdPU84Ym5SKwm8PHz4v6o2u/U9i4YkXhXT0lN
M/Qcge6IOORjSfxWR2Tu6ObNtu873Odotv9Qv19jVqEToGxwqlhuecp0suLoicaNXzYGRdU9G1A5
BBLHe5WG3ex+FP6cHI5eMgJ917ezGPL22ahHp8N/7IIK7paSMEETNC47GIpmRuFNHSqNKQi1Df7l
Lnoxn731m8a3BLmJsOLi+bPdXY6N8A7YTsiSmdzsVUZEQ4PGq4ktCoumNltJfwxLUjj5R5SKHquM
5kAiyt2+qFndbw+dza8nvgwCyEwiCSfvJeiy9GuG6msTHJH2aAxrXrAPUxkuqNUBmHEdTLx3YNZ0
P8PzkXgOQoS/QLTu8iJgn7je8JqGKII6VuR9mrZpJ00BCXnDe0v94KqwynbqgjHEg75R5Kx1+J0a
qjrnhifeYnoACpbaHqKDSptkNxMS9ePvEu1uH+T6dsklkWbs3w1vkwT3k7p/c83SbQ6tVRnX804P
wmCzXqL+l7qXaMfwAyG6eg9pcHFsYCajUY9WTXg7DXoojg7gezrEc1kjWR8EM/nbWoi5TYCy/CpE
jm+I8W+Z8NtRTgg54J7SQCqvqJ8G/2x0H12/zcZG1ApqJOhLwPkLrhOrNLHAW5IgZZX7B239rM+h
Ar3f6bhygwWk7yWLqTv8d9tlTd4VOer43i9U5313+m7l7jwKPUKfpbxjbRA3S7369MZtvG+R7ZPW
OiqXvds1erdX+hnQGV9NdGjwgW3EA82fpbM0SLn8s4cxbVkLCbpF6+tjFeoPi9t/9z29SpfJ1vub
3JFbkenxqkiXf/UB7ipk2k8oYX+hgJiCu3/DSm5EFe07CdgzVPQsJqllHoRoM96lWb+7aI1Sy83X
E8HIgvvLT1DSXBYzq9otvIi+sNlDQ+uoqbB+dmNiqUJiZk3VoY8EdJ77qXoaWWWqOHOqNwBKP2Mg
3pa0jD2YufDhQZEx61bMTnPM328ZAvg3i6Fapg/2e1tJmOpjehFvM/hNlX4Nf0x9ic0CnmPEklI+
t55ox1hfdnPAhNhJGJrCXFZ/saL5gw2LN3FJBKBZmHazSxujW354Hbg7oUVHcb8CV4wBILa7sYwk
z6uSGeZm6zz3EiA4IM7hfb/qjoMpE1KvuwEBNcrmtyyyOV5e6xqsGxYaUr5TGNAehf9mE3lYWgim
4cSUGwQpvbUIm57UIKESqzMcGlgskWDxQTR3fEkdEgI6oGGKOL8MIlklVKi6RubGru31N7qbmn2p
VqmQH8lHBHkqlG1XEXUMSSVwxa+gJq8rlQNhwd07A4aUUARdF23TNocrX+DTEXASWI+MhNgZiP2i
wf+2X4diCU1CPPfEGphbQZl3a2Gtn9MU0ukzhGEfPsUR+J+ILTHoQm8hHW2wg49yWfELEE941q/b
nY6g5KR/7yQIOXgnjHK1mismF1JBxd8ARHMgPaP4oaNfrT6KtpohmMgv8VUJqMXWjnt+AHjisjN1
LjEZ1xjWXlCwaNpZyPrkB3qadwWsoiUZLM2C0fn7NP4mW3+HYHlGtwiM1SZ5i9Eetb7OAl4/GlKT
x8W1sH9qBdNKDcqCQMeUqNDieCbQFG5mgN07t6xpGaXeIZ1++EfXULs/Q2Uoh5FcDNxFFYpINLIf
JHhMZ3ziSldzBscsBU5OFy74ubRE0gW2bkXBmu8oflsvexoSz/mW7smtoH8+dY/In4fDnQshzoZF
/W/+eUVcdY6VJNpOxHAHwDEBRXRX55lZrK9mjRHZS6xJLCS53mz6Ysz12CewgbtxdgH5Rcjd3Zqu
1TEE93lqTz/vv5yFSl9swGe9uxmCAvneKXqpVZQGvq9Q2sh6pTbSiISj5+QGGNYJauJVPuPlWp4C
DQH6h6sbo6kyw5mzOdy7bm1b0DeNrU9IIthWcOSANnO/rIjvmL5QD8w3FJ7R8nrWL8fhvGF1s9WZ
WnfimzqKHH27Rqn1IolUgV27EL48Jib5EJR9zPWVhPsHEpAXFyX8Y1H9PV6ZhwnBY26hUZ1Rh1DQ
XnjuO4DgMs4mUdkz26jZv/bid+ObFpKpyH7dHrcqq+vDw8uaERFkHrd6ELraLprCGNEfErfl3fQ/
7zLDZW/aK7wcKMycKsT01UzmcKBSZtXrfqrUIfnWOBytTUTY8/ZRTDDauA255VZH+jN6CK71Szab
xuMrPCz7myAkeWC3ZQDGGlqW18OMG/VdYuR6YaKEvKUuXHs96nc1aolfMdISXGZToeIqmXEhyy1R
qAi8kbp8+M0Jg0Y0Av/6J89olDpnu9yTnewLf4V0VPPpLJUl26S9VLx4x7Zny8Lfg30dwHkxM4Fe
Tzm9BKvHHHFwx23fsyKKckp/fMCkSMFURgP9HwRyUrYcc3ymNgNZfQpJClS2xnlHf2/Jfx1ig7r5
EPyLDEJ5uNC0sInCxPV5R/xskizZS2D4bvvDzlQYvYT1iDatMYlX2rJRhY8wWOTq/nMCpMdUtYp5
KmRAyyOkRtYcyWjJZNTHV/nxaZf8R7WwXnIUCJfsMWdOkvCpuvoKtk7D6DsKpXnTAvmSiq9muFl/
Y+MmOtUcp9ALqo5RzU2sqvApbzkanLRgulz/WSuqsJvrebTg0GIysIb7w25zOQikIzbajl1IiEp1
ryZ4yao8uSE0YOl+CGUrXIxRZpXFbP5yhrmB4eD+fk60wQXg/mpyjKyKksnPpgvUnXY0XaLAYUQ5
CiiKb0rquCNdhIJcW6BBXMLRUGi+4G5WJJIDxi3KZBhx95t9CEgQ5IBccW6MbtXbojIYfhk+KOXM
/ZSe4Z0ZPBtzAwr9e1MOVanH4NlVEG6K55iHhSDt3lbtggm00H1DqjVBc0J0/88JgOOw5319qfxk
I0dGP4v1EXqQDyHZBhoxkbmCHg0okqIEKo/CEM+Yfuga5NLGPEIwjrqy8qJh+d4iEwrgsK3v4Pq0
h4NnJhS/onC/6IJWTed6BezYdFBcqMFyI4GTP/k4Eh9Qqb/iEE6k8b2Gk4HHxZ2LcRHx7nEph4w7
OxF4/ZutDLgDfBE09cTr2O6B2vQPq4d5Y6omOXhgXJW1SVH1KR/FqTqQmKpQzwQHDVlFvyvVSjSA
MW9zdSjN8nX3up6awN5HBXlorAR1weLM31SghrXsDoivLqmHvJZSWyi+e6YMde5Xc/l4Ks1NQ35u
GD7zBKC1ZG13RKdUo5BuoEVHG8tSeaAkFA6jCjbk6nUbC76uhFdnaFJNYl2rPN+xcAt7fSbL2Jmr
8JGI6oufh7rLBlPXe7LOk8NzgoKnEdjeh3oXotSJaIB1SvMF+afanpfiHtuycFUak3m0Bcg9DLb+
fnMALHjJahVZvTmu5a/MNAip34A/CM2aq6rfQZLbxf+yv3q4sznxCk24/8hg9oh3szqIWanoVgEL
+LKuHJ1J3ymN6XNvhktWX6/I4WNG5gPQD0+UsgW2x0p4uSzBsdcZqWA/AqUgrWq/D5XGjnuCx7ED
m0KZLhDgKQbOn96pr+KjcfH9WfojsHIgcQ0uHmzGioUfbAZXsy1ixviFWQvlzb9WEQoUj7cP2M1M
WDrL6ZrPr6zT6asI/AvU7lArhil1LH9sza6lyinxekJ5P4T2KzhCtZLUqO7y19e2EktgJZHtDw82
aWVkncTZ5oxD4CK/2ys9gfEKl8kPWRe92fi95UMPOXQCW/zkz3bjYWAJo5BCQGYfiavOfnZybRxK
Lx98NodT3txHKn8Q3oHPFW88akUYLL28ijj9GsiWOU1FhuPq9Gw8cXTYOvPBxIAT8YiYziAH7icS
Hg5Hd8qydgLr/wtJqwVDUYoD3xW0ddbuG6FLLcKraNH18w0+ZExz8JJzUvaEqo/2/eOejgzB8k5T
MwZ/zdEHIUO6px2Z5PN+kDQ46Z061x+l9vXgOzGCSGy7i1c2t64uzeKjfwT9Mdj23h1nvJmJGJde
W+WTCKkts+KHAtyIYpULzymH9dwHzhTh/HevtIo0bR0uLoAwLWAB+cUfS0ej6gWxc3f+H8f3mw5Z
4cYgS+wlJNlJGsNyyS0BCppDRMVOxZVus7q1cQR9q7I/+USWu0Cn51aiBmKupK9JIXclrwGjQxKi
XzS7e2/Fwu2Q5FwK+wb2JbMEJHUHfhxPuvQMO5gV+qrSoSM4hCibzAfeqA+mrJXmclHC2Vsxq+c6
Dba0QqYg2DVhAdkA4zbo2upjWnqWMjFZWxlexGCp7luaUQdyvrNMoTdzQtsx/DTkGa9kjemP2wqs
b23tqMHDsEsA5Eqqda++HoM5TTgjAucTkNuzohOc8BP82CHsqtqB5tDXQdJgukOi9jS/TAVsYcB7
eUxXlP3DqUmvOeW5i7Z7ahhTsWxgBFkBLD8hOyBZTQRqAO9AHGLb97YVNgq7VvwzRB695d07E2ES
wzEiSpPAZr0R370geUmE70iHTtwdEPr2bmcc3QfZECkfbU/+zZLpAzICBQLCYri6LXAsctXif200
qrpbnsWT7aCV7Bv0WVskhtnlKqHOaRVXerVqh6OQ0MM1D2jzUAHdcjxnnvgojhrFk0yRYIsyrNXK
xdse9/WlSBOgISfUC4ySXQEd5Q+af459/tGhek35yUEowe2luheoCkJbo2hVO0AHxtPTZ7himCT2
37SMCZS1s4Ngt/c+gGTXcS5pdcvOY+JHDfmm1FV2geklfN37SzGEwFuj1KBylzasAiDEoGIhvMUZ
6RxzQK8BUa6617X6CIrmmaRcoEEpuS35KZHd5wPFYXmXCqrEMsWl+E7R/8B9XDc11COawP3q3ann
zTuNFJp+tBLMuI0IHD+5JybF8BPoyQwBu6W3ypYbOSczmaF/2FiHZMjKuhYPHQrs3i3jJR9F70vf
Zd0lhL5oCl7kdJbmHRd2yh3OpaQ8YMLZrfF+cz6yQgAY2t/tAuDw25Q2vPMxn96iTMsXn70ckVap
DPymNVKEQgHepIYC+v9otkcDhUEncWJQk6zBMSP5ZnyTwKxKPjFdGt+4ax9WnGmzbjtK6HWtvKjC
ABwbNaB0p5mG3P/QDNcjISKoVXI6bvgoTY0AoEUh0gxxNgRZGv0cYr0i/rSjcWA/Ea2TYmw0Ebt2
JYkMjeBq298qDe4U/ZJLQiHvK1f7WpNX83kcBDdC+NOzm0D3haayYqlnntdSdf5dff/XkKzfhTFk
8G06Oaq3O57kE6qPaTkjhCt4cBpCy31AhslyCQqVvIOjX4DCM439bm+NkouMhEW3v8wdgJlD0i9x
S/PyF653bK5efHQyXiNtqivd/n3PCT5JODn7/U+kj60Cdev4Au3WDiOFB3uYo1XHodt36t9P3IW0
tQF3D3l3RiReln4u6n+hiF/V0Hj3MmPPbNRf+vIJwKJO+ozmWPRUXOjlm7uTN/GC9N55u2QcJo1A
068EZli4/2tBtkPAdqQsFvSLvRBEmcMaKvH75Ct98/46Ce3tpmHtno1xtekO4BrV1iO0c9BKFTip
Q9R/V/rggcJDpWefNTnuVNGJo7LfEkh2UQrEOR7NlZyIQ0rHrRt4/BCThURmDyEr5l5lusTth78Z
7mkiNd9zgZ81QKLBEC8bGr2hCJnWybbdWVUNFinPW3i8FUL+Ef5xOFhFKFSxju0Y67wPqCYWEv5Q
/BhQ6wFm797LisAeHxmADEoLVhI47V70vSfhGqQMRCbAy5fC0DWxhVQ+9vXHK0qiCC/6lO6bPf4V
F4kBQmuXAGNVaDmZbgZR/7IolM1TXTFHqydkwWBixWzBp3PHDSFiT4ZNcrlfELSJaWOUD69cR0SS
97hLEemPKvN5nHuuHgxidP+wyVe70Cj1n0qwPwnGCFHL4FqUG9QPSGlmDriBiV7MYMh07yysQmQA
8Pd7LOHOt5eoRpf+oUb1NHINfI1ZY0TvSZQGx3QVcg==
`pragma protect end_protected
