`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 160960)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEMWgTUlbBWXai51H+tvf4Z4h+SSS8hRfJ6qRxbxb8nlGOUoz7ObsJj1F
+EPH5yrw6hHKgVn7DqFxAQQYHew/IdZENIhSg0BD41RnMtAxX70jvg4ySBPqZ0bqjcw0DmlPsYhZ
6tF+3T7a8DMPoOsghE1u/3ea7o/Prbtc9ole2fad/Pwv4W+qpbhtqJ4RKkxEdGx4Cv93BDJ0d3J9
ZglnR5BMLXIKH1s+vHXPD6Si9dtd89wPYgOt1OR69fyc8z8kAE7slar35kjD/6blwWu/t2Xsvz2O
B8Y4PCUhwjrCTlR6qQ2RvCGG9KzlEqZ9Vn5D23nYNGuNueoybHOkkDYh440Rsbxz9dmoOspuj3vn
a6IZs/SlkTcCtV20KhZXofYSgMeWvReY5+zB/Hsdl4qIJL3QFLQ5coEhMHw9hY2rI5QgWaLnbqNb
ke2rrrqB0yR4pZHv8fcY1isBc0chjBPEu1KPDeA4vREpLRbpJh4KFAufgMeELQKJaeuZYMD1zbh0
7ez0iwfhn/9dsEHSkgG/LN9NRhsTPch63j28GQVUk/KT7vJ1rgt1ek/XDEZwmMlqyL6jTOtGRz6q
Pcwx//LplFurkDxpKE+jvOlSsZ9xzbdztKRvPkfN+mDZ1kfqnE11GQQVQjVTp8lDgNMprS5POkhG
exA5Wxq7WEqQ9giXcCOPTeHr5rZuip99q3HPQaPWeZaEQcZZKlkCWSHBmczsFSwIJ3FbSaqLmjca
8+T+GDsdaRc9mij8zgd1ZgWXPlOJsSKjHDLQ7hjWZkFnjIm3RG8zYdjESAmo1vBnnL8jER7zVy2d
yql5eUICSPr0LHgK2H1jhDovTvQ9/V7G0JaLBG5H2EWPEXKs57G6XjsRQUWrwHShyI6QvW97HZW/
E7dp56ugoKnSr84bNSFY06tf0BEE1pBrcv+JSSJx7zcXK+j9ppRC79rjxi/0boZNQrQI0s0+X8Aw
+fso5x7lL2wrrrOyfXQ2yrr6vKm5Ze9i7rNJEQu1j8BoVjhYcWe26STFa1K+hXaDqC3lB5eH9JUV
9NvAzRykauL9IYu6W/xy296V+qHBQObgpBTJ+kuROGdeSm4PvOhO2TEYoROa8Bjc/++m6z9UKEUO
umaoDHk/XIAthSRucLEREaLCnEFE/eQFleb+5I4+rna1/aETCIwqF1igyPDI71QsuhOLD7o4QSB9
3YnFZZtPzVJ6mF1BORU1pouFrXWACg5y5ZXXoDfLuHU+sreu4XB0XLzeksxWSqPvZo/88/l5BuZn
tGkPxrnsoAi7epVjHophLe/rUASfhZajBC/XhpIdC/mq0OZpQASvCxxfvooKL+gIiZ6HcGAgfqSk
AUknEva/oKdWpXXgpQ7M1VWx5zeNU3qukYB1BfO1U4J8We/+PfcTkzR4JEb4n75lpuECDWH+Zkk+
JZ0SfkTwxmFtGnntMwnV2LSP3IvAzNjC4XBp9IzCDJAakjcKOYTWwiLsYs8nxCvBCMArbgwiE2rn
lw2zrY9ahqZbVsM9eb5ezMAIhRtJbCxhCpZtKeichAVArSIRzvj6StFEbNq0EF43alJQYtI8wGXx
XlnxLDHgj6gJsAgLVZWyyQG+8IElg2jhYthGfmyxeDvqNmVM0eEwFfyetnaHW5Z5Mxd3t3R7reZ0
TjzPq8m7FZRdJJAlg1sniwmclNJFbmQYGqsKqZa/M144Yw+MaOki8rhthyA+bTUFeg53C9RAAEoX
uT8o7nb57I7Wo8Y1xcfpMleo73L0bODmNvkt1dYLi4ZwLJb33Kh43VcPM/+ABbR6uzlE2nYwIAmD
FvT1W9sWUoa5Bv+8BNuArd6+6oeyPMGu+d5gb/HLqNZHwC+fwU9KdEe5auD4gARJPGHXi8/+cj5z
xjz67ifTrI5D5WNuB3f5j0w4kcdNMZetX+R2SC15MWEi2Ax1iw4VSSwhrPplLO3uJMoUKYlbDPdV
3pf1vCn1+fliGWrzMYwpZ0ThLvWAt30Gcv68dyO7MCUSWH8h4HbTWucSCh80c7G0LvNf/rfw0UHL
nvfttMEO9joB20hidQEk2hQHJ2WDhoDpPIdDP258qWf2EMEzTZKWOikqeMHjayIc5SKpudt+WW6c
w+mR202X8/fp6CK1PWnYzE26UYG/k8ii34Fs4JY474HdjJRk9zeEGl8BBvmegy/FZkLd3PYvHEeV
cziLJ4F0OnjmFdZBPn6svnjsWGPa8+nRB6vzj33faMPRHz9QSTBouRdn+/tMClZ1MO8L7XX+F84U
JRjQmVvOI704ziF9IB2Bc7blyIiC+hH816GsVtrvmQdfvujATemHkLnRiEo4EF4AM5qFtBsJBg3r
hwZNUFEkacBnDRBFYjuVw8D/bTlWRyb8dD7ubeo10gNpmvHAjYoDBy95q5AVmwcFzyGqmwopI3Qt
SOSb2wGdaTDVCZRv7jnvZnkXUwOjtOkiRBqxDDmeXtAlJAbHqwWvKceO4lsPfyOx4dTBf4ou18xp
MJxFjLssoJeCUI5xO+o7/Xg/fJbWizD9qo0y5XfarS70LhHfoRBmBceAZLPcPs4ILCVo8W0oxCS/
pkfOaRLVSpX4NrU78rM5ofmm/8bReAvHA1GUHxyOLJYb7Q0VG8d4n9pPLHO+ZSfrOOkAVMaiAWsz
7SYCIYRfG7vpDvafHSAc5Otcs/lupYm5J80ErYeWjpTbEDwW6WaUJa4GGItwskWl2/FoNlVT2f9O
YQ4tmSPDWrXJPJEyEE0mAjUCvbD9VwKSJf8PDqwXGU6+kKrM56wu09UHJR4VE++ZfCLGOUzUNk3Q
6mcukkQ2KExISlinqnggN6g8nKZXXI7SvDI5Lh/pQ6Apckimcu9pJXtqSJxyXiXi3anapMklN3R3
bNfvz2VQYhTw59KGL2+/FiwkpaASEmH6Axs3R8EJVsogU4z38sDAkiRIRcsWrqqI8rEfwQoziWxr
Af0haiJYmXof8AUSvlQPXpy3NFi3XY+vD4Sn9JQ6NhT0t3faP3s5OkU8sEaYwbnfzNrTdn74lymJ
YHAxa4B4wxMxcm4etwuizmJbnfWh+ZaRjBfbSlKp4RtFLuylXXWYCwh3vk9humILks32/dJLC1Lh
pV3/yeoU5JbQk2oO8jlsx91WvI0HurM1BDKiS8JkJnLBGtJXg/noj/Ox8i1KptZHr0qAZRqtLDFl
br1oRRcWyqhZNJjsvFeGr1RWqRundykoKLqAIMBK6OeMT9wsUSCr+zmC+nGeS8HlC+bIb8PJABrY
j6c6ijsfAiH/VSVlwHgGESxVgKeT1fPI0P91L8UaVfSraQWMNXNFARfDE9M7LK3Hq9kkaLyidNpo
cppEoalMBKc7JD32QGDFJD1ZvbuLamGPye+iuok4XgdzB6TEPWvcF/fb+WJoAPoWozbdsLZHAxcf
U3xPMpTFDu9I1kGjHvTrVrQgPRQw0mPiNWvYiFfLMMnxJ9ozVpsh8/cM886U2qnoveI6yg3R9lTz
8/qhhr8GZHV0s//1iTibaipQJjY9jcKcesCWdxI9BzxdbgqPpZOiTjJRgUmOQZl0N17EmXGSbMFf
kZV41nEpsj2I1he0KcBt1jvK+0GZL/tRTodmAb7NqH+E5pa8OloWwyL1FiWhuQSJ8JrFQ0A6BFHj
ZAouVhHse4tBXJc5Lq1kBMEbvSzhLglLJALWuexAtCA5ewt6HqY7tarzoQJJgQUdcBfChXYXawtY
jLddA+gMqKtoCIhfM1l0DOEvF+MWMahc+njxR2X7ILvQc2vukZplg5w5i8PySgGqWK4gvWdlUFb+
sB+5YatwA0nZItlwYjTBslf6ZkMsAwWudQZaPvn1KNiOcJC1Q9mmNA71RIB6MUUTO3zbWHZanb0g
sRsdtyZGdmcHEuVxg5EQP6S26fGyb+f1dFJ/M5kRPT2zFPTZgU/ySAy3iIvj9FZhWiLUuM7sd+mR
tvQ1Q0HOoC0C7Bm6/Jb+WjqfRVZQpJRSP1rsb41brExRf5R+PCR+BmMpNELU5bw0S7jfxFRLs2Wn
7BAZTO7hupv5XkT1R8PotGxzvoPdzq3hQQFdLiyklgMpGVcwkeGwJssD7AEmWeZiPmlCWBKgrqx2
M4u/4CLy0rVe1aWYY8qQXXrJwevwDQ0LTcdN8v6BV/R1Y4f7Vac/WO9w9iaWh7P6uCYh94aMt1b/
qZUpEVl+RT/kTCmrgelhkCXlHz6u01QGzkUYSkv3G2GNxvE3qlALA2UDj63r/g7BrkHTm2YKbQKN
oeiyKpRhev+Ukn760pPm8FPNkaAzqLjJkya8OxITOpXZbJyGkq5o+UZ9BaeRNDSA0R0it6LBSGz1
BY1izWGgAEfrcBgJnj4JAYheEtYtW1pLpvvMykH5hmXefpV77PlomZ0a8J/hbEzonKWJ+9lDKFf2
D8sqyV7M6AcRv9UStsJO9v+0X3S//wZaD6891Tmxs5XgHtbmaRgjcWZfwSUhOamyB4KApILFeBd9
8+s7adaIfmiTW3CqW4I4TjlnHTpT8gG7PwZqkIAvxkJgVEufGQAUJ2w1ny0ozmv4Xl2eMBjR/pxT
V9GqKsKdfmb5srF7Uld5zAUrq8e9hQeomr3LB1nHjS5faI3mgAQzSLp5ASkTepmGhNugQQjEuevb
tgR3UxSNWECnLkpsPk7kMMw+4AfnspQKoMw1PoLNFv03UmNab1x4UV/aU89RKGtclRGIOlb2TX+q
9Hch9dgjGDW179dNB6KpQUm4LpV176A+6PlwRknKjs7Bocl2rw5MIiqKLXSQLmMT6Vs3x2u6z7ZG
Vj2qR1MgL+cKbpjGofcI3MZ+T+tABVAZ7uSgb4OTljTd5+9SgKH7qPAek2O8t0R7cA93sdlTq9iD
Z9Z0/4IkJQvM0/0ukCn10Yf7l8h9StiysOz7FCyNV765bJBPpHKReSxId/NN2zdbk5rx7NQR77q3
wo89Kmpgh0VxEXZPtoW0Lnj1GctQ5IjZAzpZKz+ujgouK5xI+UBYUEmzdJlNfUIBCVwjxUVcAIel
q/OzVND1MS8PzWyurroceU5NBK2hGWYSbRx0idssvMiW0GZMl58SpeQoCGCQKvg/TYBp/77SkXtd
UOv/UuyqdAYPZPoJinFfBQbkE0kbLjIYnDVHDZerOK4C4MwXDyJsSHlcZzo5MboY3h9p2ABJNZZL
hZWltxhP08UFtQo4GePPn4N2DywF2/I1aY4nJV7OQ94u9dLmvlg+ocRTU3YpowbqQTcQFYjfBwhI
k4yDYUO98SQ3ToTu/6XRDooKoUgLUOoggVN81fyn4G76AhD8Q4Tt0a3zHt+HBrUVpzP2ZU8mrIug
5J2fBTniJFmePTfJIseUo419+ZR3BaAzejaE1IwCYp7952LfiX9mtM9E4Rz7NX+JpZC2AQ5U1GfX
RXpREhPR2xrJTD/yngj0hUm5dGGdQNm3S/yv4IHQs/vubuPYfp1unoMUNrAPTbumcsN/Hw+e014G
zPiqcR0mfgSKv77q/XRiRIxJ9o9Z3VuE2XDFagEq39XDI12W5ZgjXE+BDAssRG/oXgGnPC7z66O3
igLlCohQkBdyg2+ZjpCK0RNtJfYYkOFWvgnuP0uZNICBxv6kv2uPE1NcTNpimh7BFKEtp25W1X+C
EsZYtUC3iI4WPF93w0Ah5uqY6CB5YpE/r2l2oPfp5c1s2GeRHC/U2gW8FwWdQmMAfdqw2yuoEG0R
HX0Py4Upjw5cNjIVbftn76r46dd2HGjKfAvWFk7NSgqzrkpHLiS2HmlJI1JnvMKZrUNK1cdwNdlu
lOpK6bcE3SK82zB9RKNCbUTdToxIFZ3T2JcTuIWFoOIZYMSXA9PSwUq3YuGhlMGCa7neX2a1UAlQ
d92JfCIOkHuHArCUmddWRhzULwyzFCDZXk6ocPkLxwuWZaAcnqEfpZRiRwhCV+MVpr9L5WWPmqoB
pWph5qZYaUCIFwZKkUxxQXwWlbzsHJR9FY6vMqBgIaEEa9HW8JD650QGuDXid5cFXTf4X2H2rAZD
uktuokwbiMXgQ1OisCfIS4oM/sLebPxZAKY3IADUwP4qqLqBIHLSlJOwGfzXkVKx8E+lqoLde/5P
a6W/Ku2npdWO3KCDxpW1NRKH66yooaVf2pfsyvSalbcNOC2QZ2eSFYhgv4iaLCDQ05pPPdrIZ+xD
H0piWrzGqypgCrmx5Qplus8KBsh9jrskvZ1xTbyQzqDjdXJLOeaRdsUSD3mFwjFUC36Lg0s9qdPS
HFm8rSibPLbJhbpcs8EgDlO2QYlnTdgPFUm4f+2pf5uzd2E5K0EaT/ZkifwM7D1Wj0QtqrgXuIKC
O4MOpQP5YqXBHEu2QlFRObQD3NlxrrlchrQXPmOO09TMJiN6UD7MyDcHWtEcVC7rDQmLnMRBZL28
Zbsk7NQt9nOW/Zb2cQgrIl0rvT+zBHinYD84Jubv907ZuedRpJ9ZFDUg6O9UX8+n3Ev/j6YfPs24
9+L10fw5w8sBs9+sA1Z0y0snroq/zm7oObb59VLor0Lnus4MqMemulyZOWvl9IhO82Ev8PIC4Spy
FCO7eCZn4MYDm5FZnfmvxZcsZcwlP3hG5FXKuC2fbhHwJuYaH3RtN0LROfBIgbomCJXFmxYkTSxw
9GEwnJKuBoucC+qa6SDmvBRRUgAlJIpxtico36GRQBcb7yQ97mXr7USJ0eWPBDbMB84HwmxqzoL8
2sxySLopp1GBVLSlFVg9SXxDboGu6FO+JBYN+JCWwu5qtOoVB2SbYOfmaT0XVaqgVqhX6jtq0Jt5
ZkO49h0HkpTyXRFf2YnlwgZYNv/7ZhuoB1XYh7xPTPV0gcKJMK/6t+hflt3BKAhBY9lN5JNWY1ce
GOnfxJvZ2d/UI+0FMGE7P0OS5oyVQV4fmnMYoq/+30CqjrxRzv+EhhEJVgMreJAqCpBgOlG2V3w6
mwXUf7vSufFiqJVyW/47yrWveZMUSNhJ6PbnOJZeiG0zkuQ5uH+wpOh2M59tPkXklUnWOzRJ1+WN
uuZxeTy3zMQP4jw70WLSIbPV5CbJNDyBoqioqa7r34EGdNI2cGhFBIIexU6oVLXd4azNt5D1jJwY
Mm09mu88QFeG/EU9KyyHCpuHBJZ0lqphhSyZjeNMr3RcrVPw2e6/oHB6obKP2Lk371P2nd4G4wrF
PHC3QugrcOCeyDwrccILp4nPDgdnBxszbvQ2T98pj1LoezIBwUEEqMRTorsSUoNKybMbhEkjpykG
xhWnlLm+vtS6CUEmkzNeN5wd+Wy37kZvhB021i8kkDPA6vq5L+NigfEwIwCUZ+nUFW9ukd9N5Zpm
0JOckOeHLh4UMaILmiqgb1hKrjt3rwjpo/N7BbjSZqDGJGH4Wd7dZdJ1DYkdGe45nEiytAkYAWgM
gpawWye1f2jMTCekS5pDOIOgqCcc0BLST5/fDssFnQf4ELn0GtZWdqLZH5CdsTQf3Y7LV0Ed+mEK
594x8oHLZH7G/Pnw4ZjZbEjeNjanY77ICSIxrTern/9bb+dpfreF6ml0ZjOw0a19tqwacFYtOsi8
NQmMu0tIoafMBX5sffAJOofXuBSW4LwoAxvL9mgOmuhzvBKxvcdX2Vdc77K8tRY7p89xV3G0vXhK
ncCxIuxq2f9ipS0sVRHJ1rNqxT1TD7Lj96OmegUmcOQXNNB+cYHJ4Fv4inMref339+JVqvtRZJOg
WYJvRjSFnmSy7PCl6EzDFXsAhIFSIsOWttLbFyyOBpnkbctkYBV8nsoT1lHR3MP4AoFkBZUxDBV+
feWmhhGo5jTqT7R89ljZnocYhRxs2kkAAhXINTQtnbk5QW++lqtamIS0Tt7h0pm+OnIyU2VTxmf7
Tjr9rKL601hE5R0sQzCZ61q1b7LGj3oOQYjTK8iE1GL52pLq+2m3RjZE7xU2/VwBjUhAi99MG6p+
2kdOUxWyoQWpImun9KjHCHP+QjohddCmU1asXDZO73kEKQV40yLAi0/dGcKtYR5uLXEdQhq2A8fg
UcZdGINTyhFp4muCjYFiMz8UUqYLjNZpG+ICR8+/wwM9yxlCgly9pG8HQJj57clt/pR/kdiYEJir
dYuahaK1O+OTJ+/DnbEYzUS3oaqNheyne7zq1o9KJgyv7BqWw6t9RCH3soO5nkLBK1IYS+5YwXWD
24Gk1NYgNGb+jo14RgCUjbr/kTZFBUXQo9osbFP3bAYx8+Q69Omd4dEUcEZJd0l+KkyWJHB93/qD
JF3/8UkIgKtk0ZT1HSBQGLMu0d+jk605rwiga1uaEuqOO8g77FAXmKAarZbIibk2wr9POcbNOVXJ
82RVqjYcCM6PeANf6ibfAhEQd5E9ssacldkWjJevC82QHDONxDtMVIObqy0PTA48uoEAjJvh+rdI
7Z22AduLjMaEjx1njczjgQ/QfmPuQQxx7QA211oTUgT1mRL6s2nlr88GApXVjeaha8JAY6ef5rPt
P4N2ojIIP+L2C+U6wv//5f8pGJ6B3rz5+Uyffeij3ylBSkCFhdhD/WR6Ylab4HLvjjlQtU8db9L1
KzZJ5XKdk9ISr34L3sHL3jlRKvQm0T79WQT+tWLbLU9c4u0fnjTTWQO5KSJ+OyDofYpsBF4DpBRO
Aq03CPZjOESRiUQLg14Jy8YaXbNkKwQOh/3JJ7qZ3/t1kXh1Pj1hDeo2kReYO16Nama7dmvFxrVf
vI5LRzj15cXzeh6uqkQ/jRoFGDrmmqClkABqNWCFgIZuofcjUIJm9puWqtPU1kG2SEdkwhTPi2KX
AFnyTtFbVcB4I6W/bM4VXvfV+6Fb2DDGjJtCSN5X5NE2LDdDIpBerAJz3eeyYv1K1A/mPmN9kHzY
T4eSj4++ftRMjKRRLRD/Mi0YMqloQcHLRGIakGk82dPnHMw9I99OWQ4Fuwj2iCcTrqj960z3ysmq
eP35aw89Qo1OBNIBNK65Q+lIEz5qP14Vq9ejNB3+F+YbHBOoeKgxHh1cCkqIS1e2FqNLSXQvLYaB
vuGi7RAjBzpm+bNyNW2gTxyCb2bZHNtN4cPQZo2s7MRoTNEwNNS7WcwzKgDdjcv7zSCfOHEXvhe3
ezdWenTCI6oxs7R0ek3Vzy3QUxrLVTiJAzOQMNjXJDjr0auuBDa3Ccigs+RbwDo7GNuUkzWbjHok
yaTzbZ7yQ8t9ffqGqCJUbJmdWVXrDW25PAvncSeX+upKS87QON7feknlKWkRHXEhDdCOctv5Bq8t
omsbWrZRSYnFIv5hcAGczdi9vwfbDnhcT1X0jDd5cFr2TQDZvblRutEUVEwb+H3blqEscxI2R7nj
OIeGDNMHAhYdLB+4NPCLjqxkYyX9wcZ3q3wzI1IiP8eXjnsVIRbZG8u3X/eNa+R/OQKnFnOQeImw
QdqlhLtMjUvccVcoXtzmD7cjuWwmqikt37ILnElWGoc6/rlkExaUkm8OBQFDQpIpq1ZsiG+UABoA
0oP62yN/WGsNEOQo3C3MPxIu5y/9K0PhH7sxYsHGx/ZswaEpr/ZPDH0u7z/U/MgE3lh7+3u2JOB5
236xhowixRVHqEdZ1kkaE6/cHbhWbFvTZgasTQjfbpP/BwG7kGqqm9+kqV8t0PL5nKaH4WUusZj7
SWzPIeApqGtcceZp3rV85WyY8iNj/47VAzHpWxSY7+PYPxERuGIvxKJLW9ouQJ2tx8qjPrvsdueS
hyIULktgd8lNRYWIyYBhRf6uz/MiBUfA7Xq6PNjGzc2UCh/qWXNNYw22C/I3WCziX/A649rnPqzz
3lQQLd6ZtYxkmS8B2g8KZQU+iufWbmjFppAfXSuGCc791PmOZ3aDgdm6mJLQH8OqAS62PEjxlQdl
hYkwCmeTwW4TX+9BP0MUK9483soybIH/NW4RP7XZ+2Cgf9iZmxA8ajAx29/nvDj8yVFSGABtQGd2
sYAkD8SiUJUsXMN3wvxGpZ3bCTNz78dP7qLfiFU+XU3CqLvSAUBApZ0U+4HEFZ+r5E2wHxkOXtS7
CnNLbonL+lsXwCYMg3teivPLywzDmeJQId0RES7lg8xn5aeoT2w26lCC5GaG462k9KrLNovuPzpG
99SQW7V6X3SxDAA5jox9wBkssRhsDWX5mkagrGLOz515fxQItOM0kq4Aqp/ipvlzGg0gPe1q7/oQ
vHU95xiXvZk/RG8wxnlEVTwrNZIfUnNGdpc7aDZHzn86jPW3cfrLF0uxZQFW5sqFYCcYaOHcvp7M
vvruZTHYbX6AVceihy4OTiRmv7cr8B16n1UtFtMpOXeFh5cMchkxCIJZWbZgXQdW1/+Xd65T7dzp
Ue4wHtzMHKgxKY0LJ6oxaQUhZ5Tu2n8PXSLmwQugJZ35b8typo+SO8cf77XnxkIzXdaBEcBFLSqj
JGNKwIClHjHMaSs+icxsYhzPxNY61z5VO/SlYI2WeOnNEDe9VP6PUlkTZAc8t1BTzMvA9dxiiVXZ
J38ccBN8DUELQngaKkdh2v2Oj1LZBSr92K+e2R5dwrt7wgChH1e6j2r8R3LsmhJ/QqCU2/RBidkz
3FhTbXSj+Fg8D8RXa2lvwssUiMgrSOUGGqSNvmotQw8zMpr6hCx5qdGgmeXBrny6SsOj5NgGduYR
gqTP0fb9Ovr/x7BD7ZNNCk18YN3vZZ3o9QU0Ek/UwohKEpTay0afIhFB6xZRJx6NaMetz3kMj/4J
HMv3Y9YOuyE8OHBQJlqR2nfXHsBWFkAEG/rCFD2voDZ8U0ks/7iNKS55oHC7AmS4nhYhVYXOiSsp
16ADCt3kpP3b9DJpcPHTuYqtQqpYGyZHY0QbPYZ9gELyV19EniqWmQ8+2vJGBFoaVzBwr3UpeNRQ
N4+6qnTgRoom517Z/4zok+TawhIOAXN0UH0S4pGk/C4P9VybXY3tg8eBsoXMVHBiAqJirN3YjWxB
rAiJTt4EEBejg55mTarqmjisY7Rf4P8Dn2SMkSjdUofI9FzKNLLBT5ZMeEEtg2JU5OYdNfeYbjYz
fgk62TsBhq759HF/mUQPQ8pIQ2ZjassyGgBmyxNHWUwphe9kN/eB42r31vAs0QhBo/YfjEnNdpC3
gJ7uGMNSRGPyZolwo2nKA/8xEGvFxJ1KRBUiO9VE4cJwwdSd2aq4nUd5RuMQ4YxhlPtIJR60gneQ
SpdRrsHQqSzYyOK+kxa1nuKa2ZxEEvev2qrYF7BMh5283RC5zQawCos60Ho+rUIC8hA2WZJwJPT0
Eps5sl7H2kdK9q4WfVcZstCFZ0bv6nOhW/Yz4Byr2PaeNKTF+0G8+unmkP4gSXJWf9n6WuhNiqw/
UYCBqaXyP19YPcM9LEKiMeurzDj/RnbhjNkKttyfdQ84DdWUHYVmQMA6hLx88n6jsnrHvnvfbxEC
kQaKehkc1ahr72p7b4FG8so5wy47+OvLuxp9wUbXc8LCXRH12s3YBpBQfcy7oIJpC88IDBGHMUx/
oAF/BwDmXA5gsLINyyzJrhfu4Ci6aaNiYXtvvn5l+xA++UYNzHVApUuMgarin6sGAATV+Q369Xw+
RS1WaFt1Z3cdtdjUBRSy6fwGbP52YrOsvo/OwUvfWVuzz/73NXEBnyCSrFx1gJKLtFj/E/MiXdxw
ohX0+R/xrh89nQkbe5xIIA3UWntHXjUpc4RBa0SBdDAyr1CGANPhvlkyGpkLYecpi6mXy3RBxj/a
gWm3fPclNE4ZUfQRWiw/V6xXvzq04P48bbQ1ObDz5ROxjjm4Y8qZ3knABBdkzVak5uVZPO0E/vUU
6TCcT71+p+NxFEjgk1Yhs780HRbeMtAW/UZfYTTi299Ap5HzeaJxsQoWCxXoH/t9maJlv5HpkdF1
3fl+Bwjt2Ybn29qDK0r1fMqs3LYi3ID4kxefHudzdveL8Ef0yxez4PTvmEjegZpPLI6NH3WYUpVn
N8U14Tdq9VT4T2Lk7koAPmd9gYov0QU8CWZHE18OF+W7LEps8k7iSQg189bTZ7vrH/S2TglxCb/k
9Z/k7bUL540zd3X75Uchj7jQwiGSGZOMaQC+Ki7DnOtBfPjwuCNX5saTZuVzohb5fKQO4KvFHS8O
r7q8dB61MnrOqryb2l5LjLOK4KRBmaLvXOaxTeC5FV/iouemK1Jx5YjLW6Cz1U8TExWooiOJ+0Y6
nq6zThMfMiC22XW+UT8RRxjOrj+BK+LHgFRC8pb3txzyDOMzo4qHc5yU1oWu74zLqUB+0zU1EtN5
mHrDUrhS3aDJPS6hAM5pnk59yGRltPWnTUM7n4dNqCSQmYMqtFzZ3VJ4GSv7GP8yD/T9X7qSpsQA
SgxSc1b0OtZquOLzKCLT/cYdsFtrnN8iRI9j/JshsBApS6tKy3gs9m+Uq/5PLFkusOAbURhZctHL
h/KtZjfF8lIaxU11AlQIgzXlzYs/4Ek+aPVuYdWUwCUEuz2pB5rgFW0KfD3KiYSwN4HrF+tke22I
Rj8mji7mrl7oPUjiZoxs5Eg9zc0HuxC6/n53oEDPxgyJnvA7g3TTc0t9WKQ/+w5ZAcxWNbV4D3ch
auRMrZOD8U/poCZ+gbmz70N3UzThm6cz1YC6i3UJC2GqRwm5Fdz2oB8cKNYy+BE9x3/5snJ7DSVR
2quOuNLojv05uwFgGVf0piDPfE+tjKJEMVA4n1ACw//aWlw0ERf5cu7jS+LNQpl3OfbBkVHxh9hA
+D8s6i7UAb6mzX883G2PJ6OH9PdtCsqxieiiqbF5VsxZx9eqvQEDsOG8f4fOfmv0+vafJ0W0NmQg
xAouLDCl0vhb6C+IsW+97s4JWEYNOmKQhiobDASHRTsKrb1yzl/NxGtGRD+4jJd19Wo+ZKLkD2mR
IyizOV1GPT3YI13SViozxPwyw/ltPDX5J/5OTHclwAYTspekOXK8sJO29IW0yKAvb4mfhIpcRp2j
/Ye/9FZpw0WLx114E2TqiBzTJtVYCIkST/TQWMNgUzBbvF88KErhfKLVBSvDGBg2axHNTLpN/DTQ
/b4nonhABPWfmsUpRhy9cjQIuNqpHaKx3EvB0lP8RK73Ib1iy7uHaPOYufJ7xCIGQZK5d4yEIkJ6
Zq3dxxxAUIRPowgHv4g4sDOZ/FnQ0CTl0z60mWtiTz7r90D0YbvZ/ovurDPHxTBcuwgebs23cawN
ViksCnMmr5N0/siD1iZJUo5tJ4+FXPBb0tUfTboO4AWyRTnzVQfFYpQLHQfTpnR6zjcROfb+ZCPs
R0wES08sM04OGKMPaKi8h5mrioaPW0VcQ9xzZA/NHwxFIe1H+rwQq4hu0rY+1W/VBki6CxoCwt2R
+Ilthdez1JkQh8vBwzqyurF5MZ/v/Q2wk9913yLEKY4UcPvbkgjpNun3udl2tYMt1eTMJa3f2sKN
idnQA6zi5pNPDDm1ukKcru7sfHa7kATlVqd1D5BKIu1Z5DtJ92NvSKWI+2tbQST8G6u4dFjKnidy
KTpHVbr8FucT77TltnUIV1bLZFD8aQmzKiee3PH/XQ9JP+o5t1YHzyEFWbfsYqXoWfyUUr+F1dLG
yUc5gMnEd5xwVwzdQcGvaKjrCeE92psYk6LtDxIiod9t8JyeaT2pTe+0c7GIL3XxHpIlAyiTfEUC
Gucb/PzjXp8FS6ohTNkAYUBsBqoeFeg35d/DVzx98KPl2mI22ZhwgW55rJrQwrqTnPqHiDv/NAVt
cG4f7kQw69a9Ex+nbh1ABWz6SxAPwUj6jZyRqhR49dIUUWoEMM8j8hYvk+9Om6+Qx+lCLG0hcOzS
+QQ2vdJQFg7WzGnIiEYTiFdAzcH5q3SECVKOaCQz6LNyfgIwjEv91toMEIWM5whftrFB/JAxuJTC
SKJ7PQagcj6crZsB4aVXNzDwin4Ve3/fPW6193fVbw83R024D+lEQxRf51eD8d2nJKlte/T1+xP7
JxI10uzSgS7RHGygjxafybkjE0LtlE6OkGbYB/mEXhWodbFwvdwg13b4idp0dVtuyOSCLxbGA+Ej
UkZU30ffjlxtztJou9oojHTPHigCMsaJe9oxPXW3MJeUBrlhvkXJD3+cKuASoILoknhZfWdT3jRS
kz2YWlcwfRfEmL9pScr0SCA4vRANAt+KNPVLI04Xzd16O7C82x1mcRoMz358M1LFNmNgWq235Apm
4g21liT8CD7060Ca2C94DjGADT8LAYasC3BHh0LzKVbwzhne5yOVZNi5UpQildCqIRpq8IxmQ1VZ
FKjHsbXl+XHlzqhDM4ElqdcVaBzk74ERz5kaObmb58U2osqOnprrJ7TCWMMBwAayZriRjxZuY/gz
njOP7QHXEYT579MtXna/+Bs2I2gKWL7YCkmIfQY/oa9nLbwNWj48w8qtUVrduGx6c3yWsocPj8DY
aU+8BOqT9FTePYeT6Wrv47ewHS+mHUydombD+NPVZt5SPzuFTJsUyCCoNuBt5594LrDfpi7W7cz2
Aih1Amfum0M93hYOXFXhdUnNQiHclun0rpBkAA3NAxg+jSO63Bk7GHqPon3ao+oEqgCLu+uyRrdo
REim1TLTZzpVqbaiudUCCrqfLJb+kMpuG6GPqlpIyFWy4lVJoxtJVNReoh6pbXk/Uq+Ng2zLFdSi
B8QS412KoMIj3bRjOs+OSlUNZcDFggpzJW6S43IqTWHmLNl2Y+KeQfAISyUdnemP3y+1HbPJ9MIS
bPqYyCln74gnUTki19+niRnHcHA8hH6Rlficqa8KwYjp5hiQPbJBwFp4rzOzuWYo7KG3PJ11S8Mb
Nj9eiDXs44kS9kJDIsdMhvqHGvkQRKTqLq1MrnvY9rhgQ7+ptXGPHFmtYPj46hdlvfwFn8U6R/sa
GkRwq5TmSt26Sy6WG+gymaSOb1+DbKEGTxcXHVPd1KkNj/Yg1up8IX+jRwWcRZdtNngxtHu/e3ZX
5Uk3gTiWH9e4Aqv6YRy4bQfQBXL6qHJQNwJwFlzZMsAggQCzuz62B5AcdK/X7rZBse1mxDWkS18B
sXwMhg8AX4RF6x88Urs23uC/aY4eNYqJeSuy8sjRd4YOAkKoRZjcok/VgPUGLw0oIfEpQMq5e1DB
Bm2nHjkIAKWEaJpWeLHIwCUjwQhOpcFDz0Um+nyqgK8W/b5hMhVR5GF0T4mtyxmJQrKtqYIaEf5+
Pix3nb9jzO4HCi4ZI7OwAgCaCwxhdAzBE1H6NBXL4xTSi9a5JEo3YtzQ9sAA4KZazVEAP6dT791Z
zFhJzrVMv7HeEKwS+fS5w5MxLRepqoG3FAHYVKrNzgnOgJkYhqYQtTJmfxk0EZIolgW7BihV6deI
UJB36CAknN3qrkhbJWQ9cG83ABkKushkTSee+X12RO1qoxwtw7mHtkrl0aY+Kdvl/S4ZuIA/POXu
BVtQ+anVo5tlYS9s1SMSrF/4FnRuRaCJSUc6B9cI3MKsPuLzXse3ssHUqDOhWMED0HSNdh0ood1U
0Q0w6XRVYzLmvBcWQ00GONOSA0/6qsXSbMDNz/FrZWgavHZC9dBM3SkbPA48x42tWIcLHj6DACqD
i0V01mW6l6fG7wPZp6xJsGc+9NrIOp4xVw1/2lD5TCnzZwwOEeR7rzLV3uV+ni6pzO3e/NmIaKhG
h6uULwtPTfn2/hKR7giXN1uYAe+I8X6PD/G0hq/A2sGKu2G/c3ZUTOvBI6h1/87ECjPMoEM1YBSz
d9QKcD2C/H8dFqtE5uhrAG5a8KYBODbCuwYykf2JJMAC2Lg24SSbgi51RQSkPAYBmshoE+np0xjz
W46WfOrPz+nCzekZ8Efk+iX8GZeTMQ03BSDf2IldGP5RGLkOmIxo/dzv6HuI0M9cafKDCFjEIauB
D+CzhvE9VJc++0rES6mPrGsEbM4x05yw5QVSuUsy/5TFkPwcLXhgGw77iU5EyBoRjz4g4EAqT2s2
YEKzxoj71c/MCYTLXBVSU0T8xNmA5PEvafXVXFOZ5rWvy3X/rU1ct4RrLTVstvilBKI+AKbve7Md
1156J8abwpTWFuGi942gUMEEuWHo5yRX6rpcylEkwZp4oscnCGOO3cx4X348tHcMi1/7O4l0MNoI
+nojSdMhCJpKG1CqlXnz7NmF4GUaAVN4KPovW1FDmAyHmvjOzbEC6mupBsvXIRm1ktlVG+/QcxtQ
CjTLv2xn0IJ+oujiG65MwJYC/8TritP/04UoAMpT0qkTVFDaFZIIFMTQkciC0ulL5k5OaNrZGFx+
QfDQL+vDG/sdw9GdXBXPJ2FJSHA1BqhkNCe0a1u9w9Mp4EK3cl2eIYfOToFIGwV8Jz3TDRG6nOrY
Nokou3+S0hOKW3qD+GsXC2rbJwTHS7vcLS5VIaP9so+QkfCIbv7u15MQuJUQahh0NB06jOCVCCZE
4POdHI/Wq3iqeHEWMqWy8iW5dSZ2x8HnF1kRXkbebFmxN740WsPvUFgQxuDvNVBUV64JDygBrOjk
dlNyHaBDK5uYHKeX9Ws1H76vv6dwl3XVvRdxTVlSNmnQmdV0uQxldIf8yt2tumZNlvX2SBtmgSuc
unyqpihnOQ/yq/fnvxPPWYGjDFbu/V3IA/zaDRGrkr5NL7fQp0jk5UGeesB/snaE9Kh4YUp+GN7x
Cumz6CRGuzeuFWBanka5NdGPNVnvejkf+vgWgcYzH05ezAE7Gl/vyl71lVoYNZ84olQYYcJKzeoA
r9pw+GQD4sCpVdjDf/CouRT22STPu1qdKF9XNPEJujg/XCDDuGboHGSEp+2SGStolw56yc0cDoN9
/ZlOnJhjdRknHZYVTVLauBr+CWrE5uG3/J7kjzeuijKZYtyxoLkmsPntTJm8Aejl0cwLbR5SEZrW
AgOfXoRfoQh/uZTaWQsg65Qxc8vXfST4duWHhajS78LqfRVd+W14UfZRfUIx+4X5MVTFBD2P/JEN
VLv1RZJUObuPhapbNyZH6yUuoWZHBgZYgmLUXyFyVixQq81x95xD7p9mXOVjJSKzyk73uV3cmmta
M4c9ktdfsFfIIFrlQNBzZBMZl7FdLcOqAGqp0mil52HUB1mhZtTZ4nNPat+VHZk3pBmhOKQ+3a3l
2DJx2tAJxKKsWpJq4+jQInni5vWi9AfFXEy87zHjki+NodGNNMqoEtgJzSPpShLQiasty7u0VWGM
mnePDgOeQVu+I4odJdgVjLK8BdmK+8J/HmB1Hu5Dv0iRxOFQQvxqPVKcyij0XnJ9gfFj8o28XqPp
ySlYeW9aLB08flbZ+ahwj/WS8Q3JD8cnm5Sgurmfi9FNZ31F0oeH8AQwAx6dLCX7a2bfNepHo2oK
RQeOb+MkHHJ8ybDIvCv+pa15YW366i8GixGBVpZKSxQuY6Gz2rZzVsVyTIqK5IEoWT1TCLS1tENJ
zYNF093ObXVkqZMRSYrVAPSAGnx97De6AbPx2g5JdDPQ1d9Vl3tSeCMKe6YsbrMVbyGN8JWrXySM
4FlqDTE3xnXktE8VywYVcKMqkPapeui7apc5PFPcsBbgAqvu8LGF0lDL49kheE7FAm2Gds0SDsPx
kO+EbRShSih9twrkRovrpiM+pnW9OTMoMKZsoHTHDTdRwn8p+DdSNqHeWb/FUwUwfTf5019RgpRG
rj/SvmGbaI6TH2zeTJ2nMy/L557Y++/TBLqx9vFzYh9RZYwwTK90R+JPiXcuHJErPPzIH7EDfmJW
voavHC385jIhgp2rscrHzdTWeim9U2WRvwUt5BxrEG4DWAo3MubrUL8vKkv43bnHEvyS/6t4eIZs
VOAB/TCjECazwVIMGNe8SvpvXPsB+DiFzSOIopncfjEPNjiOrgOvMcExa1F8u0LG6LAgarnXSaxd
fYnRybWPZF4NzTft9D0bNlY8OvA6Sn92adkjaVarjJzXLrvU/fwCI3Ll1O8kQ9YKBlR7LWHoRCDk
IzKWhO1kL4cPXMD8dWG7mk0QtmOgHQlhN5LPHn6Lps1WLOjSO858GGbGOvzZ4FBssBk+lkn8LU6c
C4vrgt8xBHEpXB/ZhZhpEcphl4hAUFrixIxECsv1Kezz1bH5V6f7at1xd5tbjvsrgrUhw0BZ+MvK
qpD1sVa7VCkmik6ntdrpRtU9rwQK3n3FPecKdRzLDuuKTOZLEgnhlQnIfVcJeZAPQPfcWP9OPza2
ElZqYEQpy9ksk2wc/km9yLT/Kow2EY2v0tnZHRlLMoz765f2VB77SuMSjgDPIJs/Re73ldwDPK8c
MeBqkbFoNrIDeuqkVDEqncXr2bhNo5Ptk/QNlGZi4zaOZQlRRvHo2+4g2AjPX/sqPwgrHcOugqY+
9hoYFGbNSGlIL6Aj2ojizy6AyywY39E016M5vkh6HKSQ1GrtnHcnGRqxKU7MUvfra0mYP4j+YEll
2TNez4DbylO5XDy4e5oLPcoBWm7FARurvdVY4cYu4ywgh+Jyt1JmwwuGslrwjxeQiVMmT6bf0jJA
Nn51VTBc2pyWoyKZsYA1RhNiNxhry2gmWO37O5ZSEGnE4yRKCJm/2koD7j8EKecFkYAiR7jQ6Hak
x+u1Gkp0NU7Ba5ZwxGWM/+JhyehLCA71LfLHQqPSOh8KyXbS4BZswi2GvUiosIFegRY6BzCCFvK+
VFHOB8AfT7x4PSGp/2sb6GGeYIXkCkrWHiq5AZgR8IbEO1ozfmHCbYEl6Qtkj4phNAKWyRSFWkPt
Ng3wSFHBc/22XTBr8HvV2dZJdD/94KLBz8jiRHGimAcojii343n6msXlpfjf6lqFdHW85kzYguJf
jkn+8npBXaX0DZLIxXk4f/Cs0iXUjpKUfk+K/omJkIMQVQBBQw9HtSeS1mqq1yywPHIev9hJDf+c
VD4OxoX1g/pcG+ipREXavHZcemaqfTwN/HQKfUAmbeoRpgipo6nV97yBaZ68iigwixk4JY4KF2WL
AL0Ex1QiKdti0VsTpCkDNHJgDaQMcbDHpkw0wJzw8dPs5KMucg4HYgpasntQlcigo3h+ygkA/rdE
M4jswL44flzh+xL6z2g4cR79jvK1KBEQxhtRqTaeGuhBqI2H2o7rZEtMVt0+dGGGVi5f4NURfntg
iRpBmZRWq59LSaLSJHlq3OD3lpqwoYidQo4BGzRfXNFOIdn6SuXglkgps8s3pEh6lWhPJKyr0d1M
KS4nuqujOpELGsnIHRM+/rauutsxR7hHln0ptqMjqHJumXSIeaVVttkIRMVIK1h5q0M2Q1QM2w1e
TiMDNWceyixneZukxostaAe1dZki6iCgmDh6xHQTK/WNkNzaJxHBYRGHozASCoUZGG0tPbg1FBqy
p31WZvwp82pDupHj8QqCqdXibqnBh3m//woGIS1uVjIRvnpjQAZKbuOK9t3edqHxIFfRc5qMyy9D
EsxlpLU8BEKdM8a/kAjd/5AKm5KOuhHdB2qorkl+7EAp9BLyUHs8q19PWEZGXO2Q0aG1UiUW1H1s
zvZt4dDbTny03klMaH/Xfmyp/fdEOjuGc/8fPc06dx4nVflLthldxHhBJfQsl3zQcTgKkgwTJSk2
mvbrNeZBkHqNtMkYejX8gFL38fZuLcteChBFJRrzB6eQZP8YsBMbR3FoTVbnfBjTMpQfrB0OKuJo
Ky+KAag0t/tLvs3RAQ8wr/y3KOggeFcgA7DoejLR2F8oE5yNonvBrFzORtXy2MswkYDi/9G+n23L
okaY/Voy3hjArur28y5SjEJK4hrRKRvubUMfGjeJ6HTBGlcIQvBxPepGjGX+PQQ2f3Bm3dh1zXP4
dEYhlOcHJzBtjl2I3PyhDyIVBswUuJPPCxor71KIWTg6tBVfPPb8LWJcqTThYWZ/2I64Af1NDcxr
5I06rgV8cBIjDZyK2CYKWR+kq8UNZW3bw2mEaSwRzmFZyDKUXQndCBlduY6TneBv1o5Ds+eNcQrd
8W/mEJb5x+KbY4UjNUM+ilQsuObaUKNYepgCCGQbWM4kzwS1MMGjy/OslGGaDhzK4PpXWoFg8FRT
B47SWipzTvEi1WXUgws0Ebd9GFJ4WwyxhzmadTABwOYH/fmeca0ET7vWsEsgPBmZmmmOGgVlF+m8
l4jZYNjfgi/z3oT54iIZr3f6lTX0T3DFUCf3vdQZ2dwqPUXHf7kzmoCfFqHzfgxiCC3CY5WHfiNQ
GjmwhZ3PnD2fuzOL6bdFLQctWqHbiirAAZrAPioKX8ZvbfSCTFpGv8kjdC3tmKehVvh4kCQhmfHm
UWSVPUa+wiy1MumZOCcXg/axMc9TNNo7v0FxtwtK+QKDQIQQ/jyf3/AHvgU7Ol0AEnWdokDf79AJ
/v1IFbauqnA7G144IMojm58/yDtheVIMNc2XLbBknb9OVzuNnfaGyfJyEboEmOhoR27QXxY8F4m9
CjjddwfWeh9wmHnyxFzuAaUDbzzogwy6Q3cZWIchDWA05IynwfFRfWDzF+fAZcRYrkaUx30yw9Zc
8ky+/w+nySIhfGG6FSnkkHpfpNNfKSBUQugweKcO5mw9A/Pugw+JnKSA+vFjndGw7ErNNbgi8ZOH
EYSqTXM6zaEDabvTh7SZpZ33YtWR2s4T/+1+D1jIKUZjljnHmdjn/aqZdE/l8Vix3kkxrpVGV2HW
IAHuBpShxkAKpvxNZQBLfd9bYwFSWEcAGIeZuydSpc8+LI3t/8C/b5mlA1vo4h8Dx32b5k80dBDT
uSk/u0zfdxKmzFhSUm1zW6B0ii1sa4HpHfiMMhjp85PfbZUKib+j7Exb0a01QKBHqCplQbH6BiR+
RO79+HiBNqyyWkBKmF1xQ5Paw81Qyi/Bgs/JzqPKU/RedD8Sd4cg/91L5VIIY8NvOnDsDHPtGTO5
xlpi9tKES7FJybq8UnC6jPfr9fiw+Hp1ac5SSnirglmyx8D6j9mxJT2/8jFrF3TDYJszf8rv8tqX
6lDfwCZk10WdJWq80LBgNyAh78whG20enL2YlvaDc3nsQgkNg08KsLwyWBvS3pLJkQzExwTpbBZD
pUKUPc897/lOUnqY5j0vuJshsZ7WOBh7FYQhvRzenJzlg8ZZbiBchLnhRLmB+0Tkbwri+YyR2cQa
zuI2r3R06lkD2jpoBj0j2rrNfAunNNNDwqigqG2yT4yrYV7+MI0W4lGFI0Rm8363CRa+0i4OvMx7
Lqfybsi5og0+nlDA9nDJL+wfP1LyqMxkhMSXqUPd5jnMp2A2IFUuEuiBYE3v/QVqWZAmvkwPqet4
U3X884zlAoXJEWg2vXGjD5/xWkCEGE/X4KEqf64/Sphr5ylDfRSySWOTLPNaVoy/HxFLqrjQfOHi
aR4ukS7ZIkGzn88viOkWzJ8iFM6RGEMA7kPGOWo1NIhzmQ2MqJdzJDX2LtrTkar2hLrcdgD8pcit
OnKHPFYwbp14+mnhsW3i/kXuvu02pJJs4v2ciEWsgPwqan8hzfErJKEr/kMnpGnaqI/CjaZPV98M
R6hxrV3t0ABQ8JUeSIAdaYM6BN1PgOE1XCHWCazzCu14iWF92+um6ieSiMp3CqOI4ggc8YXOY42N
2J3rdB3LGJgHL8pvNFA0r4mpyPpQKyOutAApTeqnKsXlZupU9cAbyPJO+Tr7WYcsNwvnaHbJTrzZ
uFNKAgqk0h0DCs1heiHMANglSK7jE0GWA9bSBTslaTX1HsciKo/N964VJ++WSYuM5inecvNZq+Y8
SaR/J10QNUJhX6FzB2mPUQWzL2PGuGxn6/6MTI8cnBKZMZP/GjZMpyZwi1roNxC/nhf1OI2qQdZT
dDOPkF/fFPPySzgVAQByaaXT4tavTmt/XZhyJgiq1SOyMsG/hHnYSOJH8WeT6CpbEanU2Ulerk2d
2SdHpDQWDIyitGzKYHkV0spByakSW3Zl8yavFiPLiNSIC+wgQoejrZKbrOPay8scvf4RHE2ay/sq
dZRL/DlItRcdzK280Lc/5sI1goD5gEW70yg2jZac4Am+9pVT+yoB0qjWZsvsVKGz4hNJB4OB2xSM
ptNAhFc7w3T3fz5M59phKFHAA79sdtljE0pxjMpg6gnzoN6KcWndWuCRMS4PgH+7zw35Np2DrumG
7uvAUO9DN3gN4fG5NvxsNtIRaPAQc6hYUL1zfKuxM+8ZD/+F/AZ6UDZKzCmfsjaclH1mvk4xko/Q
QPDast/3DBqcErQTjpjTDKVz5Vjkv5Ku4wQdvB97RWrVnYNW/aNb19+fIC2tmYJAnIfquQsLX1eD
WZbn2J2EWnd7ar6Y+2M2AWWC2ef5Xuy8RNXh8Tn3I6MPZ19a3daeQ4bEeZvwf0M4ES+aHSsFv6mo
iv86caRZvzsJmD44wvDh+4HjRtISP8VK32jKd6v2zQdqXqUXadX+ND2Gzk7DQ7PdKSqjjRGx6Phi
5b8pqZzfG+qpEfTQul2niRM+uYMr6fjrSxIs9O5uIxrQOXgawRpdywGJjI60g3Dxcof6/IFk7sVU
OvG31gCoEBQkWswzNLEC9JTYB+gvLWFFo2+ockou5ET6wvWkYQhWwcPXDp7oOiLV8LVgVijPxU8T
GuS8GX/UdkNeLNbXJsBUdgBGCu/Z/GaQI8IFG6RrjoFV0sGnBdxBwhpFx6xhMIYat5SN+AvnQ/Hc
HcWqBDYxKJWAbevTUVj5QBnInXxCuGjAHh5031ApOH/jJdQg6pl3ubQA54zvVnKZD7SW6uvfIkj0
OUDVKBCw0PIh/D1HMwtJfMI8nitTO32t3zR4RkvFqkgMaG37rG4lqcpeqgAIhH/WWdS33L+jfBKM
VAlDTgKoGNjopDV7w1jYqsmPRx+OkPxrqXrt0rHoBU4A4ouBJVDhF40LVARA+f5kd3kf5Ays4X/q
X9h8rT9M2o9D5A2YymqVkzo6upc36eOOH574vjzUbqjrUO6juItJiglqpSLMpiOf3t2Ran6NiRdw
aFe1SKLpVOtXqobAwOwmcB1hHLjF2nuhmzsZSHmB+vreHUOB6hVQDho9n31JZqNWPIdRvVOa//5t
Yxlhyj+i1J8I4aFoEuLh35ZfBJ3EDC+cx8EGmnuAoIf4t1YZGRncEbyFepFnZqNqOWBkZSKnp4mP
ruDGCrsC84I78UGzRwZ1ktMyuPdtThAmJIQsRAjgKCbKtuKmzbTnIhLwzgHhFOJzyIPhAEvwI80M
agU3aHsNjnm75r/rDccocy+M8iYR5S2XUWVqe8K3nkkrD6HsYoYR6lAlHRNukVGulWx1itYylaiv
Hi8i3k/mc4RjOMRYUlkGOVuoSEqhU639vesJPN65Ghg4Y78epjzEwb6p5zWtDL9W4rryrtWinC5M
M+v64DAXAYe9lFJiQC0A4EvO7KjGuVfwKzcKc6vStT1S+nRwY/umvEmmV0jl8tHMiCZVGu7F67BO
arXFlDWRcEELzT95zKYYwK+U+LqloC4s6Rwn/j47oIi4PvCETx9L2GGwTZNFpovMsGeK6DjxE7cA
n63JsFRILSBHx7/G1qtLd+rSxUJ0ULifN2lMUMWsfhRKUR+V/rQ7JMhB/BSFjLBZxSxSLE6pqyE7
5xclSWxyr8Pm5yFvx0Z3HnZUMt+DfENeUv/aytP7rTnYsTp0u8U8V1KQWCCqqdOMKDPwmMNBtjc+
PkIQGQkeJm/zcCPKa2eqHwWLjpYixtacmyeTJW7sKk/6QX8u36vjRAaSkohR0cWShwRoI1fwUjKj
j7i1egu2kMn8xDSZnGnvSkwGA/in9RKIqPR47703s1CCJc9s+X1yiVbPlUfS5TU9551nMC+BvvQR
QhfLE4W8uVjIQ72nrUX6mlZs9EA8k8lzzxOpchLs8yqpsycoreZPQBjXDuWd6K976jQMga0W0ORb
CN3ZfGKuYPYpTUWVDwYfw87J9+RHwVquExfob6KG4PjgA6R5dyZGfYHgfgfYQnkrSPwirpCx7h7N
cPVGjPYEeTAQF/HzUIAW3YT/ysBbM/LjDS9GStVKVIE4PV7j0McOtyJ+Gn8zDiVvbo5HRVK5C1vA
D/iRgy6x4F0db0P5nD2Y4eOWQ2t2kxTR/aZ8bthRoOfTyVLaFU9ZsX1ed3VhQ14Gu3qCbxpBQU8j
yS0h9h+br73PKW743ZS8dvS7sieUeH/EbnHgGZEt2CK8+4Tyv58iDGnQOBb9zzJRjZ22g9Fu8hGf
t2NpXqrutroJXqXRhvifBpG76MoKfVMl3wHEnNJ5ag4wshk1+bR+kbZNC9NG/Nt5jTuinZNdgMVa
G8Ho2BWEAWsFV2dqmd6HJcJKVRFv19a9ovSQ1bO9GroMJMjlPzCaIGRlXS7KKZcfzEC0BYReJWnt
RQ2PhLcBZWbi3DNMTrzVJO5AeK0BCSKPJg5E+fcyBTrn4EwdZ+zl5eL3QJXc3YMaS4yDzK9vk28Y
1gLVrUbGaR+ifUhYD2juiVsWoPiuB1/o/T0fEp4sjE9V0dYBGrOgwgmRa/C0oA/uW3JJGNaMkXdB
ZV4vg/ncifYfdaRc7OCuGrVKQjdiZxwuf4qi90JzbU6CiN3xKTNJUzQdKTWEKs1k1N2CJscRsJFH
g/GswOUUp5d81nV2PppuE2nE3heyk0IMcn0jR50UaaUOSAp0Ex3NE9ccEiXlgE+2GwpCItJNdecI
kc/r/Kf+9+Wx/wWGnbsSB6biHNMjqCx7+ar7J3ophCwYQAFewv2ZwUfX7RZEYuY/jtgvwf+kVCYI
idgzGJ4eGBJwqhs0vsIbLYHEv1yhvQrRgqohQQMeeEhuqsRvgW1TTcD1erlktrne6hpwVhvEbxJK
P5patWoPjEhiFMBAwmx3vfAxUMRwKnfeOvbLr456BU7cp9LQJxHkxZqEcny7K71nKfV00dUjr5dN
su0MPdN7CTxhqlJWD6LsFYmZRItz7aTg4DueGmpi46qlMgHtkvOUgtsUhzwTFDK4KydTuraErNNi
bxUKui+1t7aIJskKAr3SXK4U897/JCKW4vMPGsOPyYNGB6voaKv1krLq/WpJY3LAzmGZ9nT30LhU
gZXt/qWvgmnxGFIYEtd6HhOwgfnzZE49OW6CkntoacuOMhoGOVmu55b6oy0ru3sN86J0/g2YcUEH
xYiwzBVvPtcY5cMMKOa0OoVdi68WiysfUM8sni2uBLQTH1Pofo8edE34oxl3/qabaDk1aVCvS2QV
R6ZfpCHss6Fe3GdHIQOQ71kAL7tJWK0C2LrT6rQTwF7KW1+heqYtNkgytB3Ap0QuGSXzhUcbZ2QT
IvnJzNpvh59GjbP7QdVgp8TK1MKOWMHUpKfDKF7Y3TKuhdBWhtZquJoj14wUwBFqs6a+ERxkIxd0
SO9tTNqIUmUMAg2PE8W+P1+pTaH14CR9BaL1B/KHOP77Z/VPfwWb76mBK0zBJ4A30wN67I9zNqCw
SPQBW2irDxvDqZeViLE4oINe/WbCFbT7ciABIubfznJYNzNttyOHyrP7Z/f+ZHxa9f+AmiSIHxtn
QsQ/94kD7ffLWitpzkt0Vz8WwAXkiKOewzexrIIQ75jYK0oAnmaus0FpLdyyvvCjarIhtMJa7O1A
0D5TKcnOvGR3AYiIcLI8lXmKpKzwN4RA/+Eo5LI73EzxdJjTt8ZEdIILYYvS3jjdUnNuaRmDh/zD
dYptmsw1bJilmmGfPT5OMVe4xcHvFoHvsvK12rTsd3f1W57rs2lEB2xJ3UCTcngsYW7t4pYYwqQy
qLvDGLx+O97uZ0GMyRjCC2ooxkdM7DwZEXXNy7Sue6c96IUe4kO+pqzFjFB3v6x6ZbU910Gh0n69
EFALuVaRet8awr734CJST3VnQtdZcbeQpbXiPUWfUl+Xp/mVhaip/bsCidFLeWMZRYolCDTM4lzD
XL17DV83tPGkLVSn+TTGe81LAW+UJ8ehymgEcVSh05pTgfqN7Jph3NRefcUrh73ALnRDVCGqOtHc
4bjz+nLOWZnkrl4gKpXxQ4N041LmBUazusyWIbUf2K0KqsgZv1SsaSar1ERLwo9oF+VTqqbE60c5
5ncmRcq8snn+yIUWIPFfyxcEnASi6W2R+K4gwcDx6qnXFfPtn04zw6T06B4xrSX5kmuzTk07Wv9w
X9kxqo7nyw+DuX9aTvyu6hNYrIHJy8ijdngPSbqzbJZF5JI2vjIpMEPC3itfN8Ksjbx91HP4uvUg
JjwKYR+DaNe4cZ9yqJJzt2V14+uDrwrg3qNDa+CNldPXpUk0j9z4uFMyAFoZAcJ3X7HBs7F1KO78
ruGLtjqiTeECSri0NSLETGhvDUxeR79Fa7ocwomtdcwDdR+qQ78AAHxysSwEnJSbsvEp4EUBZNlO
xe4c0Ns3QG8joYoA/3sSreM0IzCLfhTXABSMLJOSkKqatW4FMCNhY0XAFFKQp0FyNZHDQRfoeQzV
bZ0cGP8KKteAPyfq+k1rY/uXJZNIAPdO8hh4/SoAM3Ky7cuId3IJ30jk3In81Sw82OQrjpdZ14b5
vHiYbdSxy4/9i2UIaN2y8Sn8gD/gzLSK0Wv2xdqcAOThiJLrWbT30MW30TUkw2ef+ohU79jQj8Kz
ikvQ+gCRNM1nGD783yc1p0qgs6d7qmESr+lpfblZq/kbi08YWNR+tq1uC0DWyDH6jDIeiTVv3PSD
DXMK2YCQ/TwJ+eJKAnGq/4EMt94o5gDe8ZF0jhFDZAjO09Yuz6A0SIV8WMMcWe2DVaXG3CtkcSzB
pglfjPXCHrbDJwzs7SFaDnqq4h3KtLxBuMmtOdAquHeReEgiqoPxV3gLKxSK+ais0cWu/tJsl2I/
zS0QmuABTMK767Szb2NluuuMS63nk/oRGRLxObzhqMIfxRyOY1Qy37Qk0PMOqLN1RAwIT4USWKzU
HvQl8kTn++MZ85zhwPh9TmjjUemX/UQi1YRGi/DxvdbO03GHHtTTHAs08P9IlegJsZe1ur+yifvl
nP/RGtyY1ozm/qFw04xXO9dxmKSooGhTt8hPfHtNGzTSgmNjRUK45Pargdo/KdhBdstYQVN55vDB
FjEqNMu/WfBoyBXzMDykkK3Yp7miZHjRLpBlEyf0PNcb3JbvvCtFKe2ZsT7OqSfbqKBjCpt83DS7
rl7iIEMyUi/Gyk+ZrQObL3HDgV4oad/7CkYoYP1ymM3n2ZEfKwcYedJJGh+H1rlifE5obw+5poQP
9kgWg6OkpsqU/ZAynRzjoLQAK+d06y1PHw17jsoiP+uOdo7pa6mHea170r0rRlv4yCIZFO5k5dQu
bYwrjSA7Q/N7sfEj/geRgvwH0s95r4Oo2UTACzKK0caDl6t86se+ArjuvrMVojpx4ibsMRX+eP6+
CL1rb4hGhNf8o80cx80MFUhe+uNtXIXMBVtE+a5WsDOkrW6Fe+2DOakL8wwI2kq8jeF+Umybvn0g
MdlUhE4YKqs9NTSdnpYm8EB7/GJpCKbpPp9f9WOss5WsgDvQhURYRrkdjYcU9G9e0fLZ0FO3bDvh
Jnu2Lqi1qsFav4CwLUGFPL/lwGKsVEN6EMb2MFi0ILMqO6fgnIvxbZ9gsRSfkrKU6FyEcq2NNUVo
S3tsME8iKbwQCOAmT11agmBwtsbbjvaMQRh0pGxQNUf1IxEnj91kqfeOoNGcyCPRIQnaJJX9OIcj
lGYSY/aLtgY2ygWKU91AKvLFI2wzXaM5oYXPE6BAlmBMNpHNexUTkBxMX7rWmjRUZY/aQZCM9yf2
A2QI3vc9uLQiUtwI9m++t3scFpZ63NPo1Vs2peHmQD2m+eylslhrwGyvYbYIhYkcA3FCuzFIoVLv
rTK55TzwRdp2AU+llJzPQt1Un5HapLYtttkpndalmvEQAPaHBqE/4Sr3DImPQtzLlSwaQqRG3sDc
5/lx0bwiIvjVFNJwjE74OUEPTJvKrcoFJbL2kEG6ZR79rIpBNnZSBNvqhN7iSyZ9edL7JsfBxkbu
ttT/Oi+ATSRrKyMK13Ks9v3fafgtGTGd4ro7m7sG+ndezhFDfYfw4n0T8v0XIsWxKKKCB7Uabxad
UEVPbQIcRZzsFQyS88DVjN2PYuIeQIqXCLcnU7l9jOcnKhRS+WftOujGuCORB1mJJvh97OJQ+knv
d1quUrlKTEi/HYVeLDTLGk4VA2FVu/48tR0+a/NYOfpsvXD+4ejfo7i3ObGCCVkmaRFSafq+BJ1J
5gGD+MHHnv7sCkykiAUi9Ds9UxRVzFDb4PBkE/2eQ3YKv++uaSydapdFSaCsXl+l1cMde/G1wIlA
/B8sjsP/B+3JZp3wmiFG5R2j/ttkSMUaTH3FpVXW0TRg8Qz8COVkl894bm/AmCd6Ve8gm5FpmBrd
Hco4fF/ehg7f+VrFnAfyAATbcE38AA+3z5YzmEJPyShl9sT2/yxKpW/18TdOk1mxc1tblAn/8RFl
XRvQHH/fI4dcwzieaSg4ERE95XAVQ4E6JqT/bULs3KGmNzk89FNk4+t+DlA7WzRxhDQnF40M9y5M
Z9P+7m3AnEMXJzXzfdKzgpE65gJ4Xb760OLSeYaJy+iyQnuaqYDulJAYzafdo7BIqIV3JL3hXKY0
wPvd82HAILInzefwadYmX0m0ltBXoH2oIRAC69O8IcEKdTjqzxwWmdE64+O424IZohcqU6S0bodH
zMldUHNpDhMLeTHCxIsNN4pJflwWC4MmisdUdB1DLTQDYGHyM956YqHjhxL1NUAXcR4P9HoqjhrB
/JwS0PeyZszvfsdwR7nkWyOsIJrC69/itIkIC/XZeMbwErjzLXv8g/YgErUPmI/vPVHCL8mk5ijK
Sf9wh1yPRyVzOQNbCeazOSkoKmUkrfYkRvuMDhL/j62WnXsOPLYd2rjd6NVvnatam5j9Hkz1XtRH
/q9BMgooexS2tKRX+Jb4U5UmBrnCJCGDiCFVJnQ0/Fqz94iLhqS4ySSLkRkuCWG9UVsIY7tE52Dh
WcouitflsrJqqV7ThJe4Izd7a6msmxwuhoDz0FXiAjqvVUq/I7n77/7Q7tiUm3yKTj9nwuSMVFLw
srxlL8gMKsW1cVpgH4meVvNuZlJk00y0VXJX2kLN6HBs5W8Mimj5XjZlXZf4Kl9/mZRz+JTOh9WM
+rhCEk3fasUpDjLNxFz7jxQhffrHPP8F90SI8Qaa58JbiDDP/lcyyhiGaNOSuO0niWZKP1GvA/3g
Kj/ExBTh4OZbOb1w5CB9yNk5/WR10LKp/54hn8SmagWAPmujG4ZICZlvagslfqu6a/c3R6N6ki/0
3CaJO4aS6pKPcgjwlsw+ggynqztLF6BiFRnBB/VMSx9gJ+bIryWe2WW5HVc1c33UL4N1XDDJgiAa
GpxgRH/KhyrFNjF6rDAjPY+labue5R22PUkr92SVB7LjHil20gNtp0Oj63sxNsKkscm8gIjABw+l
Akb5Mhtf5DLalVgdSmqG22FOuHm9Bu5r2nmOAhW3hiFH3YaKCUXjENS4X6HsMd6KVs1tM9o3tb/8
AgsBGbaZNhTpXoc8maxSk7flFr5Ex5ICJlLKhE8b9ed+Q369IsDOw5vMXS49yFDpvrX3XylhzENp
smXR39T/nKi08i3DkLJwcqSKZ2AJtrbb2DZQyfVvCou3fZQydqzJKwJ+LpJ+nxgYILkWYadYaMtb
LjFT3cG3nsf5+bPQpc2szza5zyce7aCdgbHE6LUv8awrAOa5N+KbkT4FKDVWeJRsaUujhAkIGvAF
HgxbkfhCosfYIBOWidZ9pjgxJj2hjtM4ZZlVRAgRltySt6spfnueZytksSVimxwSyZRCSmUjZJjC
Y165DhQ7rH4ptFcOV6UF2gLq//sMvNnfYb5ny0RjKSj+GKE/CEIQRVDADxTYV6MEE8PQPn+J2clk
PSvJbb8vkQwpZWKvJKmYCochrZ460oDv6oBTWEyuJF51+HhJiSf84FyCkVF0X5TAFAJXKRbXMdw0
6w4tT3OEEBeF5kSJyyIhBCifoNWea5dv0ULweaq9lpugC4sqn1CnBXThkvW+5d1Wq1sFWiSfHkp1
ySzMdgMiHWLwahqUhJaYFSTnHyxiqD2oFIHOIksT+H5/awXBdH5ZRROFsj7Z4TvKl0jgCOVIfV3e
a3j3ZuTBUemFNN8vioLUndlndKjMbbniH4eZGk2cLtTfh3lZ5SE1yntpxIrSEv1rEcLDqxL39esl
f04jmknF9CkLcgdyzmKybKRkUigO9ChX5pUx/oOPP3AfJHPEeRD17/z+9T6rY7vGHNSYwi3tCScC
8xyJgZBVpTAwDpkE/+TRdKyoFCjVN9tYhRkLdB2V/1sF8FlXmCoWKFAMiFGNc1+uBbcXLTluxfRl
LddPUue0d0DDCo2PifY15OV7j5rncWl99FHUK1nDk9yt0KhjtrTxtynPa9PexF6VEGfmKgMAoAyc
q/dTUvd/1wQXcIPftRCGG6XR95HYnRBlwjg9cATXeiwgRNjZBTI68GtLSiNEiTLHgqeeVkhNeQ2N
pAvvooEYVZgdTnMXZwtobYaUaEqPcb6wvAEMw9/eDX8rk5BfA4edFh+w88vPPau4IYE21FjIzaQf
+BYKuRX3lcPCbnIlW2qDoZeX8f6Ao347JJqQ1iEHlBmUlzTUdKBXjRdHr2RT5WlroDrvvmOQgQo+
HVWCD2OStSqaWkhO6rRiOh7RiRJvPIQNAWVcd8kDBCakAnfN4TYIi4Ncv2Y/GExINFWyrFEDoEM1
fMFTsThFlcGM8Pd5qmyrQUyFaD6s0YADPEryHPmhOjaB481zfwJMnV/0AqNscRB3E4dXo1y29ypu
qtvzMtV+GUPYVjLsG5zo2hx4tTOYLZfQ2PO1Xh2CU9CJYYXuMUaxFzpr92T2L8lABao2Com+Wzx0
a62aISWlxNLSY1jqSRHOWtzyNXtBUevDmuB5hWqeIELclOkL9BEy3HxXAXDtoDPmpATg1wzHmTOo
koJ+6MWjqzHXlsTq5sw7PI6QwpKAExulvPd4ApEmQYqkcQm7kZMRCjE6fTJ5zP+k8cXrHDQz+RrI
87qlnqINJBCu2ViLABmE6Gr0lnUY2BdjUN6LO0SN9gvJdHil8LjOGRc9JCbZDsg2Rb1CwiGP0JrE
h/Izt1uxicP2zl4kH+A3v9eZ3FAhz2+2ktP+uiHNd2iJWG+e6smc2gAzyVcBWrBLMy+nvk4ExhZm
3tyVgVzIMUbgt08gMX5bYyMM8dutSNDYnYwpuUtUoQdMzDRrb3qiyJyK6hhZTdeQfTiT9AEGHAKM
oJ6lrA1jPgCW3qrbB5bdqldYke4BFyBs2VkeOWNzzNz4qwi7/gm61fYXRXejVMUUxEGbNj7jsFmY
111iScypdbil8JKQnz2hgK3o7VdEV57h3UmeoKtPHZoIQr8ew0nioLTId70wyuLNcBqTVfmAVwpD
rmbuzeu51qKYfB5pnE6VM8JNjMipWpGxGcyA+1bcKcMmOj39Uk5Q+09CLSqfvbDQO1tNVsT0Tkbg
x/ydK/WfPLGUkMkb79or6V9Yk+aOPea4a2OMu435HTR1Io4iw44XNXcc7iXsOtFBZ0vS1aL+JhAE
+eabD+1YgwN6WEVWmdGbHy2C0IGuMZvsGvRt3nzEUNGhZ5Qi2+VMitofNsQImRjIg9I3e0x9jHE1
IHO6akDQXQPXGuL9lOgI6Y/VxHnWkkTMGOeSSG6gnQVnF84Wue9HNZPIB6bw5y/u3IGMBsLCXklJ
9Up8KfvTVRDrjV0AOQNg9sf4gEc3xhgNm77CdGhr8Btx35eNs4Gyd4o7K8Iz//V/ZVPrdU7yQlCD
jyRONjWUGkTXIXQIqyHZNXcTCW8nNcaza1jvRyGZJqkSmYTFqY+VMcBbSobvTrzU/MfxgdrqJGG/
nxu+dmkyWwaP1ETs6NDCriHbGcasRlZVY9Wb34+OExd6gCrdMyybOvtK30kCR9lyBJBF04g10Nzw
QIlk6q9X5RXegoCr794R5cnUt4MyHL7ZBZILRJwozKTDOQYUmlgMYbqtAZFqBY2Casp7Q+GIgCjY
om1kAf8RUX+HorvT2yIZUMYZwvXuGLgtduXtv7jCdCyLtJxOAGXISFN6+MPKfY66PMiCsWsbHIZs
2PFnLjNxnudrzy01m0Tnc+BDPw6/jLoZr6YMhn0GpDvw2+VnRpifK5BZP3kmnwEsOd0APshQwsju
5wrZJT7/DFvsMrtnaEtEAQ70uWUCvpeM8pYvupeZK6BMAkkMUfCGlRE/QKxMMltWlxEnGo9C9+l1
v0qcD1ewbQENL0Fe2Y+Nxgl/PQQUHnLO7QPX11+d6dxn0YJXNGa1xypiSyejnI/6TQut7Mi1+oH1
CjvXlss/s6SaD97dUM9o3aOOIlWDGajtQ+cpplCjjezvjBEfVihGDJzRyk+uqJg7aJ3Idh1C61wS
t85xwrkGBxv56JPnQ35afANXFBajT7I8/DRCRH2MBpm68aU/mgwxk3zkpshNtES13bYIvKqVAq48
EvlsaRwdyYfsb5dbGlTKGDqCEAgQ0Ur9FeSRYc4Ux/0jMRtdkLVxPCWQ2qRzY1FOCdaGsqaSje91
eT+D/e/I85iPpRLpRuNpeMBHMlnpdqm0cwbVuqBzCAzUmYktxZieQeXEZHziwlxtPNsxq3VonpPb
+lRcJmbT/zgbBi9kvhwulNIms6W5dfcUWjxTaBed6tcGwQ2q5tV0DN72eqh4D8ZlWfIrQ7V2N2s+
s+ke3p8X0XOX/wvrZBFEKsMJ5DosT/sNhwOlrknbgDqhQQ0AUgY9GbVLbdWzqBHXI1CRTAnKpTl1
yICGT1oEeswGzFoW8RztjXC9h/b9P2xzk1kG3WLWeGlAg8wxp1zedfl9FO6D7gTNzN/b1jqQVTKx
NPA5qxORik2sRfYS493jTHSu29VoN5ZC0a4qXia3ozSBEbY+bNnHWaC3I2jUSBVnP3Wc79LKUXgq
AKGTrGoEKT9hiRxyO6Y/EgXkIr7QYuehoFzgKhg/uIGlgZl/L6ubovHslqlWSGKTCofiCvk9e7CW
WvnO5NI5YNGHFmxemN3xeBpWQqdPsHN3st297cnu1E+VH6WCxT7Q5h5pUEGKeuMrXmGfLBKk5MLa
BPHYyG8UHHY7SYQe4IsqMo4zsxKV+g0om6SI5C5tII81uKsbFZ7ihLE7uTcoVy3jUhP1EgPVCgf/
qE7lLp77F43wv499K55hBiQeyujuYMeJJSG6/6QrIqpY8Cv5Y+xETLsnSv9zSdWjEUtEKOzQZ2HD
87lnZ7sB5RNEGkEFLK8u97TVRJJ9u8K/JOyiOGMiUiJR+Ew0GQxZ+t9Efb9bzdMjx+hjVEvN8oUY
f+5iigrMNPqyIOz04WWRWExowNrf+ikR4s8oPjSj0D2JbY4SIS2wG8E8iJB44swc/1hjdTiIZw9U
S9dy3Tn+lbisvzIx+07Nm9vLcZqPWXqutH7VYbHF7yBFCtN7/quNHLi3WqQPY1HRIGBmq9cHAa+x
BNJ8V8jq0fBaLXA9op+2Wz+L640XFbTVRPXJn1P9p9T9pcttCExp5AfNTMy6LKeHnb+/5BxWHPdF
X8OcS0tEcE0PABy11Q7AlG1ESEMceGR9WVcCfFK8vCmemVt7fNzKIaLKbNA2aqyNsi7ThWpZLC+K
xJZrq2aXnU2xWO9vRutk23S1Dpjn8if6rtppMFmmwomTaZyyCmPeXId/XMVM1wP/250Ai72IxFjG
vN4MzuYABsloL49aYKAP0qDSk4xpY0VtDew2GOekhTq4gJCRMSIQDEHKZ8tz3XRWQTdsR/FIf981
/GtCbPTjcNNFEwuUCzSVDzZE12upiNQ3eUmUMtanZjmoAckOjie5ZEFPK9US5DuCmidwL7HACsMy
gkl+z7VgDXGS27M7ksD7757a/kRDjQPf3V8cvTPmH9TUgJqAUoRdhvA2pRA39H6sTLfUpsVtG2vu
RzBfvCWAMcvrKaZk2BtSqXhpAqZkhn1+3VSyw6m/YQaH9RSZ/vhUQKCMIoWpI4Nyu8KNacuIyu0D
6x79m1cd9BqOBmPK0SICrbG3JcMBjLE1CRiywLalnUDYcd08mvFLkwsKj3FuGcZL2ky+t12c+iRE
rmEWSrKqyBfSFdIIa2JReDNVZYva4DlbVlpghexj2/B1erJD7ReHvN51+Hq27cD1UH2hbiz89TQ8
OxiEKIbH9vapt92T0hjtfiD1GWnn+s7igdUhxV/iGk6aeHWkLlvzvUxnAtQENSJVrrnXVRoglGJF
02Wq96pedPx4jcBtbcl0iJ6iYhFGepZg2SLAr2dqfwTgHUQk/WCT3e/LTuHILX7w7GxTbij+Hdg0
OsOJFCME4auJU13f0DhPGwSPU78GoOdgIgbQxtZEeYbl5OFgPVtan6OLnYnzGQXf4BErITgiY2Eu
8n2IxiYAfBzPGl1Oh+NYMSgSQkHzsfyOrVXqipJqm7SXBgyHCm61S3mAo2vo/kfz2iHydwCgz0hU
Z7PmwMMs4IMC7ISjS8Hd41DX78eC2emQed8AbeuDiumPkwBn/njFYqe9iClMQ8w574EMj9oFdG/+
IOIU0motxxNFjo2U9sla4GgTN6ODBR/yufu8tl5AHqWHtUYcY6Xuc2cykCLaZBSqH0bx/09ULlsE
n5BVxNnp2tzH34IjM9aeeauDoPenW94yegCvG6/Kle8GuJwa433NqSKoMmRspUzJJGv8exHV5i85
9Vm3yZ0zqoExB0mmxKsBhBIjS0liai9hi828LQHEOBnrEll+DlhuWV8wX+9GohSgH5YZwlneRMjS
s8++MC+Tw/9fLWILoMgmNJGWXZLE3YQqVJ1YyuxRIkvsTySuzFR1qrXamJG8+OAqKANJgQey5Pm6
8LA46eF2D92V9a6eVWwzje2jV2uL2KXM3ELYAHWsKJVhbtMAM4X4MN9kAZFHkOODPkqCq9Eg/B7j
31d3mAyLsfdTFU5D4OEhQGC7BuJqQH9wnuv8g15tLJNyjloNQhA7p9D7trePqFCZ6VdtObh/9W8d
znBSnL+PVZ6xxIU/5he/r9rmBDtKGtmrJxOh4feV66LKei6DYz5qg64A5s5LstEdiqxV/BDyfBNK
HDxqRZEbdPhmtaYCqeKPh7wARi5+oasLm3aPs15SiVa0a0JghrKvFCoEKluwLQwiLYenwy+3bfNo
RTf6H61Q9daAOlystvEBMNwZ4Sr4jWd6y/eO88hqT03NjJ15OBWSStfR8LxarumxxYXMvD+pZgwB
GgeY6b2UYYmCrZ3uMe81nOULhZzYIV7/1w+2n65t+Eoy4EhufDuIDED7kMM0k1xmPFOvE5DcHuAX
UYFn0T+29TumyQV5k490Z5fcgrk9AIkkDklnOwHKPIrJM+U3xc42s/kK5lIIUoMcnH6TBf2RZJct
ywmUvqPAcw1DQThJQy5ufCukSPc562kW0Q4ZGGmvirgG61KT7VstPNgvRcTp0HDioENHxNlGX+Nv
SPcgmmik1jRQNATx9jctKB5wsDUUIT6L7g1oVjqdpIj1Cz3xeUxQaRgrCpHTAQ2LC1WmP42kcnPs
A//FoNJXTpKX/PC4vJaLHWLXDbdz8luEj90I0VYnoUFXOjAqNhEGZEcoiBC7AFKDnBvO8hV51k7W
+hZV7RQ6lNXXzn1iBSNct+q6dAB7Bn20JNsC+M211Ku0p6MmDoGEPaJYe4Yh6aPLgZL70DyGpWy4
2+iuky89BzvZ/ZVLKCZ/9zP+ScC7P9ZzEuXSIPF2//m5M7WFGpl568MYyDi8vwT2HVsdDI+3E7dY
qB3PhHBh7Nm8/ppOWjOUJCclD/hrKFZcga2UiaNGTsUtgbuwt97m12fWGkfi+bCPgczcwkSAB87m
1OegICUQzLqZZOQ24cGRRRExhJY9vUWehsji7k8KRw7GLpDnQVaveZ6lAikDLTsS24GPRmS/nrUC
rB+SgiCldqrj+hrny0M+IyOGcJfU5whNqlx0rrem4ftcLtd8k5LqQJ4VwF6v8fLWm4z9eHY06Xe1
neHSx4uoSsAIsbQ/Uvr2K1PTtOUOqvdtUS7xpxeKFX8qFOwmsSulVYg7akrZgtM6kE37PtJHaWAK
wYboYDyEt05ppLl0kI1hN1QZ5urjvgGMK5AyZp0QfNeDsTSiM+OaJdjo1zvI8mOvq6IYxmRY5LE7
ypRInZ3kbL5zMxvL0ehWL9v789Xvti/QmE6Xji7ZZfMuiQPV1TMWnrGv8CMR/d22+XqnrsOAxE1i
nd5nKecJ8yQGnjfw9vPocMNSUX/A3JQf2KNeqTFHtmTenQvTQjNx2swXsJq8F6elmfdMsNo6J4+T
67fsu8k4Ms36cxLVf7w5332nC4Yv+56JvdTS8fYDp94Flec1LbhQUHXxoNpUv/dZ2pHA2/sxUvkR
cFWTnrfg+SXN4UYfh4THpuUGKei9tXW78FOfSyzGR29aGVFA8NLasoKziZlGz7trxjnAl623plex
y+jzIaHJeuF4u+UZG8SvruGI8I9lesnBWVfvCv1nb/eghEVHV9+tlODzGEgTTvf0vYkdkTJw9IIP
IdaLP/FxEYoaQ6bKDhj5uGBC17noMw9XX9yTv/2i6i92UmUUW7vrixEqrqgFkvSdM+2EQB/oL+Ou
zCFJQQQqtTteIuRYxFIl5pDW98MxCHdKroKoIMe4FZUYUUqfURLW3dEoF6/vySWRS6NdckjlgeLR
Rk8O/ShrDt36PLlmFDPznwm1P/UzRBfiej7Ia+g8dbA6VMN8vH8R/wV5SuWnkyZLKHfsHAikmR0d
U3BRZ/13fSZ6tFQMUf66UPIY4vmyh7JUv9EnphgaPUDpNzR7slRSjOd764uXpi0xydkZMxHbBGIw
Qb9gU7RPP8hc3GyS/KRc0Cu+27geBedGwvsASa2QpEcDMzr+mbydyQk2DIsPCAIdgYsUZzic/Rhs
NqmFT2EOmoP5yhJRGChp8ro4rpvvMS5yxVrUSJ+ltQaITh1IZp58/aCk/CBKgQ3z3IWJdJIDL40/
u0lNXd92AQqPKz/sXd4mm1qmmZFuLiOU/2ZRmf21oX1o4VA4qFZ0AAmrhygi5RGdNbanFH5lR3y8
HWZUV7oD0feCPBj/C/wyxWXUERyeyYNPXYWhBMmWaa7h4jLuJp4iDrtodV90Hdg5TVMyUm38EjLj
u0kZxqTMkU2l2j3836ivSXv99/HMGscvHQcHNCS/CPQ+8Y6Tt6LZEKJsD0+AFMFLTUtG9651grjd
IAXOz0ku9fsWvAW2vzKYA/ovL2pRID7tsqnGazVFBOsLiQhoGgIvz6P+cUTNkxJeOnuXKPMUgGq1
nAUqjcdiicvdDqLb8uuw6rfXZ+86BeY2uPK6mnlDC43bW/1/5sGG40tqbpHHTR05bPDc09WjpIpq
+61uVUlNxqU8OLfWHc+jVSpG9JCRMexE7hxHzfip/slJN3Kl5O36HacMGqAe6RgWz4603hpmi1q5
6GlOoTsnc3MDr1e4ZJ6Dsf9EM6xpxxojSGR+b1ZFI4TRG1UGy4wkTW6/LScBDmcDnUKhiM2uF5Rs
r0KUpIj9tKOkSN8shI1fwrYATZdc5QH4OHPTU3oZsOXf9wAJQBOeWNOQ9mC5xYJCDvFx0NmKMmg/
6pY8WggEiIMD77dGsNwISnaOi1blnQWntSztw0lK5R0GSpgpeiGRNE1k2HYyJgr5Esa8DksS4V+g
KvfJSTwIuErcyM1uzvjg3hkbWWnoKRq/lLIlRmF3PDQEtVpebZTjJ2pOWAGR9BfMaMBeHyDCfNci
Zad8qo6LBfsbRDSyxdzkXZL2VJbR4iaWCKIPLNs8bXEfB5PczG/s9bMRnJkpnFXTAQMLMi73WmwO
wr1s7QpxfBZZYFujblNePkKNbykCLngCCoup5QrSd6AfAR8MZ7YF1Ats1Rru+VcEKMpqCtK8qNGj
8YVa1C2HFvnFfgvULCpc55Uv0DeWM5RxonN2kVSA4nbSW5i9Jar1UrQD2pg6QtDb4nZMkvUM9qFc
G/zf5QsyyqwQFyRpgmmPnGy+HhOE23kNBcEiUTQ/LscuYV3HyUFRGm5x0M7AUmsG21/hl9Kqk/Pp
Lch8wXvD6KRRWIUOh+K9sEfrGQahtjFz7oI5bOJY7OQc8zG1R59n3VakERPKuil9Eo9LuaQOLqEr
pUT9cckhSDxfEKtbu6UHuqDaCM0aKjN9bUs6VLDVCOM5j/EZF3/DlsjD4FW9z93vzHH6Eun9787B
VBvjsx2976GXdw9gASWXj4Yoldf233D855L2Qs9BevY1Lo2MNXgYun21Fg6KmFZ5Fonz2eHBazfH
1zfI2seQsswLb2CPQRYL7XBu+yoWA9Dwgiuh3CrD3c/5ydN5Vxcu/QbSyGWU9NTwpe05ufIz3tl5
DNnNKrimBgqhjWlhUoN+pEeJTwdD491dUiqzPNQNAhqTM8csytAL1ZcgstemMOex97pO9L9rLtwS
liXngLpWDCIU8ydb/KfORx0lv7MIh7ub6NcejBp6JrQqtzI8Rn9UcveLc3VsWzfLzimhHhuezExW
VsgZsvyG5o5VoUh4FNFykjUe7f/V6ZvlqqlLoirvSTm+4Mj6b0eTXqLl0f9j8n3miPHc9HnGk3RI
YZDrfaMjCF0qKQuam/U8WPsVHCIC3/E7DcRF41gPE26mRpo3RGKb+TrZ8JqaOtG5HMvjvGzfZKHQ
YgVKojl+2KpUiRfffqQL711PVkOD/Gm/brTlFGzg9GXMUKZZWPBswGl7GFiWlG+k41T5JVJ9HEoX
KuYxdJz1Fwa5lZyJuHDXKUaZ6EQAjxDgxbeEKji9NTQufxfRvQt8RVUvAP3GZ3QHdF6cRzgSbCw0
qDsRx5IVlyL+kso8GyMOWYApz7NAPv6+Xs/qStG4XQvzFsFVMDv9uk8n1Gkt55i/XrHitpol8HMm
DM6RbnWXBpwWESsL27TmEez9rCvcQ1b9lW/MXyKwDVEXZqfiu0QdTObEd7zGiQbgKlahL0InGl08
c+Uiex9s6e7OXy0x4MqX/5I7g1mcbK9yMVZpEyOVmRj2RjPCniJobErgRRjyLtYPtz6jKp6ek6OZ
37Mt2Cn+6UB4n/kv8NwAW4KorUoPS/AVEbvzNn6zhKI9LCQoX/68Gq9V3lM4UbnirVKl8ktSGD21
a1cbZagswEK+QMdPUPcaHqUljjAz73DLPJOiQRgh5Ebgliy89D+YWzm416QFPciC6zcVyscGOCL6
QmtFpOhUXNYtz42oDxoiPDltQ0ZHJPsFaLRebTt4b2r6XxYPIb9ccEe0Jhlat3Iexua9qjrnTfWt
dlWUmfl7/aOfZm0zQ2jfowrEEW5ff5F89J+B8eb3x4lzN0YOgt4C/F/D8L2BHrAMg9/v7R/cbC1d
jPy0XWA126v+NF9eSMmi2iabZW3kCIPSAaFxu+JdXjrUD5OWXaBjjdqTKZd6iISgWJ5AUsN9KAnq
9QOa18sNmRE7Q5QeipVzQGKkWYYKSjdC2mveLidwdis2WN5/DG37qeIobslIqhcEPkHu+DG8GICP
tJbikV+eVHpwFdY9S3UqoEIcC3ysI/7smG5QMFt2Klk1P9HDy+cQKUuPqw7rDaMhHyFipQqV0nyK
wgXOprhL92tk7wyXjL2WhWRHJTEqLvjRn0UAx9/WHRvq8xSZC/uINgKP7u42BWdLUrYEb6kxPp/n
bMu1U6an4su/hFi71u0YHjCmvgJgL9pyQhNn9NOoHLrwEl8k8eENKqio46kEyRu9rzky7KHuRGU7
0Y6Lz8f9RdIVHuxxBhaOH7Fhy441H/I34UVFqMV93Bb27mkYNgG6PCxbgQubSganKWx/Ie7EqP1Y
aXH3XFjvedwebeGivxRO4a9nG7sLp6emh+0R03wfx3kSytCEb2SzeaAW/Iu67QPh0lLoJN767lGT
NyjFTBic7+Cl/du73RPyxVp0fiV6Tz4+hpqjl9/FIy8sflVpNTz80SMh0csPII/LcsVgtQ2lb6wp
ysxoZ0nTpHZwZvsd23Lf5AFNgTN3EBaPlZBITliu2KMw+cn2HvCOO4kBi+qwR8vVXN9dtmyXnXct
zL3tQwZ4iItMl/Y57b/P864BtmpKcgu5nlDWPpIgGgf2QoajtPjDvEtPFOJpEeYycc2Q2BLzKzZv
eUykfV7R3EHYNoydq20SSSaXNFWm1zplTMzdg1AHVW1KmooxZefXocYFaIrhZay6vXSIDonMvL/c
jRnS9is5YVNxFxq+d7hquMsY+SAdxjcYPIR3qxJ5NiQ85fT+zTmWWHsDOAwgmQeV6zUEn1IyMrbp
tgW0yv/Po8zGBUxKepaEdC1gnPlfBNbazSgIzOOda0SraKMLjAU9hw/zR2RKFUanz0QJ6OHSBFgJ
yhlyfd4rZ4YlsuiCd7l17zpIWTEmFgawoT/s8WWdWf6CEFTi7GjZd8ibE1hX0tuTSPzPpcLdwGbw
Rq9qi3F4mPoGcTjiPXeEsZ2SW0PJGgBqenJXxDX8cnY3Vxvv8VrszlPAa547gCznvMbhJsYbFYfT
p+l/hdGIOwqOtstfGx2NDICSc9NTWikzFtiv1/LSb/lT61+rGCfOrumEJT491Hdc5Euc1e9ng4Xz
z5A7PUI6l3qdHVnt+qwWsjRHtew9tEetQQy/JfdzAP5sAkPEUa953KDDshXTfjPV3aNNOJQTIO03
4oMW3HKlDk0aCSjv3bzXtTUcYg04DDNhv1LNWEeaNHPbZ6yjeZS/xKFEI29OXj/+eMrY9zyg0ius
4Ks952se/m8hR7k204gtH8L/4RqPQlRCFDJfO/cZpupd6GnzRbq0k8+Kg9+IgVCPHnQ2OAtJveSi
NeL/55DgiG2K+nQ7+oMzX3qpn/YjrDElvy1BVfR1f3z2ECIEdSFYctH+pyf4xIh0AptRcRV4EKYE
E7uN+PJ3OhWUAQAVZyeiw+24AweiwO0xlYzeqJNwSzoDC5GGwKBrARvwNU6GECS90dgf+cdyq4li
HPXfx1+3x7ALF7rBbV+aa2WskYukeD8W60wLhj08bYJ0kiXVf7BBWbYwVFm7qydP++Nvc+jtq3rQ
Xw5ocYaOwKCujCqYjz2os4pB3Xc1k2a0Hc6tJVfVbttXTafcccOau8f1kbHHVIGAXB9fgZVqvntY
STeQoaolxVJnncjwOUw8u9j7KQq8T0yRWfjX9J1oKinjRAgM3lAzCir5fT/INuPhZP/P8vntXnXG
1Bu18zS+kGcmK8ThueDs5CtmuOnOxCzyO6aj/pcj8d2p/NGPb6jN5lq5hxcV/Z2W0ublatfilKwK
0EpXc58mVaJl2aSgLHGVBCXmgt56IImQIZ9n2Al7yty2UrnRO3zwl6szN7ZIPYlMGKW+hf1AvKFK
kbd8rmwq0huC1j+BLqM8qZ4JyupekTH/Nqt8/FHtYGdE2Ha00a/kqzl6/CUl9fbbfeX0NnPLCwIE
k5+7FS9FtclApVbT0KYWLtpQl2xYBua3gI/7SGVJUQuadEiKoGvya8rRFa6apGbKgMT23SzRN7Bw
77EYjBqfk16H/cWv80pEmIINWKS2P7JAvAk+RSBJZMaGp5OSbZ/2M37TaWGbG7hO9jX6lYhHniKy
QcscAMYGuepawdY37rC1wP4uVBkIXSJggBuNs23UhqAkdBhkrQyBdRqSBencJ7OqMruni15THO7X
2jnyal7qjlvSaT2ki323Qv7PlWHbYM3fFl8tpF5nH8fE+M3Ma54bQlZggi3uXjq3qP6KAgvU7f4m
JP2iZgPbd4deat/jQUQyPxbZ9mADjOEzc8+OGSKAJaQ873XniRFXPykx7rvWTvUJrc2YgMYmsfom
mdSAy1KcX0vyNt9RUgBGfAznyyPqTIiL1jy7W+8ikjY2zChMMuT8QVPPI+HBOaxow0lkhhe36QAz
ZJlDzx/YTH79d1Ux13Ln9yWmCgKkTNBYqDc12rN3UQyaoVVimE5xZOc2KQZPnwQB0Sru7MTvLPuP
pSnIsXcmh0gSfEtDXFbsykDdLFURIMKdd+nF1LvxfivjXSy5YUzCWlrHFhWFm0wUpGM+lJdYkbA8
g23r+OmYDHdqizfsix/VRnOY18wNFacdtv0BvQmDBUkJpX/wSCeBXXb57nl1R6lqJVfW6BAicifR
UjUf9giKfDQe8ycXnZa4DeXqUv4C8DINQqNdfbjNVBHNltK1Mp9gBOQAQ+vhTFw1UJ4ABXP9Uopa
zBx3knvhnvsJHZoLHBypXMYv+auE/DVKq7WVUuickmQ5rFbDzULJe5Aspb+saG62YK3Vgcza2aj+
iRhrBo5Ok497t5rI7EhSN1b579Dbf2N8hTgnjTrboMZLTADY4/3GL26kxPnsetKvJUmghQ+CbE0r
UewM+m60eAMh9FNFfI01DFFJt4byJ37Ahy1FNZQ7EqQs69xqMOc7TyoYIqEFaRc2w5Jjy0NoSyzg
525R22WEXQ3CYFOryXH2nZQR7pU8vK7s/ysmOnH36ehGnwgd3h03z1yzwH5lp1sBMiEwIflq99Nr
yCF5aa16mM58rVsf8jl5dZOIei2l2gmZ3Qvk0VMLalXqHg/AFvPBF6frX0SZsOPaZYyhhHwm52+v
/M0tmObQryfkuB+eip3toTcRKdi78L+Di2xhvTNf3D3p4HHZZHCgAHwXQw17Nw20gI9IMS3ubaAW
1aoOvdNFZHucWZTrXMl1lDss/RWMnNwAmWin63Iht2E7nSJQX++4YHZr9OYphn1oEZoXzOPBmSRE
h8c7cXMmt7fVad0hM0xsCaK1nYmDi6FAvsJGiJGE5KE4PJPtL2KdKCQ42aC+EnUOHN9OKJD5LZsQ
YwPsltxBcYNqjtenerAEVcWwWzHgkfr0o+RWZpukYqwTmPYT/hsH/yHAVNHGZSxvC4/dcHsEV9u1
PZZuNC2yTyOyEA/ZZuYDt4nZ7i97e2jFKG8FND+BYi1rHeA31geEkuJc5IIaw0xGX2JIrC46AzBX
DsXrIu4HPDUeDEjhon+ltryNXvOAr6BoImqj5IEc77/wtc5512bz7K4lMs4z0TSrYviDvGsxYZyz
wYZVB+3Hqv4K4B/fiUdib98v5KBSdl8Q/evO7Df+DoI5X5jEaxLU1KByfdZuakEVm6W3i+3yZnPw
eI02bMsYONJcnKiglKUf7/9Qa+t3SRjyO1ILx7U5lIvrLqd8pTbO4YiyNNlo9GYAa2U07Qq4tStE
NzwZ82kfTeo2DX1EXw3Q3btPinMjQyjckoPXQzF+AuZDNweVDNRW+U72KkbUXanEkfnhYZKfSotp
Sy4FqtVYIQZxbVBTfo/Qm89KoGe6YOMMPw5atlgN+Mr+5SbYEWv+FACEbb5+9M16SQkRwoNkLV2Q
CntUeF8j/85DseuTfEvNzhQr0y2wAWfmppr4/b9doglQbtLI1BzUaYlnqPq8nEIIsyJmZ235GIIp
zapYxXN0mGf5zNCZ7jzTQVVThktLK3zzSXPiqEyt58EkzgoWL6gLxKjtlgd5YhR/cNE0P/P/dLEz
nPZjsr4Vt+g+K7LhHhbnV4MtBm44iWHQTG116rdopqBvzZvJJ35cDFrna83wVBMKGoS5ANMhZV24
QlD71T8N1cRr3hdkjIgm3aNwaN3NddiLjmNwsmK/xKpOrYO46t6h9R+n47lk8CMz30RnTgAupiHH
ZTAYCDx2UCBwfNvZlAmpIQOOVyngrEPmHiacswclLqpDIfI4eSaSOaSJ6gu4OGu41pZhVqClPC0l
kjKVu0F38irZg2JSQO7/vlC4tBl+nKk6MWnQZ5XdtbsJ6NQbHJHUKjIqC0zaony850bAhyduz8hR
g25+xe9kzd9q4OjtBMgpxxN4x7QzFMkT26q+zk5uvungmYkG8bocZ6WCf3z7GjTBhzOa7XEbmfPW
ZKyw24lMmGnkbUX033u17ByRlfDzVzr4f1vKW1qQQgDCx/4A0dhIv3FKsyET8YQjQBCxc2XddixB
OVIOF489wTy0OAUMYU2ZIMVJtdw9SuvCuDQblV/XawwNhrSSNSv88rXBn9lILZDENJ5ckVYVT6Mf
1FVQ50UP7AeRrEKG9ZK7OsUyH5DSdqXVF+J28koXNj586yiv5ENpNgk4yy2tfTPQLfVla0qWWKUT
j0sDfWgMdH8uQDalJWfbG+RmhBzHEzj4NxlU0Qa3yNO9KFHbS4HZGMlwnwXiyX/oSbB5cylQ3FTk
r61EP01kHG8hw9T74MTMS82Wf7+GDNATgcWAu9EId4G8crc9DUWZSX+bpEcTU+IMMTuYkuzkuFFn
2dPg1jQl1Xk52HNS8n4Lb49QVtTV9cjoUSW9YtIRmhVNOhK2VRXOIFP2UJvPDZqleA94k/R3HtqH
P03wy8xGkBLo4dK2iD2uEMQUOLZQJX5BGfTy8nn3KDJuuxseD1MxboHUM4xSdUhehXE76QUZa+aF
zKJb9e1OXuR+Jo44a75K64qc/UXFwXypviAQ6KxsAoxBvKlKefHkUEHNFndas+Eyw7UcjnWzmBL4
1FT1G1MuaCSyMga4q+pLWIzF6bWWRzPWBEeCA7GsOh8Aw/onh3dkXLSFESLmlE8HEx3uIPMM259L
+u7qjH1vt2Uek5anDqMx+y8gFFipBcZZJgk15kShuNFiphEMThgtbRvx4xZUSVL9V8un2TakY6fa
JjUHXxKeEw7y4bmiSZT6gZUjjYrH0+W+FcrdFXdKgWMLU0ZtrGoNHUhOf4LzIKddwhjEMAEmrGnj
K6JI+uAgOLT+lmK57JKEHAUhWPkeTJ9Ydp1BtLMcHQYIMa1MKPEQzYxnm/M2beuJ4GZ34npR1J6O
YLq75zyMrSgT/p6KMld2ojzk+7OwANCFYV1XktLasZ0ipLFR3uPNUExBXT5LaAaPRC2aI9id0Gr1
19WXqhi5Q/VyPABDw4bdgQfgF6LJmIhIRwflCwZsf4oKEdsNma25u+XAKPM6PPyCCU9ILrkMrZaA
wqEqEU864Q7eHv5zpVbxO5rJoniFSq/cceOCYqX1sp9qxYjD0xE9+toDVJANb1w2M9BHXz8JDnb1
A9f7sTE5winIsm25AdFL0vXUYbGTdhUvrCXi1bWWgQi+QhqbsxGHPCScknHuyi0DQNnyTki+1S1W
nUuIGecVLLyRGnBbCDt/pUDL20r3UPSxBmTJKz8B9ek9yZyixW/F2FqLXY9KS8g1JLD1D/LTGvA0
OBeXXStD5K5J89P3CAHrYKkHveNyKNKpBUUcWWub5U+koGn+ViMrJis4NeNKokPaQCHOrK8EZHVd
h/SPtqafyg32f2f9pCsouforSlSCdpAJLYsBv4saTqUZn3ofJpxcHRXH5lCkm7DYkNbzOyp/nI/K
c2JdysUF5QG/27EL8WF6PzuklWdmF8i+jM6/0zDLCyF2JnhbeSvc6xImvuPW1zDcsvSFhwoIE5NW
ErdW/2IMpVqFh0hOmP+RLh1xdhKVYl9lCGRSfIYGRU5GzSpYf4E/hSb31jm/hIvX5NnX9k4UHoPc
+wwtzBah32tAayMAdSuFGiZDbZ+zqkyLZ9thC7gzlt2l/GbKZ8+deMR7nIL1Xwu9gpG8Xh1LgJf8
+R5tj10ENMUQbKRbyzYI8c56KGA1H+b3dTYQi4PHlEro0KtqBt6pLrTiAoAXI6ikcXKjB4W+5fnB
BMl1TXXFlATNXbTMgxVbL4Qn4QMSY41if2VX8bHQNvoVy5hpQ22cgUM5LcoDdhkX71kl/wq/BREn
iJMffLDCF6srbkKKqs5EMivmoFK5FKQeQEGExPqmrlqJA3DHah/1mzFbtGthO6ATDcALueGaB1Y1
NdqwiBP/tXUAgqP1rAr4jYIPglxE1u5uC9vSWALlW4Cr/zwS5nVKTfV0bQmJoTc/n6mga+rHjwhh
D22p5+U2i1/8ItD8hrJd9GE552fXmVU8A5ptjIs1rYLm6A4uzTyDtg+U6qJIQwaxNcRovhnqNZBf
ZvKPHVB5MFdfWR4uw1Q4xLM1sXl4rww1wUBFNuylF108Vf5Vx6xyrhrWwhzs47qfys+NKI9UKoYb
Nf4SLPA8A5gvKZiXVfKWwBQhi/ly8qpvXRMXQfEFERyTYdpRbgDwO0hmOp2i63VpzT3YpCEoAbrO
pP+97JvFEGTqnymZN9ndwHrKLeObUUfl67E45qvDAXLzyDafLpaY8bGA/clGNJ2M7xBkT4591/3N
KQC55hVGIUMlcd097iTfbJ70fi7Fj/tPl0nX6t9UJfhWYgd81/1ZaQOOz+QA4amABVK/c4sp7Q4q
XwQgapjueGUAd1ikGB5AHTehAL725RP69AfZ9NDJXq0n9waW0ABUqHpeozSJUFj5fDTtULPKvMsv
bTytJdvtFCO9HKe0xr0SyzX4ZTsPkc7L4lXlAUbVe8g57E3I9/E49+7suWloKpDTnKLjRnNsf/ZK
1gnVZV+FY+IA/S6X0Ry3mgF4+eYzaMnv3jIYdG56q8RC6Lw6zR3lF2FqGe1ODvSvRs+AxN0ni7oo
9T9thsBUZsoKfvZxnUmCicRCMkwBWmyEunvWHLIUupFA0OtRL0/yq+kpX1/lUIUbscx8FQhjdvIn
gNOtqTHB5GRkCqFJI5fJBqEjbPmNwMgbnmC2Uo6Ewij0nJg0l0/X/MXTjXPyLrEnXMMZAR/xcIKn
qdY4FXvieCSHCSI0XMlQRVMNJZ/G5J0aigDPBEf0UK4t07T+tKySNHIGqmG4MVeUFAOieOEg1bPS
qWmlRT2DF8Uar/awI8SHY5FadPhKFs5V2ztCL7iqdj2NOQiiUyN0bf/sP6YTQVnHkT00/6Z2mCHO
IitlvdL6DQLpBjw7n3vJuO9xqW7mSiSAq7DZVohE2Ryex6//7aptRuGYrt0E63ZLiMKNTv4Vvins
soYAhuEUQk3yYRkVLf/GJEnVD4igKV04B10h5xs+MvPT2KLV9JL6pBAbwZoJTNocpoAGC0QMtF2e
jy3Zb31NY00n1z29Rsy+XPXLjyF4U2h2h61MIqV0sVl6KpyohvF9ivmjvmZBDYLZ0PquixD6sm9s
ZMGIHtUNRVGcNxdIxA7L8evENJzVSSPBX3UBAQQH3d5hUn58w5tOK5Nt6rPyICh4FsV2GDEkQwOi
L4cdlol8ApotJFeHtG3O00Iqbr06r/2bVOTTx7HWeWqDYQk+jAg/u7M/67zdgblT4irQz3NafvEC
88HgBoyndCw0zhlS3w0LrXThV7ZPL97YP805ld60UTLQkXVPILEnRj2hIQy30gYACzcWEizGJTYC
SpQbePej4Mzdijvhlcux2EXphh3tDVyEmqSaje4J5D6h1BnvcgNNxbpTKmE4zfOEf6sAHUoXp/P8
oKWvCiCeeIVNc4rhSlGCKLXZBZyQfem6m1I2omAXJZzGuvCKnPWNqQKhxM71aNpGkL+S3uj4LHPx
67E20fY+BsmoACLBF+Sm06V867Mj6JdHNicHcB2tq9cvvmFee0TTcQlC2l9UZhN4pcUSXrahwCX4
Kq28cARlS40/CoEbsozHeXIehg3+w/oy8upfPeb/kut4lRDmnRho6v/P0WrneJU3Mku4nqH6asfe
a9tJnZRChWWbWXBdyqs+V5UjCaGrxOS2uswawngufG3dQtHaV+szHw36t0Sig/RpF9LAh8E9qIIa
oHjTyp61FOe55fciduNOXhnHhkhcnrvpnCjuZX7rhuzh2MDRG7mr2S+1xgumXtwOXolYI6mCKLn2
yfsDx27SlLjIPCknjl61jeQddkrNH6cXcDwBYAF7XE03KZmlrYS1/tNw65x90ugwO3BDsf7oETLg
XcJsqFI0rgEdhaEHhsR7pKHNnDirbRAnmDQAftsYbv0Z7+plR3mHdmtHzs9VO/Zuecnp/jJXowOD
p1WPa20zsE/g4N+w+5mS7a4kvrftsCaclbr1KJ5HkLGQBLgyw5r16hYOxiPyDJxwBpyr9Z9MJriQ
cWc8bKiEeBPycpEgELbp1v2kd8HKQSl+LqDOIbVeysZDeOINg1LAOyU+iiZLST/2iDGVwmMvGf5b
hroX5DYpT6Ml6ULAbUzE5YAk+s1Nafh1CNYh3IYRAIBy7tJjeWhzSx2cI4ahV9E5bEWZsaH2O6lh
yljF0RlhRCmSa4bSrIVbhxLHIxCorOkU2rNyytQcgJAe4Pg8HRCaStz9FPDWHrlyy+ezxsoBsaPm
abigEdu69E+cZhbIbgIzvcg039XAv2L9ve5oWOJrcjYDborriXH5D9gEh7EaRtW7SAv+It0Nx5h9
VSwEWkJgg7SXVBMRotFuLnQgqgiOi8LNzPpZLdb7GSRpXJiuhbhrswDXlXMVhbVkUTh2cq2wqsLS
uwSCxiZow+XKWwYhVHAQd3rZYnnqXXy0lU4cxFhNe2RYAbhWXx5ykwI/QfsOjJss5ibGJJNQuUGC
wMINjBEWhnru2ZE9WQRZSFaE4uMX/xrQ0ygmmqU/ArzmwsRR5BRAaHNVzAPOSDYKcNsbpIww2Rma
wXlinaES5XBVl758nl+L+2hYIzufIh8GIwWDSjpDrvS0qntWK2w9NgDF1GVJP+2jZMe/1wijP/BJ
ul3G0oCDTfjwQbntpTAp4lpj2posqtTKavmagoiSZt0bP5rFtehynchZkL1zlJXVPDmq8tFlbPsW
P4WZwS4hQTfd7K6V8qe094wa+iWYE46hkAsNehxYD5SdVS1KD2Migk0sqhqEA2NovDIgDSRMP7Qz
e1dwzoHyOHMqsnINk0K55CJeb963sU5+eISX7kFAY6efLrTiw89LY2LuNcM8XDBMDfrwjxXKERnQ
C+YZrIZAkGHo81SWkha71hFmF0SI37TU1JQaVRMwcNi7vr0L++7HeIu9I3490oky8xY2A2k6qS3a
RSfzEQqzA5zdaZrV0dvj/s+eWEQPU5lTtMLLbyzjRtS4j9kmBAFd72WFryzXFVgvDkVYiJ5m98hG
qsJMW9vPwwupoON1fqZmL6VJGV35ikSiftaaxAv0SHeQhEeicwDHRL8I8aTSyxOV/BKOexIrcxIN
VYINf5P/Wr8E6zra4dTPq8w8aQvzxjCA1aU/FJllVeYJHnKJmg0XORUKa2vgPIhOZP5mJdJj/O5D
WHIy5JzJSkaLJUNbqGF6xlUaPv1aqcSxzfiyM+DSf4PEUtMmFD6qNCJbx12n/Zf5SpRlUStGsX+2
QjfTaXRTg+khHgS86LVq8osrcZDPavpkkbXKQPC1j91LL93QFZzxmEzyasCTpffr4RsdZ4eHUMw0
YdjPTrxO6xpbpq6LrGXiSmjuAPvYNrXfmeyllPtVyIgEtJWwe13pjzo0Vr/bG0aJLodf8wHqJBbI
flDUr+pGgqoeodg9htEaGFOA1W1WYwz3CY9nU+QeKFFhy6Xc1QyskCDfRX6xzDeLYwLPgz5wcq8I
UYRBTi3KFzPqkD3+ypBFhzEPZwtYm6dE8MtJa5MPsoUGBQ/3vYRUfIyVfF2pAz3tDpTTdBDKZJi1
7LhEErSSLG8f8O9AsJEPFbU+Hrrnr2F7EwtgHjp4vTrKWoXQPxIhSSY/nCaGOvrwCoQCwPeu0ty3
tBgCdg3oWL5Ct9eprG1TUr4J733JjV4AR9dY1nM/Zijn1EsM3wLos5WTRimra6wDwRgD0j4AGLZK
1HjclNbjOY64Ix3LjTvhNmAfVYkF0hciL9XsJgQnTSJLDxdqxHMIQoaR3Mk37WI2gPVW+YmSUkxS
Q1KD554UaxIlbRyg6ZZhqsL/JX6XY0Mu3JvfcH4LJWp0zhiKaphXCesDH2mhq/Sz46JUetD/8K+P
YcI7gy1r58d/uUjaKv9gipxpgiYaPG5rsdAKaysFbVopEuk+uHuNmQY3QREcfasl/CZCKCBgW6hJ
L0MKRbsQ+2yatCaysERt+JVUQswYvjbPeX5I/2c6Tswwqnb3uZVguWHoJ+BGxe2VXauoqum9vdaV
DH7DfdH6WXcElT2cAKFuBbgHZLXpKlYaIpZ6AQV0B6LnXJUuF06GP97Mq+KJLmIbSPxRmhgnzjIa
tE8+Ie83vTqcf2HkKEv+wR83IpveBh8CBrmLLw1yIwnX94/EvZS6VtlS4zvRqtmwrtI30s/aA91V
jo1f/dFqiPdJR/J9h7TSKe/FWkGYbueF56lLbroeaFElXPpQTECPqId7mPz3wqfchv09YKWu9DzY
6pCMvfZwTAom/2aZUzPz/YRJ2CLCWsqpmY1eH5NPVFSZjDlnCA40JiMVmoymIFj+AslR8RMMlzMg
HhVvGF3q8LrpxtyjQGHJ77YNwPVG7d1Axn/9CrdHixtMiPwMQ7IOP5136EAnQiKh9/IKR43eoSE7
PsMedT3kRaA9reYCgwWF5m/jebFvHZ5lIavP1e1A4znqQNDCIrY1kPQGDs7i9qscFBBHvRSqwCu8
QaU4rUuJ21UtX0CwiXJwIcSM3sTBp/XfGtw2M1jPgxekS5hwBA6v47qu6de0/QpT9QlJepFYL9n3
SNZJKE0qy+wEBx4ZkWucMKab4MYzo/EGqzTUxVVzULFkLL0L5ggzvyLWGcLZFFdzmO4MG5HUphYz
gwKmcCsHzCucJ6CQ+0s7tKz8JzIQ1B1fCEVoKxCGPCii2Mpqui9hOD0wulGVYXG6f2TR7hAzmB+x
a7toJY2vUim22Lt+yEdMofLDidqVNyLjJAUH7Jbjnz3EfDcnMUeATrzek1oxxn0393brwQ+xdPnE
eSizgPDXXp1MwQEMpQWsEBkcG9/fkefoQozd4y6aOptUuF5XlGdX06KhjkI1+ie1tXLRu3NzRSj9
KhPrmHN+UP8nJ5Firp8GOilLw3PPF+wK66n0m+o6mPsYtZrOtSU/iiCV1K5eufpdolXSnD/9e1KS
IXLgMHrmqyBdQlD54baT0G9N4xFoGqlEfUvaR4eJOsA09mGWH5OoG/xpNP1QHcNCTu+giRQOdB12
IrJBUNnTizNX9iYLChcNou8HT5PM09la129/fnDQIxO68CgGpCXeJzX69ppi89ZvmflOpEvssKhp
xG6EUkADnl86TLsvatHuQL5v460/33y7fygfHoyKepVE4ze39jRb/vS+JWI9alNrwf++csXGAS4u
O/wT6VvKPnPq88bsPu46sf2NU+C7nyphbqcom37VDda7yOmYnvdPBpG8AessJJbVsFsD/4Cg18XR
lJ7fM2tOytRMBDd/+OsKmbUL4CaquyjivZKwpj6cnsgF6Yhm18pMsyLSHqMc3Br89sOZnUuRb+nC
5cZQFXjYPXTJnCwjGiwscoEYXkMpUIXu45D3cvkywG+0fRI3bNqS9DbQS9aaS7uw44W+KZOK0t6V
aOX+8oPxPEUGEFRzPslfs5cDaE70rYABD3NO6MzepSuhy3Rn9evMQdp1vy5heDGetZ8wtfKVWWDV
VfZfUoJkrVwPHSUC8C+qU7KvKaA72Do63liu9jJwy6r7CnuZkIzIaCjwh/ft7Tbztr4Lhl2chLNt
3hMoW+m1pY7iWQkS4B7Si2asM2kr6K86XGptXdEXJW6QGDd1Ov9tnJ0EJpHDGkgpO8qAeGKg6tmi
TxgIsBEZqkg0z9kZpzwSJNOOzOKzPgGovUZxhbj41T8eaoPHJh/T9PNEn5XRGHpaTTZ7MxsNsFdT
+DaMaX7lDeSl7T6zI0d6KsgtSaPteRDgpcCZNhrEvGWhTG2PILDweOt8xTKOfmBjtf4YcVUhHdc5
4iuPwZvoHzyX/ujCJba4E/anDWa3raosygMsjgCiFMpgztmyNtJQ1fw3OBwyiPdxjJm6ShEG71s8
VDDngR4MkzfIhALbs4NRZC4BVtJYyCI05P/V04pPh4U5vcxRHXI2yRoouBOR61iu0mFY5kvea85M
cKBP/Pw+MEzLmU9mfh/E9iWjAaccstl4xwJxmrBsi8/uCY5CTnPG+nWuKxRMhksuzznOaeqEo0Ja
5RBuDQRnQF+0HtJb36LaSTRBPdoGkxVduRqXF0V9MwdfVc8q1E4hU3N40zfQXIkfclsnn/GnV5fc
CUnbDT/ZGzkIxUEZMZaU6bQ08IWCg6V+vouqGAgmANJp1s2Lbreq0aL2Gyif0WhBOn8N5wLTYfkr
dJZDfe1uHwH8gVG5PfjofRrRLwvN79M2Q/c4yGYD8hzN+NUfrqU4MXjKwhsvfuTOVbclVwUMHBhM
3j/BVBkx1nPE7TDAhSteJviS0mC3hQb5ENnqnn9JbwSIdUvlWluEjBEJakFok2dlRda831i/YcJ5
qKDmY36KEfBua8lWtJA3CwxfhNVG2r5KcseB92gOKyIDV8m8B8f0Z+sWgBhytin9Jld0XDpMfx/1
wWLSKe24oX4fKjcb7yPhSlj1wARzjNf6w1yGAC6Pe36GTLOOIVixFQbMYNo1aaCst5iHzVjR1qmF
B2sdYUQcXNsTyC/7THLec45ZFklRrkqh2j/BHoTqZZg4VyrvmZZJfIq89D74J7T4qmC03Wcu65Sm
PsjcWxt8uBniD7hNNE5Ku4enTB2UEgAbiGhsNzh7+x8gMiFd6CygLWkkwknj5kNmG2C3mrJCsQOz
Bx6kIBqnVwjtkELAePT+GrIOfRbjHhX8MHd8yXKE+cCySzTd9+pEEQSSU+ByV6Ca9NyiBx1USYk0
lwRMlYjFS+umJlliPHufZ229NuFejc+myEmouK1THwYjKjt+Ajo9gKp2iBLt1EaM9QLp1vLm4nOF
3Qp0GWdlX5wxuV9ki8CTncIqWlqNdxUAxu1whsOr+H8fPxeug/MjqNRSA78BdQRlDiMIiaPvhKZL
QGPgt8476bTb2VE/MQMQkQTGbBooZWqjTVZcgsyUqmZFCgQ/Xc9WJcvhszpbUTb+RyEeL4ga01Mu
28qshH2IWa+sSpQmrnpZgioEso4UoOzWGVpaIMLuLrL7Cx2YuEXkm6AN3dNSjiVJk3QqEy7xayWE
xqwQy5OJhJrrvfoGCS2SS8AhjXOTRITBdIq3tLUBdzIa2+Qs7lSB+0ZJxFT3H/dBzTl5uHhtZHM0
ooqe+TddDrH+QIkQShHTZ1Fc3S4p0Zfr4Z9ed1pe3pzKrCjl+nIrb20nuNTgjOLyF2Si+Cve4k/p
92xbx/6qsZCDOTIaSoKOReS3RiAEaRyhEweO+Zt+q1i+JKmzU/lH9Uo93faSKGRFhU47rlvJgEt0
H1wNxJA1wkWV1qgwOTPbCC7XSEIRCteEtMgNonVUtzsOoclZ92v6edtz29kkR+Ak82EFIVpnY/+e
h5okETvo8SKSWPr5AijRft8McuxyfhMMTCX0nkhWvxJ/2VNwuFX3OPeirpvEiu1QbCNurHx1LXub
lX4kJPwHVGIuTYUBquVxaOmq+rPfAGXJafHgYOmS9yA3PfQXZr/7EEawUbvYda66TJqzsOc//R/p
Npwv9q5RGMu3/K4Uv590SdngtW3X2FYQpfGO7F59cGlZ2eoLqbuSQM2WkNDHj00anPE+E5ItLStJ
6k23MvkdH5GvfrUmLn1lhmcOkbAbo+rLfC8+nRZqEKjA/6UGLJXrpijFo92GMz756I/gyYFs98lX
hiyeMnmk7vBiFAb0nsY0qEW9WJZ7vlGRVYatRAB/70Sh20cTZCCDUbKPXpxGOzKZbETP4B0SqMOL
cuaoqdSLJZ1RUNO9PvB2HuIrrSpmmwVOSR3HgYavt204juzS/yzZxc8iGt+bbRoof4VFUPk3F+vp
B9C7inZr1+RwsR2djXqT/UJdS8EjgCjzYDFU5sXdd5iGSEV5unwHMnQaqwZZCdXfRmqy+ONI6rQS
+g8ZU8YX4PsfxHblKzUHNAZ/4Te33bAy7h5/J40HTMBZBg9etEZSFSAToGDc8aSEh4JenOPDnu4H
fbnyp3Iyp97EK/pWkHBHDuvDsAGrhvfjqLtKLzTZzIn0Tuud9/fHy26YhOSL7ae0OIY4Dn2pfzzy
JsyT+0dtf2srudq6SOy2stgp4381R9YBegWyBehJp7iLFE4bGzO68wE5/vH0v4B6aeqRD9zbzUHh
USFsh60rvFoYH/8hO2Rx+Zc52lYqNcXsuGWICjZxMX6M8pI+bLpig7z+BJQyiVJCWPAhQgnZhLJB
QICju1JssyN9wXX6VJ0hVuFLycjp9369MJ9wajkY2mW1IXfIQlRdFHsA74kbrshH6539IbHZOqsH
HNu+GYcQwTzdqZPPpejxe8WMr29lJMIIezdLAGUG3yB8BInR0PXaNnsp4xjbZflUpmvz2a0aSZmS
3mFopZ+mV3odNlZ09RlEKNgmA+WXGzknjk1gv66zilpSJXkmnMEeNku2haB4GwUUeqER6n9FzPOf
L+7YfuAXb1q1W3QHTb9uGlyboEdqx70QCWV0yUvh9FLOaigzkcZuVffzjRTrStdGoWbAdbVUzWQt
k/CwjEh9o+AO8uZ5gMfdl0eiwVkLP5dW6SWsIpT5MDpoTj9f773jPLv0w7+Zt5X/VzWFcICOiD0b
nXYaHt+qD3BF2KBlZF3K7w/eSyEpYm1rjUVURHmI5WtMSIugHUxIMpqzfeCiTZTiP5zWfelAUVG6
MKErrOllsQ7OPHh9mKVNbbb5+iWPbgCh3KQQWe+mpiNqaoEfSVha3JkBYJjcLtmM3sqYLveWSAji
ap42Mdl2V2526XSFeNq0gzb9M6Z7wzxjeVx3qmOHkEKDgNuDIsDFqph/9YHvtGcingRiCZ81D4om
5R6LIxiS2lM4Ue2AvQMxHv9OsIsbVH/KkiCPUqW+FPPIz9coCUuL8+QBnEGKYIZHwpaKuiAh/EvC
1f64j0s8/ce9WxK6KwHR5K4u4oMmgwbh3lPfiOdIzQBG5VqBUeUJXM4dU4rxMFMf0R6/wE5J/Z0N
nYuNg+vdno2qdQtjdigPq1Ae/NXwUBLFMwDHOI5s+pvYCieDPiNpLnrc0jR5YvvB9JU0YgolD1jJ
AzZluUPw00EiPhFGyIZ0wHNcS65HvA0C+cJJ16zReC9uhMfAVdNWx0qV8I/+eEhPtiNmi5dUmgRB
577jSk9QvPPLjjiKIpjKFNGh7x/fnKcPwRhLX1ybNn1vRNoiTIXyq5sTu1GcGbLm9Qgfucf/3+Os
Lz99YwFBZ3JAP7Nm8FgLq2J78WZWn4XM+7I9GWh8lajEO4kR9Pvg9vrQtu/gT1IFG7XBrpAHew4P
QBRwSYsGSkX1INjuhTxSzjfkj0kZwhmsJO3lZknJFAT6LosIDQKdQB0fyHTpoNAYr4Bqt7zvWpc5
Rg0WW0vww2zIWzw+rKN1+192cNok3BP5ZPfYdZg4Z6k330ZVsxl5yyI0WmI6jkdROBakMX6R+m8s
NwxUYE6m0JcVPkLY6TNJy2uM1gCghNKjp4rj0sfo6tkBBkSFEGoX7a0UaV7MFNkxlz3ZmenexB1D
4qko6x+sU8HncjFGL7cFgC+WSxfnTlqmdW6nNdpXbEvvFYl02S/KE/OtvLxOEVjRQaCPZJSXNfeH
PQu1/hZf+L5AyjQLWxWl3TWP0+G9tncjAV2qAFcp4mBuwNTFCElztz3epm5Z/sH276sCGHTmeXBm
qvWKUJBTY0X86j+9LF/0YpyOfvJofxupY49WmwcY0q+N1SS5RoF4PxprJ6QFbLw18Et98w3FHKpE
s5eCGDdIW8q08DW7DT3cjwPJ8gyFECECfuuTuw42QFSeZTD8C7+rob4rUWxZMP5PlTjm8reqUFqo
MnlzYdb3Q0A2uJs3zT9j4M+0Nv8XUXvJakA+JjgmQsImYtkurQdvi5VaH20Qef9567tzwPngqyE2
JoC/sXMoI+YG4gm5Iu8QIXf8pDA1QlplKcF+vBXWpg0AikdD6P9mUokM8F/qg7O0zZ11O2QXGtVI
h7SjCrcnJDiTcZ+rdP4IhhgsNcPHqSgbr3j1HibZSA5pczCKZ/OeuMQ8663Q38Num0cMr7/RvJgR
BmGleH6a/+QU64Xgki6bI5F1ou9oYRAfteaHXGRfOuWSRu6WMyZB+Lp2T2Lj3MAh52WkBQDuikZ6
dbnVo6OAgloKA+goX7CefQW2KLtDMPl+rRY2aIefZkvp3rCR9mqqcJ2X4TrkxWAgKZNA8JUEaf0Z
dFr8ROy3VLJsw5x+FnlUL5wJBQLBsxyCXgbtb/XxLhPhzkcfvAJD2QM307t/xiP4f25WFawA6e1s
QjSC+aellaBvZXr+2xruRm6e7jjauZutb2WGW1puTmCQ6Cv8YEtuHxQuVuvgEDuUCLcuAmyuBzUx
2WyUMAvOdudyVNlW9fg/neMXdPsUuR+s6cTadLw/6SNwxRLiMJmRCTw/pJe6i0CXRQsIWJSpU+Of
+tfKT10LwRgpi02rpq1iBEQnmkbKXjlvv2rcQxhdFdamdSjfn52luWgCnxQIIGgfZaEia0tAVLW0
9+BuF7xTSrwiLZY9tDgueDTTqzTQoS++zMxjK6iUTIQA0SIxiJwMJ5dXK2+1Q9v0as2EmynRukR8
3WMlKrYQVgwIisH1FrUe6XtoTt1tCtE58eP0Hm7XqWZTd/J0Tb8XkIugbDlbB2EI+60XWjXGILyN
dDQ0xt+87Jhi+BImewB1xdr897Gwn+K0TnNtf+H6M7yO9rA3I4XEVzq3IbZBZudKDTbdRyGNpIfR
IJ4blzXqWe1/v14fXrGoYZhNk1Db9QZn5ydjA+0MI8nq2mds2Oe7J2aTlzXqPXXN2FOxm+owyFdr
m/j/sAsqq+OftVEf9AVMlDOWSS52YG3eBVT1/hHL33bIVBCeK5LqbAdZ5PXBQiaq5BqzGyItpk8E
pubDxJty9v6tk8NfauE04yhWRYJROQpPTvcOKRDanqUH2k2zQwH4SGL5OOqF6kuwVZrM2pJy3liD
iWKV1SdLNT64DRJ5XyFkVuwUT6s63BMqV+qUIxn8qZ/kWS1MdvKRyW78GAqLFRkwINm0uQBgUWfj
aFLZQGActEmhHy3r/wTu/d0vbEXpMH9qjWATkfG2nIqujLDF8VEQpeI33ceHPnbYKYHPixvCzD9B
93Wvmroj0cXCndjmSWSOlxKY26UODzv1WlyK3POSYfx7+vJHhfrNs97qT20DcC4oO/zFB3kDDmlJ
/nchtvyxOcBKwMyjMFNYMO9B0Pwwj3UJVrUXa9DaWaK5RgDQLSSXk30qEHbLji8cBYl8d0wL2ctB
khZfG4YGBfzeHtltykXtny+UN3cKCVndzn/aBt5u2/s5p6HPtsXtRPew170p8FOhC7HTMblJf2PY
Fh2CduMVTmMX0SsehsQTarHW9KfqEy3eXvS3JRMrosRcE34C9PtDWnqBdzwTmHtZoGq8caQyc1oU
hsbFyWR6fofSWu9KhM/Jrjaca2H+oAiAs+8rORA9yPXHZO/EICqE4+cDSCdR/SkHVSZrvP1pRVej
2Aw3TFryRubFNV4+TzYb7VF4ZmW7AFWHaGeTMARj6+MwQ7CjY+u0n2ZjVPhG9MqhPdnQTNFjYs8D
uH///o9dTJUxBfpLQ8au5K4C5OhLK0r9bcM5LFnQ7RY3lxf5Zz5Tbk45U/JKCFmmmSNYZDHuRnKs
nwcndq7NgFe7ggZgzMOCRbyNy7yOxAopuYPoCCu6Aj+BjrS0uxAdWDx40rFYtHlW5PWoIiFec2ii
+8mUU1vSp3rJBaVbaU+S/1ylUpWfnJYeE+tnMm6WuuId0XY0ggpvdNCcAwJdo/MCmxU3zrxtgbWF
uRlBXstCpFYXBlPRIuUswHNjcrWYZXhSYRScnKC8/dJkljmGLsdPn5fnZs6lLWNV/+gLp4autaOz
JuVshEDs1nPSBNWqMVmYMwRU1CJ5RJ73ZG1F11N3QmI4LUTo+BTWGutzb2s5SmxI7jiTifS+mIn7
ulcSy/AgTE24MeJZtpvxKH+eSKVHnwiMgGT/eeqU2qrLPqxWcJU4NSAiOGUEwlSiy7ZwNphkNcoL
u3SJF0bThardU+e+n1gbiEJB6tGlcmieQrD4H5d0MZXER5r6TR6yO0zFy0zxiFaZHJKVRyvq5BYf
a1gXoReJ38TQU1L05oCMAduBcqcAtguZHp7UTbWLUjTW3nntEhNyONJrvJ/tDr6595cdltTc8qIs
iwvcjNpSRBdQUvMBF9Sr5YuaP9BWqfSbKBqWuxbzY8ZGLWK1TehitxnzMj+Of0t7H6NrAtDDfKea
F256AeH9MwXjKuhxNaKH5vNoFAafDHQOR26LEdF6xOvQCfRrNGQDui/j90s4ON+CjOOhl8tWMKc3
EL4vJ9hrUHRsH6CGVev5nEP5y9oj53y3UG5gke/OMxad6ObdiU8BQfw8J2BW2AWB0XmQ8FEY1MBU
OwtLK4DYsgn6+57zEvhKA0sQlFRPB/DUzShbuGtgvQH0HHNrISvU5OHRzbGfK7ernz9nm32mdJUx
1NvBGnXOYdsgEOEfvx7ChObXeuXbXXor4+yBNz9cyi2UfUA+37x7qeFWVaZ8DRqazZ9Swe5CJsLF
QeoqufF6VaHPSOtPJa+azlc9alxyA44DUxBCvRsWFRdC0bTiBxFfu7B//amUarDd0Awj5574BRRq
J3qGlhJeGfVis6uIdNSEdJpDXriZpd9kN7lTH1/KG1oaV2SLeMP6AHnAsXKQMTMUWYupvRiX3OLF
QSpWyshBHKF7OzDO5eGu4m+379vZSVtHLsx059dV+XOVfpZuo5jhnCTIbERA7oVyiox+o6kx76KV
JZ55NXIZuqnwYUohJpIbX7wYCs68GZYKyHqgm2NvDMfQVXyWruuvwEXm2eJbgcC73i0EIHy4CbMd
qBSPeNoXVIHPED1naXI6JdBGLrWzf5Lq5yK0jxp58W1ueQe8J65rwXlLxW1G+6shzDEv/GWk8bHd
cAuQ03Gl2pQxbLesBwuU7I3jBlLOyOkkF3uuDOjRR4yY03C5s40Zf/Ofs3FAXEDunNIQpRuGXOCg
VEiCYlTOdIjkcK2REmbWzgpWoFdjtmbz57Auyc1zDDPGs618I+1ET9hvrnoDpDrryiqMhaHZ6ouP
+BVj0Me1OQjwrI+4ML11jQ7HbqojGYRAZJLFmgorjA3nxMrBKNPyI5NjQGiyXQ1UknGNmJxn6e+i
dOxugLBEobdsnt11GPjb+PrgSECdvDMoRjBcwRkNBq+yhepNn5XelnbyeO5dgiXpIAXKhrfxVWUp
jN4vkNV7ufqsxw7WL3L54LEb+sy6VZpAdBqgmayarCHPdFJOrKz8xHkIncbogGgDdsYRiYoLA3om
NG446XkiWo1RD5LATwL21GzPS5qgYRCvyfTogqmQQHqNNg62PIZseOQIfAG1cq88naiL9ybKddr7
Z2FiO6ttR+ztBjG+c3bYmDZ3kZdSa+aoas66J1dILyseCwiGZG0OHrYn754JMswscOtrhQyreFrG
6o3vIQ332Dumin6Hh7zWxUMSbecRmQQg59aP0vIP+82QZkatNtSj881G717l25Tkm4u/llsYZ9j9
JQoHlgrPiDfRWvuhCEkJJbzQUq9R4Z3B/RgIo9GEcbKigN58MsWVVcj2V4kWGkcrLgw2Ap/cqSIJ
Y9zZ7dwJxTDmzw/uAkPeSnvXxCJ2j7qGoft4u6ouXhuFJwME2mqhRpQeAdCf0IajbnfYjPPtQoJY
yjsvdhcWWPMf3L4uSA9M2HRiyIQIlLVJmX9K5awvrK9tcXvEVWlzSE22LtPrah852IsZhMqZfUaR
Ur0FkFEyFpczuvn01cYOfLdVpLscByiTqwAK8NCscbAk1Y4J2O5iD1CnRnrlpHhP1XRjOSbbG9hg
AJpPMjrubHrvJImHr+WBzsiWKYL60y8CxwjNLDlW4NA7apB32aXtCFeQmKifMy0KnNB6a7Eximaq
Ea0n13ybxXudfnFKr74nJvHRRWq6H84RRtgAWjNC2wFnB8Tus2fKUYC1mrjl5+bqiVY/8AedIXr4
dL07vbrRzLUJBqD6CuQbs6ceqcCY5u9U/h4ZiAMbPtXXkqKxK+T28iRs+67EiPZuz9Npp8IvdKhW
tux4GhU7xsKImucn1wmhm9Zgb6L7HUyGF14wM00s4UfhlUsQiYQrmCb7miC+PdR2HR0pLZWAmkm5
WYxXA3nGelOwVx9adrcxRA+4DVOxnyXBaBwnARSjFu+UprlKDpp1Aik3SM6n2qbfBQBM7FUoYUyb
hTnWMerJijPd2d8WqCuaHIfaeeohLwk8f2b8/fbaOlErwUUakE2NDjvScTBhn5GLw1ny3hvhTYFO
q7xSZWyA7jZ7xGjpQKOdP2FAJHtURk4QMpQxp2wPYGN2wR/XdyaqovUpnF4KAfB5CVfF6YwPyw9j
uikeHv5fJWg7w+c0ni888v9McVhPX9zzHSYSM4RHMrvzzwunUUkN/DjH9EAJYjxobasSNVNIEkX7
W2XYH5PyqHAvO6g+41wPau33aY1EKpjx3SLVEwWmKpF2Adpy+iLsZ9XAua+7mRKORC/q/kAJp2ct
hg7hkltnvsfTcKt2JHku0YZjnlI6aCEuOKaRwNaGKU5TlBGUmvyW6yaL/6FqPAAh8XJrB06C64un
kGVmdgtF30pWj6c0CC9adxTbkSWpVZWE1ynwfkIaSkcHwkUdfS10MJKWyurNqNoTHtZhidKCdGVk
ZgtJToWbE23o5U0RYFg6FIi4l6Krs1kbCuLPHXCiYNkirftm3pvfJiZHsM5OGlDGdrmNbBOr1555
5pL099EzgAMYPq563ptHc+3NfQalU12EoY+emomVpwEuOWDIczDp+sMOtV2qf6uv36EOzlaZ+lxe
YZwWoZZg3pN+6gNd5WVqhNkDgv+hrdcPpc38NvgwE29u5dk6Wo8UCx/cFKcTvRfuzPlt3YzlAJGl
0hflhFuKGlHWOiIJBsi3++oUf2uoAnT6vxmGr0DzW71lOQmBLioyt16siNwD4VVvsA797gY1FGeC
5Dhkwgu6PElWWM8/OkjpDR3FQ1Pshk4YWwqwsi7dXQ9PsOvcP4g2484l9zPCk8svNSMLCiX03vaE
9dk4uDSFkSL7pyDBl/Q2tkORWwOGXZySaS/hn6ccAX5bEVMOFWgtAXTWuNFaKFebYKk0er0p0gKM
/V99yye3+N+xu4iDk+dJYMbmyUkMQQ3KRyhbD1stRvzt+EzRZrGtWAZQ9ZJSqcTq12IDroHjA86k
AWNUHgXPPCmhV1Dg2mkPOakL5cO4OQ7HMHRcDmxtFWDQOHjnxooOvVLqjbqnuZCiKQVtcSP9spM3
NUnyPC1uFAdzDeHY6SnAE6lEWU6SNo61CughofS2GfHJ8doTjfSDY0Jd6KGosGwao77xVYEYlNGR
mDA/v/plqkzW7n8MxTYZsxQWP/VH7KqMFJZTTIi6cmfoQrsnwqlb/8Nrgy3Z3W6d00VL0LPIrKFh
yEvzKIyEi+CPWFo8lIyvsIH7u5eXlFMiQdkSa/L8VMVC8HSbkITUngl8Y+Sa9XWhnIX/XKjPKqNF
eUpIZhqyE1oUYZhzXH9N4muabIyGEXRMQBFyRvzmtO9ty6LYKeOvD7dXvAc7coML7ARj6J9D1OV0
2PP1onGp4PnTymfAItPC8vLbEVt5e25dijo+roUo/RbMw74nI4QH19/QYQLkwWeA5RQVvYN3t6L/
tP4IL4lCL91FivjWPuAtW3jcEJSq0fPtSEcPBDsGAtCB2Fnwayg/XnFNUgau1Ap/slGwesbbjHxz
nUt+YJiXvAMkrcTrSLXTgb4VfKTbdkGfp3tdelMNuc7rfF3AN4mL9uq6bP+MI6JkuxbY0dpvlSNL
7NqSzFGBfLTLWPh9WcmrVzOgLtpQ6bU+9wHgXEamHrNLXQ1LnrTm+JYRRFLDmOW656tP8UAVwDYD
g9mWxOs0VvBbd9eF4OTAdFjxWvuk3BsgRe+0bx7nUD/ccllKjM94KSH2yAkFq8mRg+t5ESW/e9Sa
O5QriKO1zpIOEsiSjyizdcE+IeQ9nLa2Q/sgxVSM9nZ1h19Gk4TtQUgWo7be/PE9ND+7g3po/JBh
mRHyl996DFLefdYDP/pF4HF4iVJt5Ry0u646/Xwkz3j7OwbQzQPywsroQW0TtiAFVC0V/XAvtV1a
GMXWHwA5Wg8PWCv/fPyxw+P5HmEfW4jQuUfukfwGOAzRU3k4PeSiqlSkoQx6mnxBp/pPuKML07iE
XzuXYF/yDCRP0MDeih2GzsonnTWfhLxW6ijKpMNF+C+DroSlwqFwRP//LFHNFDlR7VY7FTje1r7z
vyykOZyg6OVgr96jxJO1KE4N24pdozUh53ZDqOdZwDudGUyJkyCd/RhrSnts+/spCBULdkMvV3kc
UPDkVyhaqTdeQJztRBQ4G2l3gezSVpWJQImcWXN/KyKBqGxaCjEM++wk+fLngCafv8IINKCLDXqd
mwjgtBn5Fb/W3uOAoiq6v1r48FSo3Hm8zuK274A4MikauZaGeKBfMMIf2uF8j9sbgIhBJ5CqxRtX
ONM/IphQlhDfvj/Pq453x+elgysOq1RPAUH3XJiVsAT9T4cCT//1yG97bh5ebgEP7jJwV7gZNc97
ANtZmnBLYyj0DIZDTH3Xg9SBPbc0sDELANeSy7ga6iLTZSi9MMsxsESlTGS4kZSnRixCiXZO/7Sk
eDDWh/tXuwu6ZMT81YY0DiVt7deem7SI4HzY69ll+J86APPdEeuJpf6YYgYiVgTK2+4ztUgWPP+R
Jzo3Qb4d9llUE7eu/EjFU4n1+aBBzN/X8OnV32Xiiz4EndIApXV77UQN6w9QXEuRgyB7yuusjP9h
In1tTzuyaivYkQ1kNgnHuVfji94h7lCj7GFd/REvBw0IOEO963BeacqfVGyD5U0s8sHqSQo4ca47
wbXlTkPlSxhPPzRsqguFNVXDkxiN+m/6dZUQNC33LS9JpJTXyaFDKZ25XczIZ6fp0mlqd3r7R/aY
eZX/dHqZlEGyfKk1PvQUohn41Bx7P3SB9zg08wYwuGr9EDYaWukqNwUS14eiyO3UJsY1361QzH/S
Dd7msGbcLM6WsZ6wiR9VtCiq0n0hV992dZ6glB1mU/YnHxtLzltXnfJgQDNN19Y8dveh0qGaPgPI
6JIL0Q3OkWnnpDsmbDbaPO39WD7Q6FD5097DAihxYEUuZdud81bopXK0A1Mpm8Fcoc4EYIJ8pUGP
BKyt85sUap0ddaUppQwKjOcPqWrKyJm1X8wMaEch8NyNaEIDl4FYS3k8e/p4r94TbgPHZckaBT8J
6HoECz+Pipyp+on7o8hG9XGa47+kN/Byu9/jyRu6ThirTSjAtwIzL8lS91lOjbFExYBzpON4n1I9
/XxF2OZBY8VInPfVwh2B2Gc0ovRq2ApgikprO3p9xS66SwTrvd5gLhfpVYWPytYUvZtlC+7K1A/2
jRTjWpStP4nEOyD9ST6NPo1lE/KEeKzNqzVt1e4boNzuZREY9zLXODsgsL4lCn6QaApAUDf267FL
qI41xu34MKDlxuisux5xChFcLs0MXUFTDEVuXJeyKbwOOJ2mWGToKtfXKchG2hVbAExj9am/EM+D
sj7pbezuvMptYvD+0P/ka2Qi6CdQnVSOrWnm/ex+4pm5FxlrqbigFoqFD79DdlzVjz4OsAok7Y1u
QAaMx3+BgClayBclo5/RGd/Wh19T0sCSIG2hV/83ZYyC00bIBKjvOpplVvuXqpcbR4gdqUklzXZi
TeWQmWjg5R7QBcRLGRuL8mOtbqeLQoNCqGO1N37579F05VB7+WwJ8uwyxXYGYRf6c2n8pM1ixoIc
Iiz8JaxmcPfrQ9GyyNSgaOhGnlmsI/ZLFR2jOlYrBZUaHsxop2a9JFjvRXfTUnSXWxG/xLIoKg5l
1wJHMVXiFY8UMpYTnfrxFUCbcqORZ2NCbMchjux7JHuhMMXUGz90bEc1h0i0+m++shx8VEKZE2Ws
sLbkOd5eC9/2i/yrAJWQkfTrgxT2xe+UDgIVzlQZVK7CO02NgY+yEo7QDXhoGF/mE503g++OKQ1f
NA+1/2n/qrwKFv6E8aK++usHSM7pZzCEX8Bnl2uZh/aJUtgvzyLLsRRWDCWO95DYcexNWbor64Tf
44LuuxxR65rfQkkUBRjsQEfWhgVCrMkCFJ68OWckGzT95Dgadh/LZyelktm8eP8bRoUUsB+95Hh8
dFMKzoXUgTbaTyPyxBvCPcInu52VktMCm33ju8763SXBmqj8cvt/Nn3liwblRuywOr/BupTRAQhv
vvBJaKscfMC32dcfK1F0m1AKkjpXM294BlevmMGTnjV1fTzW5BFN0PowJwZRKJIj9xJHFTYiGosA
EnrxSxwowaMoBIiWlN9a5S1LvzR8kzUbva0E+RYTQij9BgiAsiaoOPT054CSG9yTX1hd2hNfIm+T
O8ybHn4w833fQj1/IAsdZFV3YvZ/igJqfJdDFzISTZBV7XtbF4ADhKlMwS+WtCe/ttK+YWOZ6v55
qdRNSTLY7smB8NcjaiDOMd9JX/CaHAkoy8RCU8X4h3UA9YcZZlt5WNNtiRpS71B6SEgNAqtEeP7T
zY+JczVV2wquqL09nJnTlsHCd71+0EatjvS7A5EyTkR3obIe1o9FkRVfHpx+Srlm7xVwjFyVLZ49
XLOOWTjxG6URDBlmcV4sPZ4DPTEjxmHFgEKukn+fTKlgvaDhtHUUPaCKkDoCY7RR8oZdt9YhRBch
8wddyjBFycoAYuLwqRBhQ0S7/w3wqEW9mN82pMcbD0jDlMhZ7RxYVLE1Oc2cy5aBqMAO5AYwxTml
KtY66cDwZrvBkh1n6/sheMTpbEStrauR5CUpXxe+RSiE2QieKjCUi4uP6xSItKHWzJ3B27AO0mLK
MQ9achTXSocXZp5/zLpKEL5PpDNW5YdmD2tVfcY1CTe/gV2Jm3FJ0E2QN8KEcT0BlxT3aiHn0cHm
Mc/rsfiN5Z2g5wuXRuZVGTat0kJZ3WcwlK9hGFiv49bKsoerTwcAFWS+2K58QfH6CQrPEdU1Juex
yblwBD9NbnUoR14eVTwQ9FG2uIuROYSxFsqAgi4rl+7s+pZIfYKaZnLA3A+PovHwqOk6NQpkN1fj
tcisAnxw9759hBzqkSw2/0D4NjmFj9VXINtqcDu8kOGRBhS/TToB2Hr3jNCRLnA+UlWw81Wvldc4
2QJQGkJ3C/QAacP8wHrKC4/jlsI9cdC/+ZFHL4pgZyBTtA+XAzj1T2t/L3lRZN2FqQHVK0ikMKu8
CeH7o11hSxx7oWCV6BBvprCZU7+PShp4g3SVeq3EodPF33OzVIgU97x0O9/KFPw3MBzp9x0nRAur
EZhYKRjaLBOCXGdXGyhL8aWpVVgLnj6hG1rkJDL+14cc/NOwLLHwzu3nrqa/DXuRfRxx6WsUdaR6
TCOGOqCdvEs+VNInroyZHGhNdQvYGnOKeFv0zv0KjgQVsFlH4TXbO8Lvu95+IriZnvSrY2yjS6NX
Ohtxzs+IWjmxyg4mNC7IJuWY6TqiTt1tTu7ll9MQchk0ZRxh/WBiMZgObGZJ8YxK33+xFCNjas5v
8ehuqF54yXzwRnpT1hmQGSGj3UBAVY3SPTMbOOa7E8b1CIPJUcgZeycAPuf7KHu/VYR2vfXiCRwG
jRW3EsOZx8/p2y6UPOgVA6jfD7xTQB3mn/qb8mwiLw6Q/vnHtBoKz5KHLW5VXcPQXKC6qIkbORkZ
yMf5MgWgO/xWl/160hB6/CHl+8eMff9Um5FFZp+acNRll0aakSKygbT1mXKRHPR/X4jTZAohniN8
RwRCiVO/TlBz0qIDZBPGB992Ce2PY7eCiLgSbYpnt2akcSf49p9uJ3xsA9elncqpx0YhFbNMh3j6
mG0oZpL3R/zVao95Hi2aPb+ymUjZYVLp55xM92nEjtuhtr0Qjfzv/3x7i7mBBxo6ujDRxFqVcn/L
6WmcyQFaUKGH7tSEZ34kTWGI5asgmqwr7rtZd4nKNMCY499DFD60/3s0hX+hfsH92iuaAlVQ+be3
JgrXUbLEu5da/AAoSK1yeHRb1xGTud1KAJYa7VcG30Z624BtrNJ2BwAuDIFC8que0459ga4VX110
uHobBihQBY/0UvZT0tU39R8Tl+mJVdL6sey4hG9qM+eS0rtAZsoYsg9Hcs1yugpvmMwu5TwhMiFi
zZ42jQurQwGTIN0O2g9rLXUBsE0MTlgmWduhCbJnTg5lQDWdWapK3p38D+4/W88Of7kCyqex3j0u
XWkKDPGTQdl45mVyLo6xTFnY51seEWFxSZACbZpSPDW3G8qTYqGaEFGOxbkO69E1xfGd8yx5IAgx
jiik5QsazfkdWAgL5Fei0uQhtKTYSloqVX/ihps9s0b8gA1RUZA8jXgndn7EPq5mtvLl9WixQTmC
QGR/vfJrQQgzCs2KmB5oxicyLiKd9FaEDi5V7VRm5qZp3JrBjomr2dsSFk1ymX+7at84NGTqXpZ1
o+12YJ5vksrpYt4ajqngvS9VY1BhbDUw51OKGO2RD8Y1Lj/bTYOnaaUVsbh7UZCh0GhTc/ZWo9e0
8QVYN2BBYSVm4YSuWdGacsaL+zyq5j1r50MFtExYx+h3kAjP9uPvjmguhFCAQbRCamrMELvRosk4
al+1FrUOpojIiH6kH8wgyzOUkP6eyCnGLUIUB1HzpSRowCsRcnNEJl3o1bY2nL2vs7hpPd7kW01Y
xxPla2wKRdM0QfeVtkV5VwlCImSJdexLYn8oeH2yXsjQtJiJF27XrbohJHcvqjhR5BQ07UnHRu9x
F0vFCLNPzy4th5TvCvOtnPyl6x3oKWgezQeT+YuzRUUgKj67PpRmhvRRh1Vf8HeKQDHcSkB0Kx1R
QdVTqBd+W7SF1pZi8bfb7GLVCUI5Ctx+ozzf5mYBavSQJXFljJyuWiAUZY3jFR7+DEdkhcA0ZbLr
4ooh/GmxGtXIvE+l+ugGT2OkONtngFTPwkukaZZlmw47vzeXQGo5+ktuGtJzHn5LIP0e+XoVlRiF
hQ3qZymUnBbxzzcbidxxvXxyNkMnw/gJ4PbZ4xJEjOM0AMN/AEpj9MboJREleYSjVDr5vuHBMgro
B2t5O0A58plFNnnc8ta0pZ5VDZ0lL9CFSONtVgoWeOBagkjewgvzIe+ND4a9V8rq0gIl1GH5mNXC
i6o2ZZP89zVAgctxkKyxeZx+XsigZdQr/axnfH2NSuL8kMt7RsgVPwzbDICQWWt/ok4Q3b9fsqXu
kYwii8IS9w6xYwmxaLqzeslKVJsNPjEcNjP3g9f0CpGWFlz3AEd3iYc2vTYLpABLJeGeJRLmqfFC
wnPMn/C4AtRGEqNra2tHG/0U1R0WZ8tJMPQ+PsfcaSjb02NJgiKtX8Wp0ltKSAqkyTyOepKJ93Rn
Zyg5+N964ZcjEK518uWzJVsi4lbU/EkD65gPc/22tHl2W268IvyEnFipEZokZtrJKt2c5jSfpPgj
rKGGOy6nV/Gq54qebPJMlTXjvj/aCSXvB8hcRRgOv3RLpSqeULUyc1WcqfTi5V1UYJ21zoV1urJq
vUuojTFY6GHmfJ+RRJJlDNhw35SGjkYkaEW+A7wMzEa9ynW7DhsNajFOUYkGnyzOZiwI6yh7X8vl
NFl4oLJ96dAWs82Q/WyG9ZSomzfTsXvVaEAUBlIrzsMQrVQjwFXPnVZR002DJRjTq4Nj8BCE2P/E
aLf6YNd1pobye8wzrxO8nxFgaqhRpOS0SX03pUH8Pr3SlaOpR9C686ROhb1WMb0Hsw8Xme6bmdMw
WJgdUuGNTFBLso3TxN1pznm7R7Qyn7u7Oeuy6qGisx7f9OiN4yTY2Nm9XFhRDo2zLsbz6mwmyuGJ
rN8BrYZsDzEEHi2WizxF/8e7QJf2WgmP8M8fncl1wOLqT91d5GEsCPFRl6HZuQ2kzpiQK0VoMvbc
eiQyvpj1YeQ/1HzhQRzyFbeUJkQ3pC6xCqwbu+KPapOq4MVpfILMCGvc+ewAyc2w29UfibtTYjDe
jhr+xzu6vlrgvYoqbT7f5LZZG8MjdLUT8vcFIsIU7iENleStTB/3lY+NO/QlbBB0vkJsQuHIaP09
3SXMop4oprY8erPOxST3vLQURIov75OqeJtBZwWwgzlJVG9zIFTRgu4XmBI1384Q9f22EkLPrD2B
FHvs3w2GM9l45aVJxfyVmrd8sTEpKX+QEx+/s8UOKsm0312SVLxF4Ghu+s4f4JZa0IQRx9ZQj1wr
N6H0YvChJKFaffvvuci4xrCoaQ+aPIXPfl9W3J2GMWiXdq1AyNt+/PT2pwJ9iqupr+RGx9Oa4d8V
nphrhWl/9Fc1rFcWH25aUMrb2ehSR+PViVIGh79680esNYT8l+A9z/vFLjBNercoBWHLqSLp2xJr
FdZMALsn9KPGyMFD/f9GumBO4Vi+jIzru7dcpMj2Clcwuo5ntIxu7TNUMITcw3+3IFzdRAC5K2ww
guYRsOj1eF4lRuLQ85D8amPYm5rfcFzbGGmOyxfMYHaevoJ/cC5j52M/bisW9vH+V6EsDwLs/y+J
C4zGhBZBlHbmyNNs2tjIZuIiLG/mipLC4iXqLHHsBqeaSzayp0o+JERUsUIZKyRa2Rj6S7F+Ynx2
DQGlL+IhK8krsa6NUyEA1cYBx9s8wx/Nu0F+f7kPSic54UYax0RZauWuFOmzNDn0lv3wGO6Nkv6s
NcuoP0dN8wOTqSDlYE8k3zBF0L6o/lPaJ0qklMC1b33J3uBO4V0rDiX722z4jrkrWa0BsaT4/J7/
zqGVmd4H3EdUIOyJtK5r7z/3z9OSE71ehacliSOWqaV4f/QJjt7wt6jzED8hIfzFI/WMifhz2VrE
piqVDC+XzEiuzIzcTW5oTr/Eda6lQty1z2qlganxYwgORRTNVXvhoCENHWvjkQz9HnnjZ3blJ7Ip
YIeEg0WD1SLrqLKV4ouIOcpouPCFZgG81XBaDn8Lp1FGFpsLca9eOIqfy9XgxzYhhvZhSDMl9iB0
UlTE9pnBvRhluTL3dq70J3L2TL0BpmmNWAHy0P31bpy37xpabcgcVTmEMEmnBQJXJn3qjb/n1Dgc
MbxS1MfV2tQT8o1QPJXl5HhmuIvMa1MLp67CpnC3fxpXvfr0rG8/VMFo2nLYxQCYyA5iQFuXTMnM
NodwW2BTpgUYq+6e4QrRCKNU55OqjArRIHsqS7NDjIW/BocP57hYPp4xvD/kB0zKmt9RyoC80Vp/
E7/4Pq+4Sm+03dVNlqhwlGB3LZHZBzpaXmbb5MNq4FXdpquBLAYMxipGIBYHniDpspgQhamXpuyN
KwY0I6mmfbFx1pekGFXdGXbWuTXbCTP8uZGJ7tRx5AFo4aPk4R0260IiFjI+0Ld8/StEHrFsioM4
N5OtvWG3uuju+dl9GlyOlS5WJm25NxQWYTXOGBwUDESJzPMePkg/L0/hvvxzW3GrR9IWC+KawujL
i32rtZcrvQyI436ZqWclGRNUAgbk1KFqNfIdS/W7uiS0IiWw4mkShIcTqG+Q7yRk50fz6NG4CHUi
NZIdqjpVovTvs3HUm6YGny8CJoI7qm9GOGgKQWfnm51tQElccohnuaacjf9On2mD8Q+jdICj5O1t
BByCGoCvEUCp/2RfBYdZaKUc6McpdFgLgDOlr1L9GTVzHTkSdZoQHUZfotfhg3aedEbd+z2jCD1O
2bQIA9ujbzsoQ/PL9FBNrXFAkO/0nSfYcy4dMz6KnNYAZs4wYwl1z9iyfm8PeddThK3lziYXkio4
EOk7EXbffDxG6ZWOUJkl6NewcAihwBWJd+SYteWiA4IXQbYsCh/Uyagj/UgTKLQ8TrItCPGq47Ua
jSnb2IeXjDIHj3cTaFgLcqvMHuNc5209BamZzy4iOZG1QQ3ho5rmJaeCleqZMXgj6ZCUrnEbi/ZE
s7L/gDLQtTVY+rKfEzpi6PmMsreOgszSBDopd/Gsxi5OUQFm4QiXH0+mRj3FiIa/Pc6OVroEh+sc
L+zcI4vNUYWSXhCQeKc40dMITrZFieyZF+69O0foqprgDNiDYsTSWI0RdV6NFhkkKAge42FYHsRW
iYTdFVpjNjIPXmQoGUE34q10/0zMLsw/kO2P5vt/lCeaJz2JyIL0dj8ZURYygDYhcRwhk1DUB+8m
nXJx3QDyGAz/FFv9t/5XM+chgdm5r7cVZJTFGr6pQjzwkMoqw0p0FMxgfrDPsvwlgMKNT9Y7Oh2+
iget7hmNFiY8mSwrKTjrxmjae9naQgun5wfNK5+wh3f7vjSYpm0NbKNERtAIgetjbyNMyySW8EQM
gqpChRwymq86zXtKC+xjJdthA2NbGTH8OQBl+UlGdoqX4PZpHCzrpaMO2yiFuLg0U5yOMrJtQr2I
b0AmqvCUMjlHP2pSwLhVxL/1Lbuf6bhanJgZhBtE1Ims9tXRIbsL+DXYtXnDIEaLsifeauTDu6mT
VVQmfcTyQY3j/LBMsQ7xza2xEM6ZcY6/1DH2Ly4O1mY2RuQ3XjeUEWimj1kSkV+F2rVHfTzDNnCs
R8hH1AHVWNNJ/2/qu0OksvZbfKeokgu0NZEXN/F/POIUS2Hn9FtLE1nzpc9xki0iCUVt0wuzFjKl
PySD3e3F8Q0QceKUoQAmCPg0MMTnKpFUN1MYWK2Dlqkp98Jyl+MGNc6CvW5/vWlDxZ+Tr75b09PW
A3fMDFaeos/2OnXvZlD5eCBits6mfrUJiuQ96/M3fLdLc7bvyQtuqfkgI/H/EdGKVqf2lzHBHgAK
SRQHF7Qz6p4e+UGBOXn6JB+KoDQdjsiU4wBkVRlzMBN5KB8B+P/aX2Ze6sUe7Wgs9Hv++qWoz0/7
Nc8HZ50NmIIpfjQlxItbSr/b9zrnaPx0PZ4lfasDw8tqqe+82OCh0necmF9ZYRVN344nVC+P2uEM
WKw5McLAAy23BIbc9y0/5u2m4NPG0tKaXj2D/RCfn+OcIW7t7lVty5HxB7h/lmPiXnBYOzCJgZYP
7aIdHy649SeM1ZzP9meFUzQ7tZVgdYexS0K6cNfQznXm0Kxlbxiy9tBcIGWK2NhpMFCRDA67bqPl
ZC8Yyh9W/iw8ZzwvhCO42gvnEeaoQW9RrRB6EbnJX6i48b8vcEOSp7+B3D2ZhfIRwKwZ/iRmCE0f
Mhg047UF9dmCpC2miu00U0dWjLKVuz+oNlhFRZaL22l1bgVu86oeyPE7U+gqpN2GuZw9slrnYMqc
tbGoevAriEihZtHItAe8pJKIUWZ/np4B7KS9hb4SGvePZQhyXrhj8fRR2Oo1/LLDpMjOa31pZZiY
XFNAR45wpiJmOoF1XtATpRSDSt/nGpQnm6izx0n8HOPSsU/ZgU/6h533TQDqwlMiUZo69NhVja63
wPgWSVH8awlvGXYML361z8+wrXE89anMI/3P7Qr9+rnjuerPspa/uG74IUcL7rV5Wb+hBQQnIqfx
v05ca4lyWxyS0nqXzANyHM25O5L8NNb5F0foG1j+XRHWlThVkaB5H7Sb4tOImIAtCFt3Bu1md3by
E7GQ31FpwhOf876bRdDANjPw6EJjWBMnBGWh80+d2h6UQgak1ETUCDMlpQ6dr9eu4L11JEBNoECd
ImcFUFcUMvyiWsNFUWZUXC0Xng2oGndrBZYxX+MpYdx/I1jVJjW7qyi5PxZfuafd2hmuVyxr2Z2n
VVwHHzgyzHyeIs5yfN/tQ36/EXRSBxE6bA3lpcQ9ENhn56MAZDW3BVoCnxv0SYhg6tSJxyj2BaMp
gAG+PAL9xQrAJXvkjTvP/gsWG/J7NMFsiK8XIzIKWwhdtI7v63z6UhGp8cNP50ACRIeI7uduRZCu
T1BAsbvaX/0raL0K3dBt9B3hBaOiKUmvbJoDkGMPKXb7Mw5YGxTs82AqBK6P8x6SFpxwEvCljBTR
lJPzAoDWrroByaWYNQp+Qk3LkXm+O+5Bf2X6FkweQF09ugeZbL14OsyYLik/5ef33BLpypcUl92B
X0624d9TnuxsL5gXthqMIUXybmm38TGJRz7t0OvNK7tZXxW4kCv+PIsFOw9tc9UIxEBGbJ9vS/OU
dWHy7h6DADWsVmIip0kj/jj/4h6yDQ00kRqiFRmmYLDkFTYSTM34TLLn3fP9QbbkqLWA12NgrPyP
KGtdj5lp9/++rK3/+DvINfmqfgpvhsbeEQbOAl0eusGk0Ql84jP/TlUmhDWRy9WGR21tuCNZ/nK6
qx4RJimtyDnf5tBlWnUD6rNLg2EObCQ6VRHUq/65U/blkUKT2vyhlByioxI1uFEcay17OOVlThit
kVnwpwGGXYkYDHtHuCKrHUVMgcBlzDfQCfjozmO8RDbvr90/v67aYtAj0WeqUEkyxR3Kb+lfaU7k
0GgrVzMBJ1ImffXtJzkHpwtj8yQgI6DKAcS3HeT9+zprP53YhcEUY+E0MoZ4dLqs28ZKohkM3pK+
bSIEQ6OaMcpHnM/FnulHXYxeTjwlYPYW869t6/zEyD+FDJtF4IbgfMlFq8wy/2a72P5vmv0f7Tjx
TjPUfzscAm+IizCYJolBbUB48eWwsFSfDnlw7zbrWkRZ4jGoF1n4OhCmy1jO89CfccdhlHUKTBmt
1VmPMhx9aUT7lQpmYrqhWmguut8TReOOw7zvjcUYspFWtA3spWTU0c/udDRROGagjjZbwmvPpcm3
25n9ecNjn1jEsxBJU01Qcb3sV5AQiCdlgQtpjg2uYo6l8EcTsRV9u8vKH5TmXajTRx5PkpZbqckr
DFIvhGwoI7W0r4MEKFyLpUL/dE0klOvm5QaVyNBYamvmWR6dy/JOXHZ35cUpq56BZaeoLWly3hdf
XYKMBGu+gSVC90zywHzG9NRkgYpexX4zRNwdnTqUZnq9I2CwxMO6GIy00E/beoOg+cttBZcOcJOj
Ecuy1Gs41+Bj3nx2RsgtRZqE0FEeILmYpQinVWL2XoXnHOlBkm02x45VqdQG03DhRHgxWcO9ombd
Rerw5k3n4i2EZocHIShUKxaZ985qXc3bwb/U9Ps/wX0Oz+VSeI7xZU0fjUz0NL09HOqMXgLWutgE
H3QwLrAe02IEoFbY12Y/38LoXlNQcMDGWhNgLRxnm86pvw9o9rrNP/bA9314aDcs+UDNgxgZ3tHb
UO4LIbGiAiB1xfV4pHSw45BiL486vNDTDI0TqdkdT2yT78XsD0liyeII6wrNH4hrJf9TRfqCYj6/
HzC05efXv5BvFih2XTVXrNECzIFs6v2X/aN845Eycw+02UF+aHpbmxi8Gpbxoc+DSIP7BXVzZTGd
04fy/mzoHKuhlYVINM7eu9XNAEiPhBczHnYIeBhra8lI8I6urqiHoXYWMejTbBIT0jjwq0ucReQ4
kKk/5xyC9bOFmyTZSYMB8yC0KzclurvhjV7uZtjqADPxmwzOnnO1TdOP+lVKcuLZsXlHT1cl3Ssz
3oJ7Jjd1sH+wkqVq6avuh6PMhLQadB2W9V2eE4dnLrAUE9pC/IIfIjiDb6ZfyU5VknlwiLOAj2eH
LcuQhHCNZ8FsUu1k6rsoPdYJ63eD80EaiyxrNs6VsRMicIG+i3ZtCiHnM8PH90FFdXFp5E83U1Bt
13FMjD9st3hjZWSmhRou2R2ZZIqTPF6ZXyCmfKIQsKjZSfuWTzIN778aZl/XWxLYAq1B4R1eeYLz
eYzt7AgqrsgdRcaq1nGCE+tLz7p+Qz0W+GA54MRfHJ9Y/sMokH/fa6hd4VO/ZFmnttkOku2fVyuf
JXcFw9ZPdVnV3t6TtWs2Nxaw5VwzYGqc3yd4UQ71kQkdYBryITl7R8Qh4DqE3zs/8wz7lJ56mtJY
SoKH9DzmMyWe2Kb2izePKZAJtIQRtpJ+8piSn2Eq92cF4wHlrMif0dzPXxNrPaWOs/mH5r2B/CWa
xVkRB4xcmW/aic4Js3J42nu9ToBnZt2VfytrDsuvVyL1AXlCC4dYoDMAQAUkLwKENhUqWxcJ1tFK
zP16M6v2S1prKH182g5qvX7VT7NFLCLqm6wyEzsnsUpbQ+KCnNBN8jTOR+I8Uw9quUFjEhN2Qj0P
mIEsdj8+d1delkDAqmLfOaEOMy6sjHyijP7sG5PaGeHnwIjqQlt4beR5uIQAeiQZj4joyl6hicRV
mfg0+3BVpGYba2PlrFAKO9F+7X54QuMUJyKTNum6zL3emk7+uvVoe1Ec9+c/0nYRmvRHWELz+33t
H+2HH6B3hoo2XICmSOFWR0IDtrn8n5bTi0qSogtlax7mVOa2l9TKIKoggTjDZ9fWPprRS3+o+eDr
2FtSQuVYf88OhbdlmyBAloBd+cCojz8EeTzYjmRoDxpJO+J63ld4+W/A2YqE0DCxEr6P1li5VGAP
4C99vQ7ihWAyMReDJ+6dzj8ZPHcExGYb3mFGiqMstQPaSwcrDPHHHgM4iAVQWqJvvKgKUmoT5N6S
jDgF3WaItIsGT0IW08thEc5ZuSvO3hVzDXUtUUo3I2ng2FfXzT4K3vOddJh1dBEJGzdw8qb/lHzv
plwChI2GhCuC3LGqTDSHlxIObqTVaA/m25q44tn3EcOMl3zHz7CJ4Z7nu3m4HHPHetMXpsBKpG9+
xw5/VataFKFwxADrmiAnoU+gn5CrthrbYQSIMZwkP37hUga4x5BRJi0WmcMufTvRxDQsB+Q5hdtZ
BlTHQo6CO4tRWobq1/0vdkONlxRt1tgpJomEORa+a71EL/K5tbQaT/6DbT5bZNjAEynac1EUwFxt
zg0M4CZ3+L9DSCgi249UEHwelQmc8xZlM7SgqoimR1VVTN5/PND9yX4AtgQV1WeBgxTsQB3TubJ6
COcy+09IVX3FBRGrDhv/xFLQIP2WLWyak/Neh7X2Dqz3UG4qRbUJXwy/HDnBS6e7YNAO0RAzwrJ+
qDv73C4F8KYCP5e3xiEKDJ7E02vNAx2cSXNueL93bP5fU6U2xZpwbY5CXTDxaesFcH0Ho74FizOp
kaRyMDvw2ruv0mtcgTHAHKCb47WGF6ZPii47uR8HFvgWIEQT1UsyJJmU/UlGA6I2WBLLcs9yGCbq
eZhuisKZKwtGWiz4NSqX3z0j2scdk7gcdKh9l2MuCnEX85XKwrfzoCY2kOFh5BXfk9NDBKkpyHl3
Ja7fZdQRI+NMONsUp8iBljgNze87beST0uIKqUirpiLOr/CheVITzgVGs814yaCH8C6yBCpXjZCU
ZTmTt5PvkY83ER6rPonttPwFAN9EMiTLMNRwHnHZ124nS5hqMsLazPpGO0OMnWQ8nLBZO1ula7cT
da+oPAwrbr3R8d8QU2k4um3ax/bOrvr4qk3IzzruLw3+38eMiM4GuevyOqsmBrQ1IgdZMurw4ton
yMiUfohB/8BFy55U84bvd/P2iMjRDyhr49vo2ZZTvsmswY+AYtpoUyg+nRwBXxAQgZQRQEhV1qe3
Yi4DFfY2jv7QdbuoCSkk6/nrqU2RPhVujje15mBByurG6dD5pSMZmPv6pP5h2hWtZ1/wHq69jS2s
YDKDQo+3DF5Is62gESGEXPlGsVxRTrh6+yAnqgcWVfQ5Bec9cYYM4c0KcoI4dAteMPlSHiD17zsk
rHQ5RAxq2Hnuv9Rw2O1BCuq3R870wLqS4T5q085X4XuVaFp3P+BGdc8Vb/E3ZA+mrdWQ3BG2Z0KD
XGOsz/DG1ftX5pniMLiJ+FPv71PHKdaeIWfg0vPxofWe09VYWfr+eq6Tt50aJL67cA6HkKyKMEzp
w2JgLHDpiwMSvNcDMkllvTMVyQ8s+HFOIBXADmOBaAUFsI38gX58N+vQJjFskdfhcyC94XRiO9Me
Q0Zt0HVPv73sDjnL+AR5w8K/36/+nez7Egy4BvpaDbODv16f3GcOzrcbYkQV9QYLF8lqMpA/cMmU
wzEM1AwmocXM1X6FztISJPfwXyzbV2QfjVQnt72exe/bukZrygTZKFlTZH8V7JZqFazkgioNksqd
vb1xYQkSE0+0QiLHA7EwJOkX48SQ38mWRVDHqVd9ZQEBQrDnhdA4CQbUkwcd/yg3OJ9Fj55R3ypS
9DPtTkxHHE7Vx+5TBVUcSiuixlDQru0USKdqS7uvJSuA6/o+4ENrJJHYoCVUroEt8VWaqsTngH67
3dRNcvCWi9G+JR465VPI1j/lFpQPa5CUpkJJZLqdq5TRL5vVhlbhR9j7Q2RCTUeV92LKlBLni5Mn
WlKmgb5IWSziCq8HV+XeEdoI+2Z2WW0ihxXsaSL1Zm7KdgpfK4NWo7hJ00mn8+8VBVtSaGvc2d76
LxjBVW26NxlIeA3EcUm0UYAlArKXQAkpoqTAcX4/1pEP2NiH/+V6sCXAL+snd6l9okFcQDnNOWeo
eC/6YQTRy3hZJr1ehlni/L2TUtilPuoovqTuWXFsIBGdAdnknCjU1cWFukR5Qv8TWtr3e1i+4aps
TYCyyyfDgC2Flg3GKzTLYt892RHiaa3v7Cff8A42xNvIIibSAu2tyOlGqDsZE4zOOfPBkGhVxjo3
zn+R7iqBZojWKpEwBcXTIBAsmzshSREcxMuWE3JqbyuPAtBfUBh2JQ0X60V5+vVuP6qVvVVMtnAW
qhCsmfFLwW4gMS2bgUkqDaRcOZJ0S1ArDPIw5Um7bbXRH/bqEPS76MAf05V/myEmDxWCy206MAqg
Q62FGQOuApU5kIYrmgkQ9dUbYAFnEuTagELxQZ/6H9KpaJy0ipYEuUGbuY6RYUFgvx/CZwrP0G66
tM4UpvHURu7wjPzK7GwH8l0bj0QYQ0nQfN0oGeKUUh58GaFzNw0BcrBh3IxtWQII7X15DQXNzEZH
WcALfYZOHY0TjRU6DKWKvAK1KI79LlE782PQxU//HvnJagxOYewvqT1S+Mwrzm5wWjCg7lFxkRGb
zKHtkXd7cYKQwNyfaxJOrM8Ka+vxEIK5XSjk168ced7yksrUdW5jrkfS2fYOo+XWBg9lOobk6/OP
GHon09ptpe6ZBBP/azVIqHlLptbamQEGdk74aySzjGpncX8lZpCPDVNY5fpbLvYM+C/yp//RxI0p
8+VKilbh8jWBWvzla+rEAH1BZpXevx+x9bsCbsPEuiUe/sNdNZyUraMOpgerzjHQVXJoAJ0JTdCA
oyTXWdmbxMrxJtYrZbYVD5q3T4Al8XNJ4VRGmZ0KkZtnXlqAusP/vKjSFqYzk2NV1JXej8oG9IzO
GC+ckbP3FR32C0USvguOVEVOXYJh2Hz46e6FvoJnl4GYXgVqwlUmUgYcGNBYh5uks7O8Xr3TtSZb
D98Sw1670MsvTC+oK30TmGemz+ScnJLaHVa2pa79iQS+Q07LoBd/TYeMnxJRS9sUBN336Cp8YGq+
bM4Oa2E46OJ5kv7Nz0EQaMu/CnY6UxPuYZzkyOMPn86dtPYh6P2OL+JXWgUuqaf0v1kDY5XoIWKB
6HZGvMQahprNkzdcAMPP2SbzTgiJ3vZXKOweZaHhaqBWr0KGoBwJS+/ZAIXO2SlYwPTW8yA8zNwG
hJBsHSvPlTRoH+acvYo1eJFdlnX7QAEZiJdALW3ZhGWcSbp88gJvM+Va5aoLpGs7N3cinooq1o/K
rBO5cby7+qIOIA96WILxkdxne0MZFFxYAx9SNcrwjjYEgZEdmxCsryfJrrvxAcgu0g4WB9T4Bq+v
IKGaWefBc4vvG5Xf6/Sp7WsN3HtapKCd1bNB0A6ngWf0JQhKotqoJnhlZw7asSFLll/qBNji2sL/
sunotQ4ujhV16LpbVLdGE1/PfjVDXyfCdxB7bLLyUVlu8a9Aasa33nie6rzP4cHSfpARAF67cQJq
9V/EI1+DWxP1dCt6adFFPZ96/awj75YGqhuW82VI0ECiRr2uBVA+KjRkeXym4OLuEC4X0yHcylyk
LB6e0w+jwD3oIusbQ3groXLwGlpEOv3NqYmSfpgBBXjKK6YW+y6HwZuYVaGNMLQVQ3rUx/C32I5B
6pIaqK+9e8/nroHsySHTKLLpBDF3j2TQejZZgXYQa6axytKZNnAbJ8Y2PsFoMuqBPAHcrxRi1np5
NxYLblaibRXGHtL3AgMh7rLUM5jUyetUdA7wyR4velED3hYvTIrlDAEL99Rf88Y66yJnuTfFjARb
Mv2x1vxHEJY3L9wy0vs9qEIUnby2yReYuqGY1PAz7GAsqhIqKDOD0Yr2j4MhwX3b7IDfo14I+xnC
A3WzciQpIApDPY8cHW2t4uKXhvQN8L48p1InuQqVDzaxZTfmpphxwNjM5u0px9i85XfAF3owoh5Q
tEVVqhUyJ2kOLX2/tQeD06J4/H6rdPxsP58EAaaLT56KGLhSYiisbilLvu0MjNghBNjeYV1pM13v
Bl3Z1KehhcVee5//UGPyvYI7HH6WFyvvDCIdxp8YOPSMGeUrLFj+3PVpXSbaxJHL45ou6t+Le/rT
T0HnIpK34CFucYoYUF560Din09Se8mqAZL8FNdEMEyK4aRfY4LN8lH3G4aK1x9RUDOGOmHytXF1E
VwQiYIBsWI4GPVqaQ4Pr8NAxM/VafVCaPB5IOizC5gGWFcOMh/wpATRjzbnmU4RJoaxPnK9WiKaR
ZfbL45PctUSQMD/89HAOPuyi4qp3HCCG1Tp5arMyFG4HIuabq2v1d7QHoGLoqaqK/P2NyV6DjHV8
jKOk/OXjRG9Z6LExaquevWqTSs11/m2ILZ1/BS7ftAt25e4WpjnE4dAOhoCQlG0a7Lb5HB8Jnsc1
CkyTtlYvblGQ9dORdS4eU4/DirKuS4qLnrHCQZd/7mND3AlG+TEVDze10NfKAGB/XiSiqJO6q2Cn
6B0pKYjMCP2qR31GdXcpS3bPyYGpVWo+wBo55VAh9M9zf+3PbI7kaFipW1DQFZQRWlAb7IewMvG3
8MWsHOVcoDZVKHi2KZ6Qdw/hyB0twA+q/zHzFljtz0WyWKwtTKDMeofAf/f9wXPX6BBUXwua2e+B
7uGGVHca7oAohd+NQpaZWmn9ePz7YZ3CwY57ZmwIs/HKSgTAnoVmAou1+ceNFVK2tz/9FOM2fFOo
NbbDwF2CaeogEkMR3X9J0YX31JFm7TA9BCE23gL0iwvWj8Svm+0vy5bgRXIIfB1Cu6ofc7+6ecrL
cQKpdl72uX+4+gvJ8A/cCxm2QQbw7GULV6e3TdV9mwYTJspYhjLdbHcsDVAbMw6JV4rJtHkOftBQ
AfCcrzxz9NmsNEpDe1uiLKEd5YEijTeLZ0yEVURF3LpMA9vPXkbYhQnBQ4dFVw7viSyvEvq+9LMI
AXbIprcOh+iSykjAHDMhkRXBIhnFST6LO4l93NoxmgP+yF3tWB230ttYjefWHjBAiYrejSRD8ir4
6ACGDfg22qle758J8yIL/HYNYu2L0xD6k2RMS8B+8pPRbTSpnCEEM+4bMbb5W28qKZIaHtANvow/
N/kLmobvd7yre6wctdiM7rs913M9hyJxDazguER4KBR0d1GE9/w96lWT+zuImr/s39/hM/u9mpQ6
oyzh1OkFzzzqlYUZ2JQ+QO4xWSrf+Lqo66TZkGzsda9vqiZuKVqtPirHKFJTVqzk5TGwXoxN6LNk
1QyCd3PFIrIAWX75BqlEz0O5kTceT+XEnB5mg1Nse/Sp1d66SF9EdqpQ3GTIn8FL/kKTchiS18mP
NtJYy3DFQVTHHV/gGgt5fS74qG8oYJcDPn+FAGSMh2rNihb8qPum8Ekkt2ldSDEFv+dNsxUAzq08
uBYNFWxHc8JKnU2wFD5M+Jue59FjC7s8vscpiobUxqtsq5OrYoFg5qg9tedMuTVc6VQ/W2jq5puE
V2pvHqxsaSyPXAUpX0RcT+9QOtyv+Qk537S82Eos3FJTrLvmph7BSrNRKg/hthF4uShvtCuTLEL3
uwphUHEIoxkTvcGh2SCEObTp6u/lMOIlS/wVdWuyqJO75GH5ICc7oFzc1j9cdTXRZYK1T882oGma
t12mNan55Bc6xs00pwjIbEcbmdlYqHm6icPfb8NsRMOOokOCS3ByWyiJVO+NWTKMnwI6LarfiPmg
w08KnksX0eR5mQklnKaa9WSGuDseqG1l4vjClTEhsTk3NEcetuK0XkVV6G6EkyapDXycEUJtr9jN
LmePaEseoi/+71WtneWdc5ojOzvCj5GzW08FuphYGiSr0ie89Q9uGLD9XVkkv2sFSMsie1V0u5H8
Bp8fd43fzI+xI0zWDLUF1FcBgr3sxYMv+VDm7rmOAgCQzhblshnKbK6DbzT6shcdqny7cfN4cI16
RJIE/rdjNz0fdX+X68pyQHKfUp0n2YYrR+eTFCH9WZicXRA597DufdUrMlWPXdwu8FBwIJGD8sI5
IdjixlG95hC0Fp5k/Nm9piDPd/tOjldvf4F/vRNITXEX2lmySwMwPtX/Z+OggKyd7nMyrDxTcNAy
gZZk8LZ6Il7UgLMTlhkqV6f/0oTccGSJyatIFL1oEOlAwNRftaTudfZwKq+OUfw5a4C+oF9XEW0o
OvCcoSa34YEvJ700IJuYylMK2eogx8yZOxWG+kI6Dt3UrMycAYzIfQXoM4k7HhA+/PwLdK/R35ak
Sq3JAl2HEokj2plSgYMjU9UDcnJOJ4Iac81M00v23FcmrSDVNuhCJkQAQi9KYWFTD7cKjRp69nBX
/zpQvm6tmf+nzoGxe3SeCAXKvIAWT2lg8vJwWvnUbhSLcQ0Wmceoo4kTU0EPPNIVhqRPa5Xlz31o
uO/QgImxQk01rt44dYE8NOSPl4RMtNB/skrs8FXy1EFu392T956Aj66csJF/84Te0J8vGYaZa+dF
Tu2jfK+A6qK6rqtGL95/8a7dHsklDEJb83/UTj+nRvZQdJ3Jvfpw3UB3VGo9EjycfQkD/ZEhJ5sQ
TfCBVUwohdRoKFEjRUlI7rR74uokvL/qhwD5XKNQL+C/mqK5jFilz8KPVfnje9G1zWXPttNy0g8X
lq0mm6oMIHre4bLc4lzw5Lg+OzJD/SCjQQ64jQpIKmDv7tHoflg0W48flQ4m/OIZyUb/zOAdVN+w
3SLeHOnEw2Nw9wg2KrFKU+IYhGDN7iFunw5Pul9zaFCN4GejOTJQ+nHB7RZk9auQia1RFd+PRAiM
+4SBRRNnEu8n5In/PRlSKHLve3bpdyFy6F6MvfkUY87mYJGPrJKWzRD4fUgt3zoAVtrVDAgg5hAv
ctonNTEGhdAB6vEGbeHsGmuVgDwQGJh0PBNUa2w2QqWDLyi+oOXBkdIUbA1rkEV7Kgcbq1eNv9qW
iUrkLK4uQwVUor0AXJ/zJXf7Mwva+MItntWFoiDtShz+1f8A6ILrosorxfogOs3RJqQV/YxrQAxN
2O4S3VhqQPCU+Jv1VEosiwC2lZFCKJuwbQUN4sTrDrwsDhyVS/3uynxY9md5MnAulT0WWhk0k417
9t2TeDOrv0lIW67maCQ2F8gYmVEbvNWj8X6HkQ3XPTptWjmvqsX1SbRcHdXObDmnLNM6vAusvFLF
mzPm18sh5wB6yDfCgTvoP9Wok58aAVATT7k8VZq0uTa2Pfx4HVhunbdCuG8myJqRrCB6MkgMezFS
p2WHE721KcDZF7F7A/aIXN8ZKP6aYo0RZGY9/wFokaRqIdLw+L4p+1Ox3mMRumDWNgDMVSAgV8r1
UCeCen7CdZpwZ/IyVNU5oAOS/YsmHG7zOzWnHhcVa7Qz28TO8VowzAKntx3YSgqPNFLTngTR8j/Y
xz+d7jXrm9mJ6DO8uAhTERHJQlfuccQ9bZWAF+VLQypWJrzKJrcRrk3r4RTE27vUPYTLEdKm5yoo
wSPIgu9T3YxYinXIzMnuUbv2yCWuoa9dy4/AqlwHV9JnBUmQ7cTktaMej7b30J+ofEmrzfsCV3hB
tOqPwEdnUc/G5U8Jdmm7QXebr3+zdqHlO2Zjha+0JzLgFSEh6qeEzf55NKda1xbGtzYotHXXPeAV
HCzZKGSas/d8tTug2zlqhraQwWk+VwVIWNPVZq3GUbOw8VWhTntPyOi7W91iJEOkT5whg8JcmTMv
a80m1F27LQAc9MFEYmtj9A65WKf68BSgvxq9OQweonjLq4PsR1ENE8ykOzn0C0PJIg36125fcfMT
ZRfQZOp7yCirE3UdTtHE1dmfiDi2ldS2vrrehf5ZatVVr6MSR3UtB0CirCJ8pl33lvsbYzhKgL2c
QjFIke3ZLgXfJKgDY7tZRqrLEeDgYJhndwQ97oEt5GAe6MNNiXU9Fla/gIP959OkJzgBF8ksj+8o
P+JoMlh1Jo9G7yRjDtjN3ceQpvvzGfajJJdIroog4nKukWthzpHcDi+HxIDMTCE3Jz+/Ls4CGTP8
4jeQD2aguJjZUeuple9ucN+7GY40C55xqjP8uFv5Q7STHZVlK3sa4QD0SgjTYh7/HyQewDhfUlqD
gaOvSZE4GmQyygaCY84cPnM7ARI8HocQv5OP//MKHhMRam0ddp8+yITewDN3lG2ZuoWwOD2sU9dd
yDny/0cetMFTQsV3gHQ2tvwEdwO4za9t0WQGKrceIOrWh/+LIYnUWRZ0e5SikbvWd6kVnBOm3+JN
K6QtzyQacQ/TQK0WUiK9J83UN5vZTdDRpaYnseRZZ3OPKF0M60sEuEkVLb/NozjoKqVgwlU37iuO
32ycvYYOs1oH8hLbzAXC0AMCq6c86JQdj787F6v718uU94ygEm13tFKzQ3k90ybPfn4n4tO9Nm7E
A+X1zdCMpXq6wJS0RTgWJ/D4spUNlSJ2xZfIgv07s4VablYPWy1IVJLav5T/93hbdlaaHcd/BDIQ
wd5X/GjNt3Dg0QHnIxHNcC/32NybNybHa2I0m1Dc5j6HAEm9skYkdi1y9pkw/FAvkRwXCmMzw1wf
BOj/aGjcqOwKPTf9HcyKbqk6Y0c2fLk4WFzr4uSm6FJ2zHPQW0Zo626BwTnMUBVqkmtbBCQMNB6O
K8yXrmbPsk2XS1p4xPaT06ksPSE4mcvf8/WaObTlWkw7SDuryheXIMFVyIyLCu0lwaLsGJ7Ie6RX
UBp1EdCiIf4wnCuJjLACX+B4bkSMOYwg9CbAg66z12GVDkm34HPEv+Qb0MSAVN8+oZGTAVCH4Yl/
VrIhv+ZVe7T0CFcIZo5aFUGL9JEdBbHYTazY+nSrd30YHWarg10BUv4BmToycw3yxtCqaTJVW3kF
IudWLyK3Yb1ibTMeBHiwS5wPMto0NubGRyHV+I7QDtFa8mTbAdLWCA4CSwgsDint0iN+N2gDCHRJ
bVJQTDkr9VESprpPj3Q/QU1whJTSYxc2YJ96YZPVNHJmoO4VhVMEYFlhc/IiNsivafGv2qcE/R6L
PC+K0gXPkvLEwjeNFfCMCz4PkQymJvo8O9TPKGyXOiaf+XUTDhcynKpl7x84mXWmy6HPeHjh2P1Q
JopX+cooRxMWxL6OeiczJt/G8kwY9xSMSDQvTIShUkjBlN/VI4w0UT4T6tWyme/k4yGfi7IVl4SR
wGWm2M1kefo/Wf1tBnTuqitIZ+tT1wIL88WMHSPGX49gVjA3jir0ef8lwxhT0dYN3bD7m6Scz2CI
opq8muaBVdSHJmMhnQ8ynC1TiR9uY2waXlkACZT6ZUMKZB17V0zJElCXT6+bX+0RdjJ+AbYwpQQS
2LgJbjmwqxcwl/m+tOECGRl6drgvt/a1VOGKnjFRy/fNml2nsrc3+GVWVD+GR43uV8noCVIOSJYJ
YnkRdRN/etuewRvdg5UDopQiW/XcG3lrdhUHbyPm/rzMgc0f+snLo/Px08EjjmjwFlbuWhTTG+vr
Ljosd4O5Lrpwv3+Kj8fstDsaI3vQUfkVLvJtkeAffrFSyNdVoDnYy+LqXhIxykSgc35rsKDxMg6e
Q3V/uKytmIdxEuurAa0Pbd9CRnsAn28SkNitgHpLIakutjaPp4o6xptM9LrnpJ1QPlaxcxjsd1dc
iXlIo/Ky6l4UZQGXlyuZ7VjLaoG0nW2lTcZrQWjGgl9UZ0Jk9phAP9uIfZx4La4c+AN59L2P2CC4
xSYZFbmX9S3PRUSvgcrkgZujsuDgxMfvb1q+gnRqhbHUQYJ+FYu9L9R4KjDid7JHzH98RWJAC+4D
Kr3n+1sxZAbc3XhaPHuAeibIv6nhEZGuvF8PVTfi63IVJmE3StAjGooDBiQ1Ra7s6M7uUAHWnf4u
6vy64FIi77y52+ysc001Rxz7uNxAW3L7vCMWBIslc4QXobdA8+1musY+fY8Cdec8/xCZirNHR94y
lLFMrUB8UYZwRHVVx5QVDOZVDCUQrd+oKHB7PRYlQdMgD5bW5GhSbjW5I+v5RQiCv5yoZU9sakn+
tri2sAP6k7hEcntxmKPx2TG+zaoOUkUlXTp+yrPSl/LbVkiiRqfTKk2F9KZUwYjaPBckeHjFWU5B
+vJpTFA9b9HDb2/XHXpZdhkaecFcv/JQfp43DBOO9oaIM95BTfhoQLttqP+uVbSEnQ+L+YgWAFrB
Gry/q5e86aysa1C4bfJGZv/jxSs09TQTewyNJePw8rvlsPTcOHFZTnEeBwTXyjo/rHS/M3iJ8mVS
b+KW/l8BDi9QSFUY4NSDRE6NN8JgEsJLaCNzDYOCbhJ0EVxljboOa8LHyrBQaQKYjYpd2YCg9oNb
8D03kkodyQGLLLKXRnmw98YjT/LL88ZTGSGkPYOs3mq8Ki/rNtp9mJwsAvTULNZyUviPgAFdXq2D
GYvwsqVUYqWlGftZkUmFVDzcpnpNfqFB0+Ac0C50gj/AZG3Oj6AM8WeEiRnawqB9Q3QXrIJoYY59
sxdOPU7hmOGplL6jQsPmh3FOp7BdJe4A0C/bZAMdI2TlWB0onrx+mK5z6zquH1kjqeZuNWY3Qyts
VeCtcbuBt8AHN+U4b1i8UfIab9H7rkc2Xk2CphdL+LV6inGr0IpiUR35Bhxfx3Jh8QFybgOicfv0
nazakH8AeGfAowvKQEpPvrUwvrrQg/WGpeQjWDPv2siqbms3cFTmH90094nuZtKXHuM2VP0A8dVX
ksrkJARg9gKtLAfzYMoxTv5twlrX8q7Qt32vo4S30QpQU9oyFct5LwQipNYwVB/0KKXNL1+/mFeL
dqfG3jdBau25LBQAOLi9gVMUip4DdfAYLh5TABQ4/b82KGn/3OsPCQ/emp9IusvfGsY1eCVMOGZX
mSo3yjrZOkLxTWBrHSDsZKHaTTK9RfDK3O2nynaVDEMrNYaAGJRw9GtxY+1eKruxp1LtgZW3Xh6i
A+JOiRbwZbszO/1gU7Qch8reU/JZvq/rswFHeW9248uXq5sYxCX8UrYTsYkmLPOEJxxhZ+Of0Drg
YTObKJK2k2AkyjYapb1rgQcDXl/n4EBagzLJh3dTSqisOW639ma079mnZx8i4X6du7W7UDruzeHK
GvEDPvo7i3/Rj/9CKDc4x/wxUU9gUah213b6FeINFM5jr1X78lddzg4yzZrm/3VwlJ7W1QQLhxTs
/dT9fqI10Bjhs5svG0u4vSULicR16q8w35g5XKn3eCUgDKm89Tq6TXURRQZ/ddsiCaoxdyJruynK
cKp+dwAivua73GPVqg4UM0/yRSmj+CbqzAUal6VqiU41m3u2HDEOEzH5HjauhIvxfwj6SYkK3yF7
Zv9yG3mTrX9gHgRGqPGXNFhVo16fDYUCxaM4+3r4z9ab+Dmz1Q3i1o96ZAkImdBjnDoXh5T0bdji
pMURlQgDNm/UXypuWAYoJ1Vr1oajheFgEkDxujShV5W2hXuMlOFXlpKBaLM/tb4m1pmpu0jx16Cp
L8BKyAl4PVzGC21e2o3nVd2GBDqnBAGnMc+PzMCamy62ykBn4WJ/kCzD1R6GS8y0VCYypijWKAMw
lb+2yEbfHowvFLrVrSC+31JBavVIEhpntIfPl/PLAxBHV/ssvtrxkE5jc8lfsGfl72fzqkdwXRiO
9N99W+Jk1D3XxLjDX3fPHl+98Hwq9F/UjSADmB4a610GjoyBB396YY9eDXUDjpo6tObMXVB/JGiE
iGGLZAk+YRpJwbztILVRPtv/UPkVT1JZRWxjcbHdFo2FopKsr1vTDsOLtP3jQoN782IOEjJWTRoH
vVAWQu/m/Bt0cElH/trvFBiI+Luq6cC6mngwg/zGANbv6fu1vOvo2haHMYiwMiaDSt7gmTPbeq7P
cDGB3O3EDMg7ZNW7UdLQkL38wA0JY+Qqi9zQg4pzcB6hu0W9K+jpMqmA5l9wiWVa+iFXqZIEP700
isLRZlWCRPbSzbBdIp5vF/BSF7VsmrUe2A10xhpVccGiNHQxr6eqz6M7poQQu88fttLt8qQvJMCb
juWF8LPbj8I/ZsMjVscdt04V1KYrwN0/nLDdTLiKk8k0mgPtez+EIYPto1kDWfbqytvu8WyJya2G
DAn6UngcbkEG4EExLZ/Mjdq0fKSnCoMuZMVD0eHDJAq8qeuEeL61HRTT5aYZotogqYt0iWH4pvEG
LA9EEddw30AXLvqTkNO1kAf/2ZGTgYlnavhHpqikftyqboMqKl5acst9ArH6Ydc5BGUMHezZhwIW
oeOT8QcLIAa6MHNiEjpWjuLOGMbxZ+QE5wdxzKxDeJWnOVbrqdUTZMbUY1pyz8yuVI0ks/SYWeLC
wJ+Pnbsvy42sq27Vm8LsAq1/Ya0SX6TOD/R4n4nfnV/53j0hQok4+H9E93gDtn9uKp7tBL52r75g
TF8l/7Qgby1HpgTJzi+EqDJ7mTwwpTfXVJfjQCthAke41qYbG4e9zCKDJPZ77J54GmyjN1f6Ywyj
+zQAig8LPVrvZxyu8ZffJBn/iS0RwNt9K5zDsUoHjTVHHoyTyKm5+6Vu2pkDM4g8HggNjLyiPySB
YQ8WhQJ4B2nZPegLd1BphmBTaNAOIHAbrjBsCxaIyJPdQUOslbeZdkHMUm51ZxDc1qBA+0B7Ms/c
JRzTQEUVk2PWZCYZCZb7Be6CyGRsAnXDDewoxsBYEoOLBdb5naJLmUUTDrTesH1NbY8zxHHnBoQL
qNwCg36fN3+kIRrvsetiJ2a/OWD9diSPEl9pus3qVetzYfUvuqsTcYVqNNNxqsAAlrv04t8e5J4P
VQ8cz2nWkzgvBLdbrAMrcDppty0vN75XsN77QIk1VrZ31+SP/JeUrkaZn9KICLMzy9GHRJxvAET9
rGGAtv57Vq4spbTXM5pv5RTbl36p5gC9NnBxlW1jF8B4U2b/N9sH3K2VNaxei++gvYC4Shvs+vTT
ss/ChEJ268SXCrCVcKdwcDBAajtvNokAmFEGXFw2IzAc0R7kmfKx4//zO/bRYRZpzELt/uO4sU6S
h/aAJnJArjM/MTzVZX/D/qdKGcWRjiQSNDR4pt16uRdd3sePChpXgv9TV4xBijlcZi1F47jJ4aGp
HVtJk8Npayq9KgdLe9AAG0ZVj7wWfwDzTrVn93tYbu4ag5146mNvtcxK8cnqsRK3UMTYqE8HzR94
dDjQVppI8Iv4QbW32mwB3y/tAHO5nKbY+B5lvloBgLIkLdTn7XSh7JceMtAScXnvBQHkUrHQEaIZ
awxtHp+HI3tPd5Ca5hr0WSjlDH4GdxwKsZ6WjqO5x0ZG6AgtnjUfmw0sys6oJrrvPohk35jko95g
3xzVA88QanhglE6+YmWd/9wCGMLSl/E42zMfy8gKgSL2qzKNhSdbsmv+ZV1lwKE/qnpH3m0kKfBO
gwK81lKj6xPCqlLxqkAZr0oVKbYUXiC55mSHDGDqylk8evIZCAAxCPnlUW/r5qOM0HZDZO4f8RHa
gp2KnRsYyR9iEl17qPobP1APdn1OxWx/zQsQcnYm3uDSaJMdDGpsWMurOHGXJ93XPgvb7MCsIwvF
JGyKC2K8qMwp1ig9ppnEAVVgVHvxS2qzFY/5egtLmWpEWtXtlzTzvX3VwiRMzIIs1A0I5TJjwBgx
kLyFJjpCOhIWTQEQtjOGw/1T332b2e82kFuOSGWvY63M8CXHQJPM8Lq9piIzWBEwM3grcqg7it1V
Ol/fFGjTDosbblbOlWkcGLbgZCeGvNPGb/vK9pyfv0+VpWWv5tc5BcaXXSrG2BzA3+xtXbCCEDbw
UYpXJKjK4XArSwBHU7S79rhm8JuF/ZlgYCSeVDUpnlxJxdxBU7NZnZ6TIO31A8HKQfvPQWOJkgVq
5XltAwPK+xfRZziF1X8QBEdYHTo/ZtJKp2Ll3GzgOISeCDyCyoNy3kT0cpZ26/471ashEWNdVx7O
ubRfNG5p1Z0FyUTiE9zHBqc59vVrW4XtLRR+kq897hnsQUP4sQEP7jT42jK+5JxVnxd4h3c21t0C
coOEhOLETVynqHWDKq/jXYUSJV5+xqkRnCRmFd67vvTvTKEkbcoXdL/ZpRmbROMvD9uu9YThF0er
+XC8APwqRi5FkAf1B4toS/4VU4PvREfdDSw4xxeaJJGIOZ+19CqpKSW+g2BbUtmxvq0qPaK3cFcj
fZ3ZBxrX+xiHfhEyAUSl3Z5rm3eoyYX2SJ55KAzT6Wd3J80XXNbaXPjNrcHt5M1T29yKlqHLj7a4
gV3/BRXnG/WRgyM7FQYGx81NcOJ/SIOs6qinNnlCGX+JlMlZigS0vy1XXOJyJMbnOWqWoJTKfqRj
Pra+XpZyawf3JZKXSkhDM5nE02O3pTsjCVrcgOOzIB/J0TJkfG8bhXSQqONj7DLnRcHvQXcjQwci
OrFMBKrZA5NF2Ubqem1R4NpnnS1Zk5slLJFYJbv4/RbZZO6/eifofQ5//BB20HDR0C/IEf+fmc1l
bnie8URko3J0h5jnfbqutb1etoJoDrnNwNmcMYrRDf8p5uvaLBOjs4tNdL6BBJPGgO2djIDElgBL
HQFmBUXyPe77uXIR+xb3ihiYGmYCo8w2nvvl3kI01ix9A5AmTgCECpEOpmHDfUNc88/c+M9CYxbJ
hVyA0d8Uh/dEk9rNfzfkK5RsbJcJR6zqkS3P5RRnWg6ceUVyKVCRIthkP1b01De1wbKpzuPn/vJe
obrJpidm6rzzqwPz5Kc4brhyUnqxpDjpSPjJWsK2W0SKrlqoWe3xzDGaNpoh/zQYplEs9oe0ErSm
u5u1tuELEiolJJ7AAy00fsRvyji3a2mEZX8GxxnIVTmnhde2ZP4zm9IlQtdPgwqCAc5S+ulMzLez
U88cAL0tBYDUPbEKeBeuX87UKfJSrQWO6nqoQ13u8asxUySFDpmooG8vsqiSgNDibtOq5RDhAANS
KTBCAIWpd42IfXL3CcZIFMpwJqfNNEu0o9XpzHs5N9Bh+Zi9PG2onFklYIuDg1LxGYlLjeVBRQgw
wFxILJy7obWprhWOCJLRJH9uWwgr/Qzb+Q8y+SegRp8Bcjnx24em3zlyFjyGIcJ8vLFhGRJtSO9x
kUls6T3OW/l+oegoSKnYAXS+CpakaaDIgQxvnwJchfrEI8KHBwCMOIXINmLWtDq7dhQhyvmpt41M
hQrFoEDsKi39nVTTRQEqjY1Yqlvy3f5Mz11R09SA1ZVHetNmEDvJ5WORle+Ucyiq1e6DnLx+gKYg
RCxSzOoGUZmBxwfZg8mYLkAF+nJkiF/Ot6cS3x6aKGXAJrIei959geK8WQy27hCPzbm3jVir7LaT
sIm/VJLzKXWyCsfPsznd/M1VHv8QcIa+ppq9IwGE5X1H0AxbL27/NcwnSZl4aD6vu+Qq2u4SCDDu
iS+2/u9s5VFLSv4jb/hK8AKVDjVDTAczxU12u/2ojRo0m0jvlEEYFyNuHJy0gkuvAGQMGzBbHB09
XQNYkmEnvonCVZFg7Zy8l2ezfbRhJTrNa4LHyJom+ZJt9ZmtY1q4tfN6DxpJHdVGVy4hdDLT/ZXY
MnUv+JEd1md1Du8pOQZcBKX71D6U/QxPKLzb0ZTbT9vEaPq0AZ2LXmyCSDhYGEpDzVekGAxyKlV5
2Lzq+tAMm2tAW8p53/Q6HVlRvk2czxu/LvLmVnOZXsFvtGj5cY2oOSI3JEJ5/Sx7n883JEUi15eK
dJS4uiZOc18h5KK8s5Iu9dyVpwAGtzOEnGildJvr7Li01HLsVz+dwcygxNQbNofzS3GV/EH2ZmHQ
4bLfRAxufOVaK4gLZvPQikMzprTvI41dMjvExwR+/sIKIoBVxaeNwXxnrleHx4EfW/Kqo70jyp3z
Bk7rktjLq8rvBrA37XycIIhhgKZVwngfo6RGvP/oyUnCHlEjXw88FUGBzXFiuP8p2L9vaN0QrCyE
AdWPgdkVDHdJdA1VkZyG4kTb+eWmlj8j0cGvl40c++DOAjDvlmSp/gLuNaRP5o7NNW8sLV9dRgon
s5kdW53WgZJY1bmUbbXgV4IjBYar4TAD+dJ5Nj/NFA0ss6KiUJE6d0Q4eMrczPm5VETtmcNafxXA
rpHwwlmBeQ7Jz2MU2Wc5Og9LzzWLx/+nbQhchgW+r+g71pTHYA6lSEz/OPw/+8Jr6K8GyuGqH1pJ
Hnp5fN1hni1cqVyPCCJcIj6F+pzsRj6VwI89ZqdFHZmAphDghkeqDtRK5VQpWP3tbW3xi52cmcCv
YsHqUoHQ8CLJoo/IhzMNvpkgnMMI0khhzTRvUSmlA2jP52RYmGmoec05HeM7/Ff7fyxECLoZvPVM
FzIGgoDhpHEUhi6Q3kMv31W40EV5WQYGGea9yO3ArS+pwyPSpey0ADzeUzE+AK/LTE4HthrKfiQo
gEF844Tv9r5CcUksdSz2vN1WutOVYzCom6eXKxwXuOwLrwV8hQi5ui8o0Kx/TJm3bGHzkesmAfvB
sv5CrEx1U9GvzyOdeXDjHeBmdC4c7nN3eEdoCO4iGWoBbHEVtcN5xYtWuhtsmdy38fgzvOCa07Zu
OjMx1K8mUEo7+KpCizN6dssnfNjOdo7v1U++vxb78ac25jOQIxRm1ZNc28O1gA1vqlmFrO8dbo5f
aeRPkwftK82sH6OAswQDaq3Iaw21lZ8yPpVa6F426zxRgZCkPbdn5RWX1s/bQp0KzhsMRwT4BQxc
gdF194OTmpKu/D4y4HmVe3VJrScZsQdjUSgma6hJ4G28sq+voOAxIM2qES/YDahJYSQpxWfcn/gy
l/onyj1d9CRz36+E+FPw0cbBzSewEeP+Q2dJ//d/sUxRMS60lzGzQemRYCS3l7+alLRfJNNagaWm
ePfyJp97BXyrumeBkGaqM5MB+wGfUQlMOmRLtyqGpZVN0nmXFR1kiq4ouP1D1VKR4mxW68iahzuW
usJnsxWs0MkUicK0KE58UTYYyvnWEyyGcY2fXnLoXDmnk4K2MUpjhgfOjuFVF+PSvXTSAhOgKoPt
pzefxIcR+lw8o/WXlrvgO4k2L0KEkfrydXj1uliNHc21isM00gzm9CyL6O65RaCGZBLD62Mata0x
K7Wcf/ANC4HfC8l9LCVqCfHMOQBPiUKBvwafSjglj46d0MEA9w79mzbCPilDBS1lpwfsSrxB47vh
ixUm46vD0F0th2mjQ6+ZmBH/SZ2bbmYyPucLf3bo8ghQscw/sTVwKnb4rVqASBTT9fLcwpK38mYK
t52OA/xkOFs1EBbI4AvtVC6OET3mjsE/ktyPkV+AMowRpbizJzlQGU+HjAsbzHBt9GkrviS9k3bx
y4yspwTv5M7uurso7/3ZM1rnJYFQq9BgG0j4OhO93vPTosUcgw+Ow3hFIx0YtwXIPjuFA1dkW+oC
NZrEw9VTgnEQbvVTKsg2KOwGSfyuf+N6XtRXlK965PGgJGAfet7KYycyCXnGT8dpy/dKAKr30MSB
lY/da1qEQzhZYbZb+YMpQEREU/3z0R57w8yVg2dqvShUB5m5/6w1I70cbx0MewLArlm6mEuj2Uy9
uii4wU/vniGHwk13z0IVGY7oVsJMvjQmBj+AWKN01be0osMa3VNXNImy1UAy4Id+WJsyV/2PG77n
bVl6OCCK7dRPk1LHt339Tj4k+1j68YYoEmWKupDpBBStc6wMoFVaWq5kgYfKW9yOm36LZ4wxOeZY
2bJYtmZAifj9+bnjUyZ2GUlevN5QTLDK+LNj0e7Mt8BaionQc1KPsZk0T2BP9KIkZw/PN3Vf8+2K
VQba/8rOVyRUwiqsv8qwwtiZ6OKLYsGIVUB/O3Z4Q2Z4lEJWM4HPl3A5iZEbeHicNRmtN3FRjXba
BE8TVyubeMLlH640KDISWNMXWcycHwI5iJzKEvzmQ15O4vVRytEAdl+OgjSdeJKlt01FSLahcUE0
b2BpDpQaC+5qEnHjHnDwFpXUAsAy4VAOaAIiJWciRUd4z1Lf14sxWcJYq27vVx5C4a7ELnPvYjqx
O3Jlw2oRUS0sjVs7ldF9cydTS3mibBCwzGDqp0KLqfTpIDD8oKwFDl89dYf8AsrGmV3mIN2a/lT6
QLKFjdNd/+ta4TvepRTrozWgbFzX48VuGcwnl1katJxL/OW+qY9smR+eEW5pj+XJqMdIvrO5Fsa7
Hr9EMvtj8npjsWAye2W8rGMmsNzL4H7xI6bIj9O+MfxS3bW4zXcRwhsaslPUsp/sLhGrGE3bq/Qa
2YFeJ9c1VFGQa/G8jQSjvhjDnnv/JqnFJavQrIygB6u+5CGcAQfaJjJ8C9wXbn6reX4Q+qWvAbMQ
jYt3cotO746rXCjA5YsCVGyBmuluWf4Z2r/4b7G0bNliWt/vT5VFgi96D500gsAGGDOBwgs9VHMn
MDxggd/KBubjzL5x6kt8GGSkKcjJwAzbPioj/xNLqoIfe4f902Vz8DQ6Fv/iSEyYgkAEBiksvAe4
9Makpa6ex7osF/zXDcQ2XzGQ3qYOeptOn/UAkVxTcJNH/NcvjrltV9Hu+vRxhrEB1nTacYcyIqyZ
S4/3o9cf39Jv5q6V6MT4zn6MnQJ9Ikq9E19pfA6DRadYOJNagn1lOMFoZFC32WHp3VQ3ADeN7KE1
FER4HUn8S5CfuszVziTRtOTl5hD377tvOcbO2G05x/iHi4nYKmsNXYmtREuNY0VVLMMW3GROURQA
6C/1DWInJems0d5plRL75PnoiCFGfml+KlZ3Vwd69y+tQaN3n1VbguD5UWmxZwUzx97P9x/JqT/+
DNN1hi/bEWEfzsmfyDESw1Geva96lwHyQRUHbIebjrymLBoIHKD5U8Otd8h8RxGZmTzDebtJ0E/B
Qet/cAebWh/7z2EAQNHJwwzqV9Fdi7SdtV8b4K29zCOJl3aj+dag9j9fyD1/k2N07eLMEf85Z3nK
tLxy/PksNDnCqPlhT50/T7N5OihGquF61ysptvNttCEF9AUoEC0JoG4aKFi35siwyrIJHeSkziVV
lXnt5QgCThdvVvdjhmaTfgXZ+erHbwMIF0+aMfzFs42XsufEl5LXhXf5xne2DW7QQ4wjQfTtcNvO
w0xUErPzwHy0kv5C+U7wQUcyJnowxvX2TS4g++mMr2TiQ6o6K8z3PsOS0f9g4LVimcckpIVwV3n7
UYiRzcYTWxSe6DLOp05WI73zlOihyl1SlSXD9vHrFUprd5emAZ6papdSP/JYmB5HVLNLJY9/uDhk
tWItdA1IKhsU1quhhVTFFCWej+wZS2v+BSqllNJg5JdCs32Y7q5K7IIOOEFPPWlW11e/inejJz/m
jj0qfTXNyMylE3J2AqqgDaoQAAu4xhRxXrvB3Vi7Y3PxUcdkKm9I8MUEkZnTC4cRYBzPEzyrPqpP
UW1dnSJGgWuok8S+voSNQ64QkTMVVLuGBqUY1d459AyQJYfa3P8Sx+I38FNY1YgPeY1OVXbepCiq
9IFSt+cQ5Snn1NCnMb0vz7h4VDiN7mJgFDeufUBGk9DTIXhsKznj0pGb1WBp/ucE4mlgtSDc/GL1
TR27/UnE9QznZ4tZo5NA/0CXzjMuytQrrnABWqVy6pSOgoBYQNYiUXbsbJ920TRgIzglcgYn7I9g
Z4easXiJxmHOzswCIMWU39czSxm7I0UXp79Ye/9Z1JHBTnqEms+cB9M1OsKVrSUww6dcUh9NLEku
dyVjIYneOt0yuR5m04cauRHJ3hie/qzUh9P4gdEp8yjdOXdl+QccuE0yWmfEm+xG+QBI8gxeoOO8
d9XbKIqwIyIzlXwBIXxxrARqpSmxqkpPYknBsSFPryIGI6WGstGckVqHH5G3LEZFlLegTjmIhNg3
g8y6ukebhrWwQ2qdak1HsCxq6A4fr9UCNhyXCrnDx0HP1Y/geI+stVKhngm+c3NgD4nmgB9bqyxE
MeRjtLz0Hsj5k1CuSmWG8eQRnrdffJBs9i5Dxb/Vor/uEA4E9nWJZlVULVox0ieFNnIG8cppaXbR
GLS2yOT+fAzCaVPPBhAwUfdPjYpTmCsVbhl4TuT+Z9r5jmwkRZeiw3k9NpCk7WO9EMviMoO1AJpt
ON4IuL3p3zLi7qvHOi6tr4Q8lIwB4GEosIj5vDw74IroHWxO5VYejyjLjlqeUAGr9vSAoue2/m47
CQBH8ufleqtm6w5UQbfirjsxIHULlMIqBXaYWd97U/ZEnaui5qE1Sl0v7VfzVRZRQ5nAF953VGYl
CPgwgKGkuvI3c2c0UowBZRHD+b5HKST+8+HdXDKE7bH7lgFmXtW4+X7J58/gTcUmfHiSSnpbkqMI
ibHsWXlTan/t9uqzzM1uxB9KSFBhc4shqdZPTJMkKbEgZzu+L4x9U61pnKV4Eas9BJDmgYA/ag4P
wz10N99MPSOEImuIQMOVrYpt5Lqsa+7t/9jW5fJKaFOIuT1LNx+awHEiyDbG2ssuWjuByVF22r+D
/YVkZaOXrOpwK3zHKzmIYalxUKUX09gf7ysQJE3uL27keVWRKAGBUFefaTycCqVzyOho11f9BHgm
QZVRAvPIrVdkNq61BtASemSefIUBRyJcxdbaaMw5wmeidCEZUGwJPmwWNVmCPHs36PZf3QXlt9VL
daV+R4KlqDq1SGeAs6YZsaNZIS9IH+fMFCBMSRN4iFCe2IpOS2KDvRLu5bGsjHVgtIkhZCDs+ZHo
oJT+MvSfojO4tU+cTBmwdT/hPUwVntsgehZrbRV/wLHFD/936Qd4au5vjLvvzVGz0IABZ90aOx8s
8lSKTW4Qu8bGyQzXCuXEJV//W39z7a8m5hI9JJca95MCdTuZvaTECW6Pg6EaUL3G1vvHKq8H3Wlq
j0yVRVs10tgypjCY6slzVJkdlGV2g8beAnMdYxVrvuJF/eASfkAl0QECJDVRDKW0bUN6aebLpUAe
0HXuswFwcH8YIqgOa/libt+pn75ybUWPjT4MjHQxj2IIsxHsH1oeBKXg2E5zt8o83FyWf3eQQVpy
0VdXVLCcHD4wxVV0k66w1lDQdUl/nbL33eKmKY8KHIYwLOdwmMjhu7qw4NiEeKWHPdCrDtY7kqrG
gYA70vlxq04bExjdgRLH2pvMz+FCvAZJfDCrKO7dfTCSFQfphdDIzVUQyloY5HnuBSySSwuWQMbV
fqXyxjDCiM6YFme4NKoYGPyFeFxx/43SoOFNCmaeFex0JbnyD/m+BgrK2qGZxMNZCwtl3l9ORyPA
sUrvGxGF9NJRO4mTa3+KyL6fu5kose7tffCc5O6nvbnRb0oyspW+ldFwbS8CzDdUVWOQapKrXASy
ElkAFFoKzrw2M8QgvSxq8WGuaxHLvhy57p8KOWXrpZyTzdnx/LuuhqlDVQ8Z1JaPBklZWM9t+d4S
3KrffeKO48PPmjUGae4x6daEzzdR8f0l++7eQPMpFJZ8aBAvm1XlQifqXTzMCIGBFQb2Cb+bDwjt
y3a0R1Z5cVtEsf7hKrcTbWXG+KoBdvqwc21yMV16+rCrxL9asS4xWAKoRGEKAyP0bv8EL0AqSpbc
pUUSsQMmiiFzBMyCfRm4zLRVGB8O9v6rIYtGA3SamWxS7ngpOcyhwNT8J1h4VrMhpkiQlReIJCAf
dYSFcsrTzcVQ0/UNTDXUL4QKnjvpmYEd6LpB4cdBcBsTcgjeta+IfR3vkL4DOkWeJZhDd2E+VTEW
Gd+lOSxxXXE0FU89b3uxvocf8GggFs4Mj6Du5e4BJdsCElZsx4mnuhxeMlay5bWCSWI4o2D/pR2g
8MdTrOAQYL9k/1rBoflp4L/0JFAGO1dTMJJHa+OrFH6NSY0uZX9mM+4bUDoq9o503+r8YCOK8QQR
oXhzl8HpHRxIaL1MZG8oDkh8E73c1eRduH50omZbe8DgMbHNGOlJAwQlF1BAYJ9FePAkGSf3Laja
Tbeb+zjV01JoOoJR/22gJNjoX5FvfKYzbATY1OyRF8le7mMUZtqL3u2EbPNpE1nhzsBXHJD8C59C
FOMji+KSFGmV7XlizPPpQrR1P71BA5Q05aeVvRzzkkQ3m4hmU5cQCjxUMH9IBdSdncHQWXFX/1GI
/m3NGqwqnbwkBAx8lFWfv66wFHRPdtvTpZ8axkmy7MohXWztY5Cm5J1+Eo1JXlW+64xEA1zYP8lz
WD4P8sfzUg0KPvd67NLrv8TgmQ1vGj/6S9KP/DukmWqmILrgpiJMMYca4P96yJibYuuHbDOpGOrW
Qq0Z7B2yGN6MEdmehC2o5jY1hrnvFFx5ayZuqGevjBzmcS0ym2IMp/UtK1RDUKMtmbDHPv2bYEJu
Yp/HQLaa3iT6LlFsZ5MOF+5WCvLuJMTXZWqkThSLGPy7Iu1MYWL8AfCQyMMpjTEoobab3HeLQdG3
yU2FQiUBKDfuVN1vnwkQ36ObUEZBC7WDxdw9LfPoTuRtOuyYWphDc26lFUp+Qhs3Ha8syq8J3C4/
uoWQadu5PIs056PG3GGG0DD0L5VHprZqBbhami3N+lxLdsvWW0PWu0scNN9VrcDSX0Qco7OhYyio
H8YwPcm3+VftPAxDLmMFAnGEBbCLFBIQBkwOAF8zDOf9AgjvG3vxgQe24W5KKxmVSRNqSuaM7DwC
mQnpMSI4D474ZgpW030Gzvyqm9HYnBjRjYlIjLkyyYkWaJrP4aKNhsvdglaXMj8Holc+W5VBfEke
r5XUL0BtDf4rXtDXMj6OBPxfVsb6DdHgUVC7X//je3CKXvIUHD4CABcVFcxf+Bsx+RYJLUKV31E+
s1lCS8aZgt7zC/6aTDRK/vAKJ8zMc3HeJC/9AGgbaBXNO+uglnHU/raBqehkaU/BTEqBoo5kV3Gf
U5/aGaPiEqL5n7ghEt18SOuW+O7GRt8CxxzRCXnqJcG/7ciiExFGlw1CtG4uYHuX+manPU8l/0bq
o6GRZukv7L0ZFpFHcfExr+VLzSQuVf7X+0x4jG3ADfsikUmqfMaLXegDCo7QZRRCU4zJcjqV+/95
ztqu1sQqzPbYSZLGrOKRkuvJOhAisK7vNuz3uqz9np1Z2MM89xwBtgwQsuN1tgqj410sap8CMRd8
qo4cIL2Tzwa8TIfh9dUkL/UiRi1fzZ/IiKbkuy1jHqkhp8RcePrCs3phxNgW8oHL0S5wgA46MydU
d82HuDDdtS46y6TYd9MSo1uCIFjrohtzLVbKtJ0n7XXbuSE+OsxYgG6HNd54Ou1qNcysTqXusSq9
rIcG+BPzk5eAdESGNiR9WquYFsOwfy9Wit9josWI1cEi4b3ydOS764DjBnNWim2+yPu23BS4yYFr
AxY60lut30vvXYFi/uG2FOmVLiJjT3P+v6nS9Bc6sTwCgvmPmq4p2ftNzzHnXS7zpDXAD2UmM/xo
Ts0onIJyQeFFvVs6oXmdcB6s59zd5NpZmZN/vFfaoVycYbB/Jib9xlgPA4aewxNIWvn3uuCVcYRe
YJ9481hh73CcRukMNfNuDuyalmP2e86TOhcP3g0idDnahXLAEvnB6wbhNHvO6U7cVjt336PSgthA
3QyySaRK5dxaSyNFVKVPnTUDmkvGznZw6KGT6HyZe1p045rVW2tgso88hJtDiCuJufqz2dwnpvhM
guMpRJeRQTwxZVLJODUKMBgfBr0b6pEUCPDU9jZ54R0UUCkCxot3AMpB0DWA9IPnxduc1pLWBFKy
uEGGo/c+fb89qraPG+qLVj+hBzpTlWsfDqfDccAlCLDcMHksLj9N4BR9lVMrPYqWQQAYMckHyCCX
7RsGLa9XdYDcLNHSDWnslwAAWH6JOm1GThgf8PkLUWA+a+ZqLOBL13lZJlQkH6fiqzmXAEfzVgDe
w3ltnG710Dse1gbsHVFlbdQSnW+OwDSpPfvbSsFr6x61OaoZFxh9KQN5plMk4S3s1wjCjliYXCbM
fq4iH6fQPWWphYXXn4HLhvZnLZe1ttR3Ow722uErnKk6wa7OoeVVyizhQURY/l69cxfPxPckyHTG
X2EBO/YMUkqGxc6S3gwGZ0DDXMzbKT4dXmBC+8JQMmUIMcXdGavYDfABFfGocejl+6QvEHb1zmjL
/h4rzmDuKbUEHxzaG2/gnDfNdeaMCd922x8uhi4sgjI/vS/2O5qrjNJu7W12RNNDFRadefftYVbb
Qmq1MO9jleOEn4qMXKpYFuCLY3tMXNFGl0aE+374lveN8eUfVe5d0sEusaaX2MfA+nrTEU86LImI
/HH7FibTQIo4p/a03DjdGAV33b1LF8kyPNWUjJ35Q4tntV01ewh1zW/Lcu6wt8qR5W8n0MNlLx+i
D2+Z7u9vMRO+qgxmDdXwtxkfOu0xZIFCVtBP7evHlmigzkU/9Fl+CzCBIEEodQ6PbjkZYY2D8HA5
v+4vQ4OKgtejWvb+3thC1f3QYn6iNfd5694Tn9DSgxe/4sdjaIYJx757k/wJSri7CPLlVAkYN7hD
rDr2YKjzbSsYiUXRZInfEtzzqKRSGduR1BpZ4SD18i19Nd9GSomd5tCEnjMDu2/kMzSVyGUezlIX
qZxN5jVGaFWzfW6j9vZ4J8zDS28f/aYnuYugB8slIGck4INyGTVUjwHcd1Ks4FL1LdAiteszl1ne
EPDgPd4yfU7DY53veXr3RUhBNvOHMAShJVnjwpM6yJrQNy2c+6H8Xuzy3oJOOHMpcq8aX53HuRL6
3Ju3a4HTNOLIfwsC7D57ca3LKjdARMYDWGH6B66pHkh7r2cAIYS1DyWr5b4PmCfuJooNfkkr2j5U
9eWgMUONZSPd7aGAwvuL4jrwOmpQleV6wb0FO36lK6TjIkjyb3KWJGn4oYP5DSXUr00g6OVg6DbW
NfbpvBW+IzHhvOl/nIglGu7tEU62oTg3s8/JxtJXZ93q+YP4bcwiCodcplAK0bdU0fjVL/W3h4cq
eQNz7mNsHKL5MbY9J88uz+G0s9r+zPq+ldc/BCS9qdJdHYqGdUmEGVdOKCbcADKU7YTpQ1dWvVhu
9bYphBO6qvW0xMeH7225XEXEXQmWDeJRlPu5g0mTji1mCsNnapNzVW1MNuyyW9SNUBd7gOnJOw3s
ymYOwvRRED4Aaads5Pl3rS9mUBWwZHhEwOF2tt3c0tcypn8FwlqBbIAmbu2xC2Lk+AoptEGkMIsE
PbAzInfM+W9QKfsTYTlMDWzHWg/T4xE+IUIy1qqoMsStLGa1hKJyd8tQ9L38EfAuCor7vmsQFMw4
PlKnqfFeeqhessYcTF5j3hKbXRvgcpKEwdVRocQaOefbY3nnIASrM8WsvfW9OQCbrYo4ryw+26E/
65ClH4OtLlK/xSws2riveWz/ZaSyVu1MHEbQzMLLnvzgLaezaVU+FEpEfmn28dYhI2nXWOECZA5G
+xhND2Fku/xeYEY9YuDDBLVoeDPfrWrsqDtKApSNKXZYq0yaCpa7Jz+y8z9Y3jcu14QgGwC6185d
WYlasmLpTG3wI1NTCvZLVGQWDLO9mkJi6D1LIwpX5IWKH3WXqPXQWuFdn/Kh3b5tBpBsLCJnvTBJ
Lb7pSZQhVCvLYUhVS7ESnD4OBsIhdhtGZMDfhIHR1jB/qxtsn0X4MyIq897Ae2FNU7Ja5yYpmv1Q
nj6dCgbVjTdOumIV6t74oXlYvSNb7RpdLLhHO/8U2J5EtAcBk3unKTPiptPtlWj7oVJbXPp8X5y9
2WtD5IgK0C1fy9mKfo9elxr8c6wf5Nxeu9nPLt9Y/5CSTKvQiHAPxk5ISojFTdc6+tfUonRRyL5a
dqYVN9WN5vagKFdR3MRHy4x2Z/SaRXyATj8o1b/b1QBUAQWDwSlmuQE34yiPtnLtUwPxWZYiXuIs
x7u8yC2VdWbSj45WaQPk34AaHzclrYy+FMjtz4mKSxcrn0QLOav0WRH5VprE1M5xvo3SzspqdfnJ
s9Svr8sB5hS01898hvuo0wRsar6dwtwtmnbTsXi/1kV7N1FlEsWtAfKgHMifrucuxzrKkoHYtkuv
N8mOuZ2a2zef76cPaiEqK1FfnKqbgx4mErfVQ27/GjN89yWJYtIw8htSxrXe3lyXF/7dIqBJJ5tM
KRBWKzYvJR1T4+DUvY4BcPhR57Y0Fcg7LSan/6pdLu4YpEjlNih+mA1F+QzvssreYnaRIhu6CSwh
aZjljq3iJPz0j6sf/A529fsJHh+2ULjcPvXEWwyZvC9rUnWeoiFUIvHIJomj9JXDoRWo63jguCyo
e99aYqzJapZ8SIjk/g70O1PqxsQSFb2bU9l41VB38o98Ca3iw6pYbYtJEaKfQEBXescLf5bCCJ4W
6CCiaA0WYnUPQ7Cbk6xoKgpIYIbANpU75I4ubZ6S+1915j+SIt9a0Af021t0vOyCyUaOn2n2aKrq
skpVKKmWX95PYMwzJE+rExqPnqK/ugm1HcLxhLw5JWqb9kVxo8PWLkgwAr8bGLBYuTj8QSlUZYvv
wvPAUnYwEtOy2F9whxAFl3R9sAhDM2cdzS8zeL/IUR3vxpq71cRxlLMmC368wF8rGgKXlN15mY4z
alV3vSbW+PW9JG/YpABAbtikVhF2sHaCxjjWfADGU7uX77bhRJazgssr/4WNiX/zPnsqm7EW0McJ
7iG8RkxZkfXf3ORyi8Ax1DK9gFR3sNT3N7ExhwVuFKMbYcT9Ci3n112eKUoffLu2ERDr5tL5nwGg
nFfyyn/NMzMGrGP1N6nNZVJVECEBWilyTbig3OkBgpsnkzLaTpIpG28IGwJAmdTp2Ykndd3QnKPL
32MAE/ZK0c5fZHOj+ZwBFa0WyipSpVVzaYp5CJTnzK+jzuZVZnpgY8tum1YODXsj13vBQ7uG749j
m3Jt3LWAmS5l/EcSQhE5xdeXUKH+c+7UBToSFJt42jg4xI8NBvskeJ8gS9IIaB+jYUlEK521LC59
adCWptfO0sXiRLY+9buwgarkdFzCSWpEy8fC4fXwo2WR4a2qY8bjNk7p65uRS1W+sMW8pSgvu4nP
Vpnws03GnIFetlUCTxMfQiDSN9nak4I7adYq24hK9cEpIr0XiiUO02NxeZHEc4eY4PFtrxqDtOkm
HXXjYxajoTKgq/klGO5pzQdgxnOOE7Hi0BBXnBDXiKmC5n5dDVB8jOv7w1RdZqQMYIL2iXWVj/XQ
0DERij/h3GcWxdSFIXlRbtn9asMC7RiSIwqVMIQ7ejK/2MvaLtZ1Z7ZevcuXE5PCf43jiZ+if82G
xrNog1gQwWG15lkhfdo0DeiI/5u8+hAuvK9W+L2nWr87Re8ntmIbx+rFpHhnPDbB6MLFmCXf9YY2
VTXZXcCOd+mNWesNljw+BkOLlPHG0mNg2DAhfWtsnsPRqj0HzBCLDWy2ku7BiAyps16YG9lIM/lC
vdLVm9mLn0V8ybhZ1zvaWrVOLMRp6I8AJTZcSV+y1B2fH1oeBwDP2ci4qGbM82Rm3B4TivtLlRhb
UKeU6pSAhnyDGj4Yk7O6ZJypB87GE+U5/nmQ7lRMwotzSI2FaFlnuQ0f0SjduHjM1JIew8PjVycU
qhQu8dHUcnIG8a+k/iFnNEj4t8NqEbj0NqfepgQjrQkXaV8ltlbrh75WKA9HFqMpU5eGWBsAZ1DG
h8vM4vWyRIGeVC1EFjc2614suW1x0zBsuICz0X1B1d6O6LiHaybfUZXRYQPPZfgxoqffhvSCnvZP
wH6vuN4kWlhgFkJ9JxlpXlJb1wnVBmyzvA8/52meks0Nra6O780SLXnC/Y0nfhXAB9WbXL7CfKkv
aJhjaxs0VQ1xEYFdgPicun5ifED56QmprztKoCndX+uXyn+z5hO5n83zMyeO1txks4gJU7P9Ox4M
nEVrDQx0Oyldmj21xxIpxmQVAuXMLLszPswKfEDoVN4aEubk0wIYKlHNJZ9zUeOpYtBjEwU08ky6
JEr5RDkGdCdZHR5xS2L60uSZlQjVig5KgZLgPCD275qlQ7HYjPuItf4C5ebri6yuTOkSnXx5yjnK
u2YGjsRSHNCz+mX3DHDBlkMNve3KvaBh853Y9UJSragIgnHR2q4AxTFwTJ9w0ahX2P8pPSexqbVL
uVWoL+kuPzx7Ov1XTla/kPr8vr/NQzbLJdRQzIH8hX/+VLrzo+is7+ac3PP9i6wu5/YY+bmMVgZT
iEDmU8ZTEAuEt6ntNjAY1FAPL0lU5jNyxCf0Hi6PRHRfVX0rCE25JTHzQfS7A2BwpN9fz8fJ1rN7
Tdz6BjizyRHn+hoVCTp4e6sOOHezxJsyaAkLAR6+iWPmYCK3aIyhpvqu9h8t+mLjTXgm7K+DYhQw
r51SgH2CYD5YApnoQMzU1S9o5MIAn0UvVsZ42CAWNOWyVuT90qgoHPRg3dwHIqAzlQmkHxNNPmjP
c79X5uWJwZt0Wl4NBkhly0ppqz/XQCF4Hcb2/V00nDqq2XJ/JJP/BkT2N5yi8YrhD0UvEJBvnB5I
fSsZ3QGmKvH0z/01dUtEisIZ2ZjVYO2K/ats7Am1zeUZDYCwzU/HZOPdq2tIkQg5RrEti7/IsUvE
6YV8GY3sAXPgSFt9JqMtb8lNPRGy/hhA7UEun/PfbeHDRb7sRs8+LbO4pY1NaJG4Bv9e9zqfv2Py
C4caJsE81KWfJ2pZKvDrSc1lkwwjpBFAIeUuzI+rTM3QH9TsfLHTAPwmAMVWgs8D6YPm0fnW8VuD
IuH+izp3Tj3/ZFo7GCLgRkTZil3AWx6lXghCE/moVtEqC3t8Rnav+SmrbGetRHFILsbTD/n1W569
gWmbrOTgZERHTQJQSv9Ge0EBCbYXC/wEOkFUKRpdrzzuALx6JPNC65R5w+tvbBdUOhNxGcP0C8bL
m6MbFGUg7Ct/J9COWTz+zs2uU9kgXnD2ob0dAWTIhtAzra561pBXbr3uN+aEbqwwOmFTDrm2cU6p
XYawpN8HkvrfAX37wFmfPkSo7PGYgppHyQ8zDqwXRhk015LkM9r3D/0Mc1Hcw3v1Cuu+MTE/ajJv
BepwxN3rgGWgONGThuv5tRjd9DhoUVtzGhmKT+OEBcWTeh+dJIQRwopb4iR7QkOQEejicPPfo4aO
YpUAUNJ8xhsoD1B8+nqaEWZjmzcD3Z7Iwc/uFedqzSN1HpF5JZo7nbPCnp+pHVemKD6IwBcYA4b9
b7ZxobIJH8Gh2M4xoDOeyJ9Hw29NI4S8BMl+KtslUdLWB1gFKobDlr9OCbrfcBk+q0vRsPVxIjY3
dMH7SqZRxICwIKKDNPQ5Ncm7i8qhliJpqnnmIek6FPCLlwnRZHVcFsm7ttpqVC0yFzmC+HWTTJEw
uLz3PwVik+FxQpE8gPXk5uwUkENwXim/S5PUUWktd6opx522OWN1M5wYnZUVdRRZdsyzFTm5u91o
A/fuGK4KixVHNwkck6bF1BKB390SvEa0NaL9Xl9rfjfqxaxoE+rNS9MhNLCoOmOPLtxXan/SOdWu
bMvNNbtLrjaBMa8G0cVny0PZO6gZXWvXDoYPG9WcRBeqt37DQOi/vuDpSjZzOCd6fxr2CDdAEm4n
nug1ZesGp1X+iLUnaLqLbLVyfquM2BZFQvbIDCaGQ1vZ99fjCm+kXog1aKgUef2loefIJsdjv1M2
GJxIZwUzW2AfWefVaOykJRpoyNCjavtTI/GBRux/ehHkaYhaQU8jXQk7J9Jv+kANzhGHkVP9hBra
+PyVDMpIOuMpCSIV8RC51bE3HrR5mQpVHSldhJQfYNNh26gSAEgyIijUF5Z3VBEsq37T/I1ER6u1
1Mu9MrdNw6iODpWj+fmkl325hFdT0rljIyUt9zi+/SVd+7kzVwXGl/toi4PMx0CNVuGSIri0yIpI
uXqGabnpyAXkQKdhVVw1imX+joJYFOxc/i711qeHBnqxLUBIOyKI9sjbsEggELqypYcZBM0sqBzc
2gmTtHFiYtqfTdGu4fnVNoaC1zn6mKKPVaZgE3h02LJsloxfifAeBdrAFKsPizFNyG0ex6S+sWv3
yQ+XGgN+Cbp8oZSIE63P/GKpCDftm3hD2elKa4cx91P34z/KfulDks8K0LkoB6x09z1/QYivime3
5CBOhfPSJcwnL118idL6KTtcSbCP56KQ3socaPRvJRvDrRBgA8hH84vSfxwNzgrnleNupP09VNq3
ioCvz0l2u7aUoagg5tWFcU0w4SEcgOBtbd8VKN1IkxeEAI7xx3EC0p8jAPdy9X+BXG+CgGAHoomm
hU1CzjaF8ZTP3dFdSW0gdTzAb48ErR63HS6Y277uTdJkF1GX63XZtTrjNoZXZLrO2HtXqYLZJYn1
QxXRPiZ5yvK5D/Wvx3uFMD6WmVyRXh95q1KzIyFTmNKUoj1jyR1q3aZQYLIZZA7VCTZG8OJUwcJm
IZxDWo9rJJULXD6tT7hXx7NaHemZ+Nhi9LoPE87qAY8PJrYRLusprFluevPiPtUgRe6foYDt4tN+
mo/GooRQXNP7+69mz6aRaFRojvgm5EIhkArjejodKvT6ChZhhEJr22HNw2hsI8SDlVWf7Ii0WBdA
JoEHflncWvet7bv7fw8po4PYf1tqvRvr2412R9+l5vHtsxk4T3CComF8bpt+52769d7djMmYwjrQ
6BBOC/R5es/IYlFhlh1xzwCNDgu3FE38csy0YS2bGNM5GLrE3DmPzDCLx9FRcohlH1YIRxOHlWBx
LtO/C/p1W/kNvR5F0bgnUaEC4Ynm9gcTKztBLPWoRiroRROS2HiZLAhmnw1tolCRJcHMvhsfDwIA
/fVVFiylm24rZ3OmQFBKhYHpO1rn4cKnqgJipqIas3cREnYIwlbAndVJZtMaY1wE7gx89reA9qEQ
Jfz3wS9T2zm9e5Vy73FCAtU1iYRTMYbs+8Z5zv0CD7kVWzadfpB9Vug40K3Sccm/ALWd0zEzvGow
+kC+sPW6P2aPCAAddkcjFMAFi7N+qzsJQjqmJshFZuzqJTAXcxrFPj1qVyWUMOQjRX2EPxYdE9I9
L/8DEBzONshgnIlsC6wioku8JL4oiqGqGGUrZNGR/xsNbTSmWvxcq9LBiUJ6laHf/4FULyeOTmDZ
KsVHu2N9Ga29UC+k6+gA7qx4cHJVwlcs+tUpxDaMBKBD4QSxjGKzpstm1jt0ueH/p7I1POlLYohL
o/jYsGd75YOp7uDI7tD1CQ5giianrvtjAKw/06cjaxlWflLuzix3AO+h+792I+GLEX3nhnOnMJsV
VsplIxAZZuSW4sCtHsM5mRzbUFHWLir1XiMCu1YhNQz25YY63/J/L3EFsTNMf4zve4AKzLuEBlqt
DiZJSMyCjAYBbiwo75Oh5O9h3rPcNogAgZndnSdGgbOceN1Mi89u+yM2bFcPDIL6wHdMyhwBL6bU
zi+Av6Q5hLIzcCsySvy8vfB+A/JI5W9HMGN8xn2utu4pwy7ShSfZ5IokLI8VE4YBMzoypnVhhHkx
IeESFFe36uldlElPLmwFGty64foYFVFeO0/e7m/T4J9UWOefehoPU8U7QVewL58aJanN0AaJX5zA
AHmOiR1drPg4yoHtO4f0bXMuxhbx4ou9OUjvdeQSuR/uWDv1Stc6sGwBndJFqUi0HCSKCujYauyg
0Xly83JF256VS6epn1snksTJEywnM5qe7izC9LuPyhe9i9Bcaqr86aDTBglhq7xYJKzwfXYqEA3f
ONGfBdRgNM9+j9lzMDvWxG+mxVcFQ4UL/KslmjHsOJJtMOVjec2JSFF4ZVgOhxo9LPHhbNvWuRWh
P6OLtmmgzQVJ2Qaa8vby6dvV0YP7aDJpMRFANbRQL0C2fxsjWM5Qi/JPqaz4NO0+Z7d1HHpqpTR0
jgrBDW9b9vthyL4ymk+g73bFugOQL3LDtjjxP6x5uAEY0sjp5WqUVdpg9j0RAgPNe96BLcJPWJ7J
rA4C1addVCXy8XzUPTmaURCZ05mMC1O88T2W96RkhPMuIABJbvRYRCwUcJEct0tbtmt6uWQhRO7N
gq24/hm/yPfWVkN9M5/zFPky4yZRRei3t4PhoB1v5dHSn/PrwHAXXKlTZsSn9C/WLaO2DCKKKxlE
petnN/0ToKVJwIk7jJ40Rxlss1vtq73jnMJEaH5FtgQUnbU4cWcVI6BMv5lQiEj0UsONaxHTUPZ9
Hf9VKNx14vozo3qvjGr9DWRt+2vLWY/TnEYFla/OXj2lVYAk8iHD8ZfHDbdvLC03fmdkqFFxJpiX
Xt+4yLY2vZqIddirI0JUJz6WqKe/R3aSTiSKapRDjVtGAtOjtK/KoDKpfu+DgaxzmQU+Jxx7EaqQ
8s8SL5OeofdsumJUNEIH2RiM+zeS43ianz/p7+BS8FeBmnpz+NYfOTLYPg8Q3fHfX6MKCmFt3126
kyKZOhPelTfrdFYbunU29p8kZ1bfc338JHPPQc4g0WHtpfC5ADynujl25Mhhg6xcTqESCLWp3fel
DFCtUGWmMHPUHlEBgHNbZpgM8wMa9bLRwZizRwW3siUV949OcYXePZleX9yfnHI8Q5Z9ib1pe13q
i2tbTgxWfDr60290bEbsuQQlnz/UcW+qmqEi85V08BuaXc2PQ4OvWzHaCXyV8faAAwxa26lC08Ju
90afdnZXQkf+w2DBmHKoMWCcT2EFkNAEJHp2Sw1tCY4WspW8zTRIQVZ1WzvlIyZ9F+PkENKThio4
Ko+aMrCF9Bj6xRp8vBlOexH+tZ0StHdTGShS4Pb+4Ffd0cWqJj+SpB9xKne5ue1ZLmBwWgz/kuvP
fY6a53iaZ2Id1GYvYAPuxekMZ98pAYMZZYVNeMAxMvZkF8GDBJQby5lJoaFE4azsRoIKa/I/f8V6
qb8631l9FIZKv5ld3WVBUrfhfV183Kva11WE0VDH+xHy2TECgtvUq2pFJR51CxTQR8Q87/JGcQjd
woj35wyqFMzfVjh/HxB6iM9dMMfduaYAlzE68bEGJSQhL3df0l2JfSSs88MPUJC/vn7AQSuig00R
D18W4THBRlHBSWFmH7J2RXJ7TTQhXGUAYlP5I6x2UcPFx8QLrRQWY6a80RZa1e53eabODnEUTa/i
gun20OJWqnLqses1je7Tj3ttALFmgYsDgQiLnqGHQcjY/gHFkHMkwpTxuKJzCR6g4F9bt9By5UV1
EyTqZzHbwYro6a0F630+p/t4ejJLSH+KmgjoXj4PHnyy76VzyjnrT+mL7Y7y+Y7BlxsN7DKK36eb
r/PlTBKgC7pwYttiDswklrWVwL7qKqJ0ARIaozwxjh2QUG60h+iREzNNhPJ2SUzFcfgltdtfQmRR
B71MHb1McxJu2deCzIoJO+SvpBlr+quZT+e+nPvBJpa8dLXvkpI1LfGX7dsMhsetOlfc5S38k3DK
S8XcHgpmhpjSnNVTHmEGNvWcMsJ/jruDnyaq9hzdIlu/Y6w7jc8bgf3FGwF+TBSByNrEKyUYu261
CXXUh+rseIsuP38Azu988tuHa8R5sgvasfKfacoS5NKVPbwJJZ71biow2CBq7AYxobthcYnXdhH+
ySJ1Bn3/SqOzvfEDZdASf4JyEhv7uW7hQuXbBt49I2BBcbii94kt68O3iuO3bUsuqjuBmslSVEcF
kWyDJdLfpRliJFiG4jS9+aS8LiPooM5GLC/5ppjvdZexGuwUHRBBy31Xut5lV7sQDtt0JeDx4R5/
PFRuKZyaFZJbQl4F+ubLuLkw7Lx+mMPTb9+63KjpV3X6F8rhKUFYA1lkV7bJNPIQDI0dJoPYdErS
olinMQX4xe3ZtrMKLmvoa2DgSfGjY/G8H+ellGcHXicLikAyxaGfTwLqeote4hX0EYW9kxwztUPC
RaZbZTAyBgdDv8fkzoOUQDY52TMRrkbYtLPQRXZKqRREeHj7W3Fzan3EZYe8aRZ1VWEwNT9Druek
KE+h/HYows6as911A24P0gtws3egyDvei9HFJKoA4p7Ou3bJCaSGkGPWo2fek/VAFozU15p55Mob
BAJ3/sZ3kDNO+WcJpaFJ1Z4zYHTPsmaeKfftpJpMznoTE0SggxxBm4vDt/AG79I728A84MNbjZ2b
2MHg4eXPLnFhoZRi5j9KtIlW7dKH/4xOxzGQqybDI6Lt1Pe6ozbAXIrIk6UZCaMruM84slBizd0T
0b5wNCtZ+V5Dg9q0b7S8KLYsecUg430GEj0n8KzVZXSuO9Owk56rqHmhBRnkZKGhJBSUm82lOh3O
OGBP5hMmtjUA19dl2LVWYxbSvcVrZAb+bCh4dCDyVNIM0ZRfNNKrfmxigHpRKDhuHTL1BcQKcxeE
9jWad2GO47lu9RV8hAc1ircW+AQjrDufWjH518EEA5LvWJ8+ix+U7/MapXDn4H7EWHUW4/FDy8aV
awqw+d/dlZiZN+r5SQ/QEdpiMJrsE0/nXMY1x+smpZbVH+BPO+Sd6oKLI56VWtoZoAXsA+XQSazE
IfPbEBf6/V/BRsl++6MD+qe4tHtPvPShoN4HIp1nIJJd+qoV6gD8tgBnwFi6VvJShIEz6O5mZ2DA
OjOU8H1MbCHPJgLfImAzy10ZLbfS4bswDabL4n8PWH5seqQbKt7eL6skhBG8z7TGUAJGmsemuOs3
4CRbDqbtcncnZmvema48UAjFpjsJXhqpzUXspXLZkDz/v9OSf/s1V5d9/lj1asHZSze+fGWcH3pW
pQbeIQGgLDXo/eLxlC0Z1xVcqGnVNfiORaGk9PTlMdwosWtMlSd7mkxG1GdCsHDEqrle3SO2NuO2
cB/Zx2MsHOoXy+dfNMNJ/2WHBCEaK5IJimv0HYbgfG6QExRUQbNCWf2iU1t1EnpPjVG5R8wXmkWK
hDdK2S7rkfZK5GKGE3meIywq2uD0LKbx28gVPnbpIZa+P36qSekXJXnN37dOzkt1QeebzCyrlTWq
iunE9wF7HufnLPgOc7v/2NqU22ydvlHpWGJvGa3IVGCOGPttsaBl6YTpwjfxVKJkNVuuVvxBwof0
UirqBQTijOKaN/615aTj3aUUhuntuhOOhBXCIxI1356IdJziZTYrqdgn96ULQB9rtwLG3o46LRzn
byJrl58imq6/+CcDuf7AK6SSljtzM4eH4O1Z9EKPap1oKaz0+3jzraHtyN5NrRh9YerGqlnqkZb4
kH8Ou8kuVoJxr8kKvWieliRXjiYJlVvPk+CZsxyb+MoZdDbjGeOiYzID5cMlGKPXHvSjLtL25MBo
83oU0DHnmRCGY4V35TBHKWwCWqqdeu3qBG3OFQN4/btLnZ8D0ZqGUYaSkmLWvfaS4ncI4kg26C6U
OW2XN62h+Bg9P6QB2tGqgYjq2RlthiqGtL+KBpLPG+Fsw95D+zshl9oT5D9wBbM3Ho2azS8LZ4Fl
B0RFYOFQgs5RaGraQ695U/1PvtWTBKxa54AlPcDNWuDuIaZXRfi9k6JcE4NgbJ3pLJOcB0JBm1Jm
gqykiXMSCqwi04qrbGoxLS7S1EWCOLcG7vY/cNHUWst8Fvguzj0i8389Xl1ih9X3zXYKwfzMYpjm
fnKfS/nz8u2OlBmUJlieWmaeytSwXMLScI4qeooT7ez+8CwKPBcheGPq1n4faR3Cw0b5POdOUc3L
Jf98WeB9a6rByLnHVk/kJx/DlcwdlwWli4uwHrmKzr4JJpmy/PyFHiQWBO3uFoqhOaw8coXSpPcq
rhgMqu09V18kCjW1T1XLDuKhIpBiTLiZawATRj5+UxrntTFm+BSPfhAprJIciLarJpi8deoeY9rz
F11V00PWx2aMTfdJDdz/dfpNQhCZoDaYSIfREYFZHh7SgAY01SZGAxl6kg1WNRWmidNKfk9HvQWn
ntF5EVsxVO91kIQmKz/zQ+WAkqS7BbE4jMfqLSKqffBU4ZcE0UXfpfItm/NnXVRD2Wvo3R7fIoVs
9nbvEmihvECkWkXMOSgl54VJC4ccd8gKTqDC/uWhwCprJ0N8Re9dnO6tXELrx8MnSuWyS+psjT3k
wRmg8buB8i/rPF1bXP0H37YGS5j+AUbvmHGqgfcYVUu2SP/PuF8H8cK7sx9g6tH0C0U9RWASs6zc
/qjkpQWjvuEcGgEqFN7WuAuYVAlmJZV0Njfmzcro/5XsT3wBV+qp+O92SOtGUAucjQ+7WzuKOdZ+
qS+JF4LNTVt9pYYgBQffIT0bMCwhcItrwYu/iAAzHLPnP2V0le6T5V8TJHi9lrxopK19KrkYjXYU
trJCctopobcXKrQJmK9aipgQvZBpzMYwWM55UiaGZaECwHwirZseHYjCdO8pFN8fdXUpvLHJvkIL
Nb6g2JUXD5JpjaBHTzz1Oz2aHkIHklvxjq00PY7smd2ZSYxFl+XtO9E7S3y3iCLgJuG86fWDU49Y
8k0p2RxzqzCGoqh608xCeAifHmVwU3m166GNULjJ9/vQI+bsC2G0mRQycetNHIyeW19+wvqSoB1S
rZH5qBYIjHz7RzHW+TQMGU4wkTRz7BbcIW6pvhu443E/lHkflNcGNubXJrZjwPn081lw+kuTxkjQ
o/rpJPCXXRKGHOuwT7C/6/wnR5yczfkhw3JncyMePv8iEpBIM6TC0vLAw4bKPWEFwJTiKH+C3j0/
/jWiqnU0WqgpAJwLYvAgM/Ms/X0hlV6namg08afkiLL4ap2UlntppYa2jCyp71c2M5wxkTj0OvBb
lbMbs/qaXDHUgPyDf85H74WIfkrmRgE0aj4YtOZ4viiEpapH17VSFS34qmcB6C9V5Eei/75Iagt9
kW3D9YDOq0Fa6jaWQnUSArQSYN+KqsRavsDuiZchJ8p3lbAn7t+ihyjEX5sUs7WCiYEzK22m8ba4
C5vERIT6DDO7bZgdUI2qWZzYEh1iSe3HVTQWDWQldNTuzsDSFbEy9fCnxMbc/6fmSs2Znfeq+ZB3
MIIyblOWGN/90fspq/gOAZGg0dbPWqFVVc+CXpyikZJv52JaZZUnq7iHBjO/sryFifg6m5Q9GxZV
hhFPXRaHGJf0ZEykr6ON5O5PA06JqDpirA33ExL7ByTbAZTfkCny2jrF5P+/26JkymX6N3NvbQig
JvzUThdGHQbRsZHFWd6A25btVDe4nInDnpXZViaVL5lzIMSFFrRXFXJX2avP2yMYIEx+tEYWACW/
gqLgmuQbIYo7ZnKu6GPZ2oZbOxc+EDo7XbEAi3FJD7lowiMXQuKyhj7T36C7rdKiP93msygxqE44
WXmrKZkpCKKChr4TgOiQRflAZCammAmIpHvDETmYFgIGWLiqjqQlEc2BVIFBqbJCmbuUVljbtnOW
CLKkbUpxI4bab5tIP+zCPoXMDL7CePATW4Nsnt2dWbeKIiYDmAlamVb2XzBZgN08CU9uN/I3HfP1
s5qPfrwcS2hoVlIpRZdiuJknpI/VjZBUw9rAEyVULnEmrKD89XSknHgWldm1rH3H6D/RX0S/2oDV
OQ2nTivj7JYtGQPUevewnArcCsAtV8zMrkvxiL40H9qB1Y05FAmOmI4rukxEBJwbds2rcgcJHgxt
CHexzVQhEOFClUp7bP1pfT9gtEzMpZnsLBhCwdAP39w76qjW2zcpzobMM7ucbYP+UgqvvJOH6N8w
0DGETdNsPyqU9HcmT4H9aG5qFKTj0lYNMk20+t2ZXVbe3VXx1vIkcmb3DhdBmFXldRT1AKSOMaXC
THkQZNXGXrCSjZw3Zd3YCWgXowl/6BbN17qPyFx5oGvwSq6kwQAQRhVQL2FbQCdq4gxR5ojUQQE/
Hz58D5yUxGAxZzJJW3scOMyAvhPKHEcksPT99vQZd/djLsUHHdqOpyPlXQbI4niWSkZqPhDP/hA8
8L1En4JU5rWlL74/3CKsa390rvW0HtwNqQD3GlEaBnvjufQ2PeAHeqDzGXu5d+Mo0f6S4dNppRdZ
yX39tKuyGmLcL8bSL3JqHpAZbX8fohQo8YRGrXB8+a/LcKnMnaLw66lU6jSuyWDDR09lt91Aku28
OV3lSINKC7BixAxoLpvStThOHI2DPBHpN33t94+GBEF0jIQuOOaNx/amabCZnHLtzbNnIXjmrTIh
A8raSXv5Biy1XxlxJ11146jgvjEOwLBhf5pZ9zdTM62l+WLEqILR7XRK+guCIWhlIAw7x7r8xvHV
p8i8GN7Y5pdUpda4XHq+IbwNDqGjcMvuxxrR06gH7QdsNIA2PiY4yMyMPyBag42JwLsM1oG/swFX
G762fq0/hUr2W/+0/D26K7cw9QLend7+CibHQSgc9M2f7PuJIJUNWL7NtZR4bR8UHeRleWPA/CaY
zXABQQPanY9SlEsb8WOVgkcz7NYXFCGwbwql7vec/VuFWaDdDrraE8OGtoK7J7oz2FEFpfMig3dV
KAaEDBrS+uYukDF+/82GTmJ/gQovxOjgwe7dhG2WJqRjFjrXm2l7P/fO7ZMIt7hr7NBlPZVEePaq
4VqCzFb31FQu9q0LxwQyRM6DR7WNcsKA4e8De7O8gJzMFFFsLRf/XKwKqCEGoPpugrfM5eEf4yo3
Ac3VtxzBzTz8eakjD0UGGWgi+OVRxkFbTh6O0/5VNngRvo8z9mWkgXwAfTfOI3vAC+tGvQeN4dMp
F11H/bxwosvbhI+M/0XbvDs53Lv/4yn0DzswTj4phq1jiFvKnEEl8vVAIOZWG1Qvik494NTf2MTV
ZJDguunT5oOmAcDjj9ym9Pue16r/P8TW5XvCvdzP/DEXbJ8CKJDkshPUT3zmfTV5whJcToq8g1fJ
Kqi8/MT+ot4QJXHr31BotkO7/a//Dpusjj3E2K6ewizDDixXkKAT3Lxv0I2TvRpAWqiONT+cN6hj
/6rNER7bfRAM937vv1WutpFW8zcnJKHSkMpyqFzhsEepsiHq5gnlyyDhgG3NTpfZ4oi2evShcIOK
qrfDdVg21HmyAs+eV3nQMW8nrgA9dw2b0AMSXmK+zjv0FGnAhMV+MjTejtQMfAwoTwELfOqj2uWg
V611JYIC4YvE+EcgZlsUZtIerPyQRgpRFoEc7Fl0Wxxlit9JCichoPaCzTxgcqJJe0QhiMMZ/r3E
Ze7Ttjq8Ykzb6B+ek8VCrrxt7Iplgd5yeBMt0Wb1oYkv54SLGL6l6/oXMv3AqZZdbfaik/R1RdEV
yWw/F8CUPgTV/fipHvIz4gVvkL1JXd51u8YVD4lSq09xC+cNQtlUIz8S+5Il4zbnROZlBphwL5ZR
QGW1tTX3sQP4ObW6sBrlbDHuACYafLd7R/hPdLd0aC5jShHCXOI7xqonNojcOZiDBxYfGBuhu4Gr
Xi2fjo2smfS/ZBomev3gGRk+o1J7lHE+2+PtGADqJ9rm5NCh/G2i1U4rKaiHYXQ0a6U221vrVBLX
Gc9NlRRyYthFmc0szrp6fKNeEi0AZ27XOsPOUBbFqm+F1kTzMDcrJdbUOVgd7Lz+6VNT4ei0XO18
wc0hPPHpowMCvLxKy9fhtHlwbLNe0gjliwQCeZh7berv8Amv57w0BqPO20rn/TTncM6ODx8nP5TO
abjEOnkm+8vPpBZolQOFl2IaKh41vh5ZRU/XgXXlFewVTdMpjoqsT/bm9uBQl0b2E4tkzjz15Qf0
laxLgI6tOR4xYNulX0o1U0EnpDVpmGxMpz/fVmAy1ktJQU6sykCi9zDMv+4OHn5OlURA5RjhIWaN
DPUObTPzY7PPWxCqxNT6jtz7uSxsswNWYnhUdr4E660Wxvu58QtzKtsutXUMgJv5vDG2ycQ3A+gJ
vFHyke0pzycI0g03izBKlgMl4gi2wcS+LynF/bR0dTCAhye82O0duH05QbaNsptcq86EegNdiPAX
rKJPHC5TTqi4CZl3DfbidITvK8P1G0qhwAB5SgMdQhb3sa0SIFYTW/o/q3D5dG+5A+CWX9Uk2ufk
na8xwfx8okASvWd8ZmKVrXE4AAyYFhlYiqKbJSQw4PU3wwoQIAgFkIS2W0cI3S0Nw+CK0eqfBH5A
/bWR/MS5UtoZXz4gdE7QwVOF6NB/RSySMaxoLmtaeqj1258eWCz31UKdlmsBylG7Mb4WR/lrwCQd
mvxAsKOUidNim9+y+UfrQX/YF23cCcA3Jb95lvjQifEbm3IE7UeTazy1tk8M4e/IBYsHtXSZgqP0
wvIum0qb3KZJv8inZ0x1+uvNEO9sCmJNsH7D4j8kWWzLMBTclkRY838eECsTSB1KtbqeKtqdyPg7
4ctZdDnIS9jY5hmcChNKbrPzWMtR6XbeAIRowQdpmtwV/3WtqEGSVwVOFeSJ47bw3Ur+ZXfmJj+q
IM4rb4IYLGVBeF45knhK0LtXIlVj0PDuMl6vkN04ANZM6A++ym7IQhIEe4DJWRDbqrElU2cSWE40
9rUgkis4uQ6N+XydQqC0fSJbefA1eBlIpTZmc6oHMGuRIFpdgoCGhpksb/2kIHvxiNWF+2r3pwsN
tpZHZogIl1Ag2BVM8OgHGkrNEVNke25/qsHmHYxryT7eIUv0ZHHFmp5fOoilCEFIAHr3UFQYLpAQ
mzpr3+KF2YAICxdXV5LAwoxxiAOHqRTKWoYYVERCXYoyzGMAHlPsTxqA8/y8JLZW2VBnG68UfVhw
4MgX4XXF1JpiLMtCsi7bEKbvZ0H0vDVNK6Wvzwn2j2Qs6ilpTzTKUa1bKhYfIC9jeclrMqV67Bm9
gW0c4gkPaIhFWT+Q0sZACJiuCmi02g0aGcBw4TRMZ1s9l6AfeiPzaDOSWGJxDGi19YiIrXJThio4
/Pj0ihoUE4/6hTaMeRSG19uCT7t9AOhs9YtxMbP20Yoy4RE+QeWGoAhqKEHUYQ5VToCBrFXeiEqj
+sDqEgrSIgTAoVphsQxH0EU05TjjMTifZT2AGldwMQdR4JzYmawYRfyjTJe7S6VD1415WjPZZ7kE
B08EEEgLpyjwg4TKRWlU5vqTETaTm07mE6dBaC9gZweQqV43Lj2pt6JV+yK46R7b1cDTwsj/QoR5
k0hy8p67HTNwLI3ElLanKTlogFBjjFAl6LbC+5viOi9p3PxkJkbRzwopsBirtRvou+fcoaoXEnWU
STQ7pXPXBNiQ50dZGFs86sAyChJuzdbLOr4BXehv6hAYdNU+onZ5YZJFm2yy0PTsbk3EzrO8eRQF
zRxydmPxX80uiTe5fbaV9YVOxNys/Ua12BPc5HuDjTvvggytDzuj8Z0FCZtQqHaVM/lmpEL30xQY
GyNRqAQtXJUCF7+WWYLrjSnco2q+5yHNeruS1T6LDsxaV4uF1EQk8e4qcdQpvMB4Dplouj7lROd+
xoAiPPLhlRC9RVsoDGphGuA4AX+ovi6M5Cx48Fk9B96m9ToDfPkcVc5JdQsUMeXfBRHSKDWY36Fl
pUBN7COTZmqlE+gMK3LiR9heACRUvrQt5U5mJaATNUVloWBtHOzfkLiQNCAzNgPLugtfdLO04r11
fSh2CZs0YNhiHJTb0z3brqHqPr0Sdl3OOXEFVctfVlewpdktpBzPlApEtMzndS581PIku5QITZDe
/CvcF3ksaE7KVMZUWI2FddLMk6lyBWxMEc2deTkopoG3du5T6HKNmDxbJffAVkH3HO5V7F37JECe
BS4g1U1viKbUppi1lYWz30LRhBhkFxbVAZYVEmzhxGKu6pushfyYXDlua9pQfp1ZPqXIT0tI5xHf
Hp1ta05b0vXKTG3PoLysCw6LZqqjPXY8tFW6+deqLAHjmMcNhnDCNgHk/2ZdR9MZo0l+pT8XrMPJ
IItb25+JALL3e/WtynZSQ+baP0sFev5rPstPRSy0Ee9qSsHQ2v/W3q6M4nzgxGRKTJjv6fZCkbuI
f7eRMqLhxtumDCpeffpYyeBvV9Zv7t8DX5/WOfvLEtdBLJ6xIfjJCB4Mxot6G7q8azBwbsaoMIGu
TlQVoJG/HDmJEqEC4TV6vElDOlFRV44fNXRdqMBp5RtUjO7U5pnvpCOD58OSs/OzgCoXI9WAC9Gj
JRb0MfNETuGDapaxC8h8at4dCwcELTpm1hF//1iNV2+mBQkO4IRlEcSGQSMkzOA2nh56vvvU+tOr
LYjQFphbo/92Llk76N4UhAP8QLIDoeDy9RBQWyU+APb8nSS9Op8HT6PS/PWfDyCVBg+sWASTpA1O
Y/9R+2eVUBQAimmIxE+F68WaJSm47c+tvZsHwZal6WysJXAjl5BFR1QCyifSAQaS/qL1USIOXIf3
2ZgNrTK6RfwkUhDLDlpoujNZWCoz8nvu/F6/+sLz+p17Sw4pF/ZL6jsWN3vdjwz7xesTgwNsHAD1
F+J/mKhqQ1a0Y6BVKox58Q5MXiGahU8hVlG2cF2+2FG5N68JSybe/EBzcT4M2QS1tM0uymfDWyjS
aYcC8IEDVly5GoAVPxqN7yDdN+89Jk/JowJJsUmk3vdMQG/zuoW3bEJikVX+9KIMtqcGVNTNbxpm
JtvTuvUBGiKIBo9/r4pf/DazpILZKd1seTEYjYdhOIEnenfi8kS0Um3zxifk9xLBmcJoyLiQpWoY
1Uwt/HxV004HB4hyEr8E3oGqHJy0xTGquFWTMjoPwxprtfVfv4TavddQAvFLNG0URsxMRze8awgp
rOP/H82GbpPq5agWepGmE4/znb20nELkuwJbp1hyNwZFoViEJyWxxCrpb3c74MMI+8iFNPEyWoBJ
h8MZTWb2QwaTMuR4zMindIYeTbeR8cpB5QdiMVxEEaoRYHQEfq2tenuEwuK7n2c+uTUi/wSLoH7C
KlK8OIQTi6U4XG/hYMt5sPxZkd1z4NYPtGgwt6xMBRtinCFGVJg4hqjGpZajli7H9wOzkJElfa35
5PKOaOfuWld6/zGvIE5m+s/ABFvRzfqCESva8nUQWEl231RKFyuuy0bSAA7Ty/QQoScya8NOxsnD
oA3nHtwg1tSJRQCcLWYBKMIjE1P2tt6xRxq++1UPt4oO61z+YlWMaoksgRBvysBYKe2X2V/FEHkq
A7oqiT7DoJLqLV2fsLILAxtgt7Hyf0+D1kAX4OswEezlTyicWrBgk+ECib6zz8g3L9m8Hb2RRlN6
RuvR+kSdr0qOYSsPVRXgh66f1BGD9nhZp6iCq0pTWuSZaW3cd0s5gVNTAcOYtcYlciXypJX8jUi2
TVS1J9hthHtNORlzKLqC1FpwdYtRh3iIvrVXdu28GP7ZGAlYBDGfX+ofT//gezHP3IQ3NpdCNCcI
AOkGkDfBtcO0DcLpcGeRi6wJYf/6hpL+zSwr70IDcmd+lhL1UsYlL0V2gYUa7fAlMDkHC7t3Oyvs
UBvqR4z3UGT/U3U6HRFIFzUf9l4lBaFc/igwbEgTFJlr1vSxz6qprYDKzH511vvGa4OwfR+DQP0C
Y97oY/D7+1sFV5QGY4MwcTAhld/spHq/ud5F9vKDSB6ZNl7H0Ew7F1LXmiXh/fruCF4pV8bBV8To
FF5TjuFEmqTBgggF5CteNP9oxxL049jk9Psp+4/hdVwI0r9WTg6Q9BdK59mzTDHAlGfWC3f7SBgZ
KJI5AFIvJ6cK91YwEw8XaMAQdMCg+IsplNnTO+E1ZsN3ruOxq5loQ34QbwIV0B8dzrsFWvtg9HLu
FbvlWPjQuJVDBe26JYd/FlaahIowVHyiF5NMqnyd3BvP6hnp+dGFDbIMfKO+70mj/vfGB77JWocT
0f/INMyiwL3IRTjRHDSJGdzz9xR6r7FX1Isf0SG+5G9u5mS+LjEBhY+lxx0OBFcqn63xZYqLdY17
bPMblzPlrgp2o7aXAatYM2CJkBqyc/xdBb6eqr5GoUudOF9GxFa7i72fruKhTa4Zwib9gX2e77+n
TPYl2hzG0PS7IK2k+3tO9jiKtW+NKw86tx2ZI3jgLFLByMg48fqBePrASA/CYpBLKp5MbF0dKnmx
tTbMa6G84a1nR+iC/pLkSGyBiN4edKh15lTMX/8y2HeN7TnE0Y415GtbKnI9ypYvzjsc1ZZj2wyL
7htW2t0lSnBKk7chrZzBLxl0Qib50DZLKB9iDDJW0LCtVNfCOCnkkOqKsQxR+BbKRbrXQW7uTUjQ
MncISSRjTOjEW0mQScUCGxHYMeomkKYPm3eKxC38pxbtCF2T9qb9NgeXZE89hJiTO5gL7WYqTdLx
FMMxVGkiRmQlXWZcK8PxisEDVkw9essrHO5luP+3zipbpIcZ4BhKN8q8PK4St0QqfPV/leTh9Pow
pwJPOaCylo4H2TdWbdvL2kk5NUvTgEBIR0FJSit1PdZ+v+BcCTO/oWjzcw7zyjCaI0l24BeS7v6Y
i9Z+9GIFeWAYjNQmgr0tM7A/A8dQAcdY3fU97c6BkGnMbkou9ORwXFpHebjDkUuc+je9K9aehMKS
/7KgLdrtZhSEKpc2/HYMAd1+EXhUxNTuF4ahl80XBsHjvfUjHRe/F0plcMSMhMs8n1qen2ZSjg/L
UrOlA8Zj8Tu/tIJ6SaXFSufiMvi1kpz/odL034GEPXM+iaqOlyk4h9iOsb0/ypkCEDfmRqS4cR7D
u6nKmTdxJuci9Jt/CbP2jwgn+vLG/T0uj69GmTFjYqiBlHMlGkkm/nNEUVe2890IuAZ4FqODXtY6
16nYj+T24ji9cdTELmC3Q06Px0/BgUYcXYhDWQEpy0S0D4Zsn2fknjhgdTOgfZjMNMIbyFHJIov9
ItvAiuoWR2i21MM86BVQ0/IDJ9TrALOP+otgKCNBaj8MZ53k0OZlbK9gPKoGpC0denygvntaXxK3
z83UwXxQyrOBeEkZOxw/S1OAusaj68PQxox/CNxJKQga4R+IbnVCRptZomtgrGB6lYltONEeu2jw
ApkLs3V1MHPVcf6d531dOUHqwYbUGkJS7mgUqjpsy0Xt2OcM4mWMOwUXjzj6nfF6bcZSBo9Y2Vu6
biFyTIYM1USnKsqR+91Y2Kf3Vp56pUnhlgiOeKDu9JrbVRMPxBjzUc7n7m8rF4rOBL9d2ZphTdbH
PJ1fSj6TZxK9kJZsmIdnfGNrFJ5kCLI75abORaFHuU4/Bv3z1DN3NkK13MlzcX4P0Ify/Fkh8v85
zd+X0xDbH7ybYuKBEKOcYotpLELEBSk2z9aSl+qpylS1j4gSAdxEkJofs2uLgb0WZq3bKestEOpv
drt26iQalZ6c7X6NAekFnLgiIQYE1CKIyjuXtIW5u8e+xuZiHQJpwXgjUIA3EmvaakidZxp8yxhb
W7Yv18eVMG+NWHDB0HrmI3sIBAcZU8J6VtsVVH9NT/BI+q/Q9AkCt/AG6MUY1mLfb2Gv7+C3jLRS
bIGkuRcK59VpAwG90EhOhpLGihvrN3NFCKJYUsPMPmolp03UHbewwFnZGk4HWnEQbqxeIdGRg9dg
49DYbJkQ3PFODx+jRNK38PXkzz4EpLaLbflQkfE0eA5Q9gLwiHRt6mv2t/qIQTF8WZbdyC8cnk1M
PDMAbaoDMi/6XDS1BJXZbwA+9m7NenEQpwHG/t4RYwBnVGicNAUNGksu9LWEh0fMLPpfLRXrHPH4
19auAk0ed4b7CapJGGbBDUnAg+bH74QRPnQV2eaHPXS5X2cOEC25+HYLUVRGAwBBgEnfnhTPh3cw
S7IfWYTEk2dy3NufqeP/BAEVjq18xWKaGc/Z1yzG7CXB3EG6ujzpTc3xYbFDaqImepL5sJEAh+rF
5wkl10orAsUMmDowOhJeXiFztRQCZ9CZJnrd6Dgwp29UUw0bR6KBc/nostLmlUFwtaYc6lAwwfbw
Y1vw/261f5TWv3wIMoF1HQu2nXxYkxphInq+aH9QF0yZowSX9dDZPfQ8CeCxPG8IYYV0CZZqR89Z
8/fE4oxQd+585ivt4sUdCO6RRKppUd2576jchLJWb/lqcX4v4m0FBn3b+CRU/D2j3L0XoeA+6AXS
BxB8/F53XbZyqLvTv7CRMV+FoTxDcqOiLywHHm+Z/mvY+qoyFJLheTFDOe+lOGQfdrehMcZ49Xky
xQmSG1klDCPez6hBg/g1O5vF0B3v1HdS06DlC7/o8hGO2r+3h2uP9PRCf008DOesItAia33L/2Hp
2x7AUa0urzm6crs4/ja50M0Yd5NyH5cqOfLwsSJIohpHZI38WdjQ2NLeSm46PEnMqhJ29zVIkjgE
LDd482hCqr1B29/DlNVVaUNQKlTxkKMIqgL182JACvmlf6HjTPZqsBdKUB7u+YIXt4l/KNS4FXid
GP/6kfmLKZQCm6Izp6dURYpgx0HkznVMICDXqK30lUccHrVZ6CK4mvCM1Xr9uMP1ppgH19CbuRz8
VBUfvTcWRqq/UGXI/LunmY6KT4DbAvAcnhQH8A7yoIdIPR+zh2/5KAK5NQNoWqTFBeaL2krFTbd2
AChm/triZWCxGjdOvmGJ/NiSkj0c5eCWFZlDARznr55j7mqysE2d4XTCRkaItC7/nAzPgidQ0vcN
hvTNXyl8iz0ehdw0T7oe11HMHmC5bu2uSZLHc3G/6Axk8H1QX9RQK8o8oA3fMplslhtXPBbujFDF
lT8vbaVxH7GcxWa/Q1H7TKSpGCs1+J6omN/n0yWWZ+ahcEJZBLtgw5LjTtTwNUIkfjYWKxn6BfKh
TrVHAkPL0HGHbVnyihsLiLPH2pJ/KU3KpYetYEg9i5zpKwqWa4RMswAOOV/tcYCC+OtVVRdVIbp5
8F6qKyZNsZvg2f544Y43MbHQOxTCLw2Ywe9CLNnVX+8hV7UunQfj+ylkUULzbPS2p3fMjl0lus4L
6V/lANdOs163r7gCWELAoN8rFmi5EqTyzUbKzPas1SWN7euE7BJZdGlQJQOOSu70VxF9ZexQajxt
q0nOzHIY0dK69JbnOsYpwIx/UF3dnWQ1WRRFWvbpGG3JWra3g2wz6/1V3LpHjaOw4GzLtrFr7s0r
z5S553jx8shQeYsbTs7SJ1Uz6WQLxl0lhO6pxSdb2TUZAvXzK0sZinTon0CrD/h8PR4LdhoKN49G
rXSU/4YA+mEeBMBIxZMXYW2uP/s4qKNOkekvfQ0sVYc0MCCq5N+9ADScLXDVx4zAQ0dG41mBstMF
1GYq6TITNFkdqouo7GjDf2Pdqw9UU1IE4/heIVfuilTOQhkP5Dkmpcupj+XO5svnhLhgANcVQuwG
HE9C6ocB4qIpXQT0hmAsqFK4/nLepE5uDsrX3oM+E3K7SDhydKrx8rM9v5afzSAp2Hx/yzQQ8oQt
RJWVGRI9rNqzDOaR7W33EeqySae74m/SvBB6ejdTSNxIpo4FFy7nrzKDGoMytM59fzcWhXUKjFSL
NirInHQVj+wranBYv4/XH/SL6h87rSZGyCDd8WeFTOtd9PHJZYcRhHsXrLg7nDY6760g7Ny5yEYj
XESzMWdKajPDDvvGx/dekNCXFFqkgTgnEsnRTRpqJiLJc4XjJimv6wH/pMKDdQNuVG7VaZnKGriC
EW9kgMvnefUhaZ7fc5ttRq/KjsvaZTmywpf+VrbQ9M6Kx+uklB/qQ2G3jleBA7iroOkwZsEd+cAQ
sk3IN40xr94l/0JCgGq/AL69Hg3+Wp7eFtonqGzPxzeKZdAxAosiAFWjrfwIxY9pOHlBaOHP2SsN
DOYJygsmDwvQKq3UnSD3W70ILd4+xkEMzEe+ahplu+Y+w2wNBWLBGtAgT9nru1P24b5mzoDdVVLU
YEu2K3EjiczPLUPFO4SpnmfGd5U40+G+JmTiznoNFm/scFWfXmByaE/A18CaAvuKlCD0Ta3Gvvna
uziNh0LfeXgPGDHER0aonfBX5Mpsl4QoEO9raL26LqXeLVpN/IFd0XNvPUJrhFFw7sl2py2QnJ/O
HKOv/w5FW3ciYwU9gC2F9VDTEdoIBWX9whOAg4j/TkYqEOpjqELTAVXIhLJOaPibF2o5cCX0nkwM
m12ZZqUCmIybfUlMhEhOlBzt2VFWdP2qwRDc0OffgbDaZnH1gcnUmIo/jN5oPOWgIaSLAbrgvAY/
80YqQW1TM4YLZMO5wKp8cQCTrWEGLFJf0Owo/FLWTyVPnUCEvdU/3sYImJaX4YYwt4La0S8qtrSB
3rU6Ast0JRFi7JysedMxVRD/LyiipzVpIZB5O2OgjLP54lIPm1sLWHgED+VwCFS1rW7M0X1S5qUD
VgOCnltv7nPw8zAV8J/MxYf7oUbxxz/yHkOAo8JH0zN5wmLZdVHKWJXfARPEpr5Bdd2k8B86WEIO
OT+S0ScOGjTivi1pGsHltEMeUKXJf2oMRJOkbygooGAI/EC40eDVeDc78J29fGJ0nleTYMN6IuEF
wvMbRRqQ9TR2Y99ADy/Wy+C/FLDec8g1UTcEsRXfltpxFOmpbAk3Zv7R9OVYxvOTeS1JOy3hPz2U
YDNvrGE1PjarnqGAleq/GOMKgSgtf+qgd5Nh0MWPbTXxnGAPfJZ0Me12usGOZoZQFqgKDOMFxD+d
ZUAWhwnjOGShcygUrOwHGs24FbBFOq/fNEcpkFyKjAb1PawOxBZ98J5KcupMZOC5O8QhwvwLibhq
X80eq/6BfdfX+KBE7XD/jjtd3lD2RJYoQpvEU5BRUOOaXszu/FwbE9FjQDzIrXBtYxlu2ndaDwRE
nNMO7cC4gGCwmDzWWzxbr5NVuKmTVG8iHbsvXU7REtsu+VSgk8pbWOvIFnuteRKyC3iv9BdeXigC
cmTooT69aEFcaWSGWpg5WufrCxw7r+O2a23pi790hnjD/BJaK4i7qlWWi0VWmPOIpI34zSFoEVod
4LRlNomOsIkyrVFYwmZ4vqzwpTnG1hVha9RK7fjs1B+8lIeSjeeUcsFmuumQ3FJJu3ulixMg/7s1
ZhxnN14ZDjLvkyVxup+y1cx99AaGRzEaMxf/xOvAOph09iDQ+Qf7PpPc0KZzvnAgvYmJmm922/+L
k4vILnqP0KJPz/JV6u+tc1/WP2ymUIUNmh5ah96ezC/9n1VNpDyVIY5/jIcersQrKiqtAESSjxyC
p2wdimrMWP85bW99DZdIhiIMV9/1Zc/qURU9IND4GcACJuQ4gcvi/7cofYCGkIZYglX0PnzTx9iC
KNnLUd9pRddNFtSyuFlGLMjBEINATfRh8RLKEpOCRNvn+OruJ8Ug7X863FcQ1Da3v8Z+ixoxkd11
+TTvgjPSN53qW82UJY5bKhJ8Zlw/dHMd9kIBwZQKhFX6PphiDfvanEbqXTPbLDkhdlXtvk8+VjPx
ftjzD3pu9l4D9hrqIsUyMHdx3qPzQsB7NRqOY7C8DJCFN2Z/YZK/Wtp5lAaeJitt6hHHCcLmCGJI
N3RGykJqTKE83GeIkM8YHPJUD1uOaTDl+vEgAv+Mq02SS2Od52ebpQ/WbjB9RKSBoHip91C5noyo
Ci53EGyCGWp1Udl6jmOuAIRHGRnY2+sgbGs7QMtoDGOHOACzhYFF4vpMMK/kQORXKtL3FfdZjhr1
721Opwxa2l8jxygME2jSEW23ZJDMc8ONmJpfOqHGHsnj2ByePgUC33gCkdAYGEOLuf2DOdGZ9SGi
pIGBdZjcuoX3lI80KG8NUYPfDzUH4zfwdDyo46tGNRNQ5685mHxNANxlktCS1duhHp4IYKhsefwA
p8z/a0fkMdyGLF/k87HxV0oHQIbAuR0gIUo8kvIL2bp06pEsEqmXX8jzrpVIgy2LBdc2rtioxAOg
SifzAL4pKrSNbtuFNhCn5GtziE0Ro7Wu9mzgeKIZTJSf38xBM6VegiJYXgdkbby7MNLZ9KArxZr5
kpIVNzgZ1BduxWa5MN+GVE3VhirMa4hQgcUTJKq02nJt69rkOAS6b0g64X7mbkTzZSpbUuk1yM+2
XjsgH/O3VPInTbYpjw6xfOIYaEbIChm35wS5iKqoQr5oqkfuHv50jowNiEeTEZgH/kRwcftZ6VRv
ZCkhwhOLoQK4C/OGtgtiz+rvP64LmR7byjfl/LESKrkJwexEpScA7RXQEsGIvjL4OyzaLRnv/YzU
mtL20/vdz8v53Wzy7ONlteWCOOh0i6Lis/OfuYBHNDbxeRXhqLFBA0rOyI6swuNsNRgm12wdN9CH
QVhzxhsF7drOx6mBd27WCnWXAGc9066N9qdrWDs/KsZo0gzv80jGOOAVSJLkrjzE7FR+ncZvrbIS
dTead5FVD0g68PJiFGRBLuqVakluZSAeOBzxOr6x1h3ArP2Cjr+aBsneVK7foDINPq7AsvVSLDMs
m/jkc8L7dhk0q4rzX1UfIxavC6Vr/npzSGtU2oFGyIrEMfONjYMH7CHGUBcTEhUwVg1hIkWd780m
mVu3joEa+OHSSP0H7cyPW6s0AjRR6DD+eznnWH7yOTYi+1wrvNqhvyRXBu8xoF1Yeg0AW4A8gEWQ
qphjD8uMLjHNTgaIpb8ly2Jvx/1piX8kZ0jFqZDVUJTfdJIFSaUaV9ZAOWGoeBZYjC5yb95An1Wj
FyDpXn6FmFU6hsfSHn71ehLHUhQWiwuQZHjRZfmYkvJOgDdGA3O0W0sZaSZ9slfmeEwXA/wpJr7m
BUdX3tsUrEkewN2QqDH1J1a4d2budggcgNHSnGevB5suqxNxgCR3Io57ERM8fBpdhoAmTj/fuxgs
JNJlwm+lyi7kX4vIxzdqd18qnJ311uAOO8det+HqtnnrZDntIu4XS1TF1CFKc9tq8K7nUQXzGez2
mOPQv1Dz/GNp7cP6KMo0A42oYpOFj/wOEVM6J3UyYygi1SHQL0kq1VyVFGkK1wlXpRMZVTqpRBEx
hgk2s1Jp07ERWfpQY8L5c3Z06bZvRjVCVclsb8zMnrfWAMlQqWRpBCOKIFRxfyXH8IJlfHz5Hnng
I8ccCUiZTbZ3S2fzXlov2Tz7maAHyoHVeReJlanFCYu6tQbM1jxt9m1mEpS/Ix9pX2c7oOOFZ4d/
QhYt9UKy0iescRHbC+3RE427eOyGzgweNrkeiKQwxYvDTrheZ0Q6vu3ILUNBuGi49/SV3e/ObBtZ
I9au1TrkVPz+fMtchZUiY2QfL1mNnZA90T0lPO4uRUAXkWkytsztWE8qyfXMeS0W6fQkLbGohKIO
2cyL50RngBxaNlGUzXfh9UsO/p8gvXy2Kn3vj2OfuvlQTbxinPgm1ipb4jnMX3sPemfQt7rzHBZx
xD3dKnMv4YkRCRtwMttwKCmv9qEun/oQ2ore7TyOEw6pwO/KGDLeP6jOqUsfywBZP+6wyJXEKCSK
7yVaBUc9PSWo262fvIVZT0cFMSPNfR3qZPwHJTQhyxj6Fvlf1YfsOcxmZBGenjfZml/w65+cDG4G
FWR2f4AK4hyrVWLyAotYNMwGiBw7SenQPifEeqQ7Ou4t9RTFPDVIlQjmB7WhIYWz+ThYNfke4Nib
AB3DcOoi04COOAxYpNpajwSw6F9uRNGHSrj+JUANOxeNxmY34+03SdTiLtRADyby+vkY3Vtv5JB5
BCXiv3SKRM5T5A/y/4T5Iwp9BvrHpxFxRArhIh6Ocjme5ihN00nxtoN3pfv6zobjId3s/nP9J9Lf
/Dx8j8jBEG8/IdSNAlDvHS12PzgcwGG4Oebtt++YpPit3tGCISRfrf09kpkBjzFQzyk9oxNSsVsc
lLU4lruXJ8O+UrhO41I6y+PbW1pqXJpN70bytgk8wmLd/kao3ZRL7T+Yeh5nS+ZJ5Mz3PmLWxpMj
jbhTWoePhNC2ipCIPF94oLEy7FfdMy4mghWLE8p5c2FcLEpQcRj8zoaNVt4l7UvJeB4FHtwzZ011
zDCqj62cjisI14jtXZriQGggWldCABtsK/xf4jQnXGcG5HP9cmdr5HY1Sz8gaX0uN0/ZuSL0DENI
XEedwXtTg15vYLDwpEpeTkevXC0IJ1nyueF2nHUvg6gyAOBRuw8rDCpKtOqgUctbtl68MUJMIsnT
GpYQzUbWCYafQVzts6WdIbFE/CRtQMyS6sYQteM/dMr7vH8E64XiLR5UbEWmYDORh7NWqdqobyTd
DQmSJ/eW3cnKtGzZdhbLpQa81HsjBIaFWdU7BLVAK9dkL7pxRX8N4B2d7apWCgztS+jIoiv1hwFn
9jx9hfl/nix9/MvwGir+SALJ7T/Y0yFPx11Qwf5qdEGH/GFDjRDjYj+NrwP/nrFV8lmN0b4zOQBB
jYXG357TsOP6+wHl+zvRfpt+Rw9Gz5OBOEVAQOZz03ppodpO5hjyib34rPynHeEwz8GRtBOklJT7
oRwH35EesOVyJhYI8hH2TcqAEhJIKyTVmIOA7kZ/S+wG7H+zN3cwxb47dnK4ESZw1aKmp4M3l3gd
4Q90PB97QGjncB3thOz44TtzcZfDGa+BBTIAGz3MT4FGUyjuVlDLTXrNRmToWO7rSQ3rzF9fBCbY
6TI/WZsFqkjUPJz0xQ5Q5e1AB8wO35DvEHfGvDooDDFTFlpQYDwpYqERb68Zdz1dJ6ict/PtI7A0
OChF0xcy35GlxHEX8VVdG2EcjMFcIxpAWaBE71rE6YdOB8GoXISXFn2QOOJT6K4vAAQt+oe2yPn5
cpajQGWbJ/F8KVV3jDmvF3bGzARuXT/RnoCDLiaG0keOJN+MMd7idQ06i37KuBzYH8I36n+9g3H5
tdbXymoXXHv8Mb62wbHOg07oloQ2oFYmVywPZVccQ7v9i82RmInqBohMuhFKeYaaMnL3GVnn7Utq
ZiMkDupBYL11QjdmVfN2UHI9xlZi6l7XiNKEPV8wwy/CjSlnXOdMwVJLbaZUd98sZ4t7eS1ypU5Z
G7FnErGePJV3Dgx7RKM8MAcYoUys8Mwl/1/9lMYieeh/q3MVsLupRWFhusDHMrRdgpQbeEHODTSd
grLt301hPzsVlB6kDARuCB9gkqyIFdlRm4lkPJ5EN0P3fxQtKdtZiuLh/SlEnixrGCNnzZgY3fbk
JLsZ1qblRIfAwbFhDyDOkUilUl+70zBoQNAzyuKOZZIIBV5HY3Tik2UcgiQmO7TKTY/Wwpk6X/jO
lpjJy98uoDLwJ2ZHJG0a9MMN8uvXCh3FvUra4tRDxQLFI9tfR/0H/DUygGHotr3hyLUtypJmQDZe
Vk9hE10vlOCYCJf1RrVg8Ne0g68dmkUz6UjiIYJGRf7Dd0dKZ4IdOYaCAvOQ28FcP8l0kIj+2nGj
Kn1TT6PH4HLKHGUqgxiG1dqTpeKVzisWU30d4rqUssBxEY6Rj/YlENaWXcSzVD2n5knYybzSpKgs
GAahMUfoBGG9U3eAUUfNLGQA5K0pImCW6Hgd8bn+0SG71TCDzgEqqBA6ChmqoTqED4sZ8zLdCJWI
IWY1zGk6/mU2zaJ47mN7R2vtrSSv6sFgI6Llg3fqyfn04iTS6soifV3Ln5S3EODQzORo4y1L0R+I
aVS36QcXL8hEiE+B80uEGL9H+aMBAsKLFSG0H38AWbnSRUtf8hbIfJR/UxUbvImdNULJI9sly2JG
/u2n1eJ8XZT1nr0Bzot1NtXxP/d5XAN9DDZODSpNH7sxesQZy3c4fJukS/LDmfDzz49MsJClP1k2
2qJOYz5F4ENmq72Qq8JY77O0VvpOQM9ZiQXWCrzxWH+ZTHVZkMlwyaLtPPGyWXKXOlKF3cap0km/
yBLH8610UirOw566OU0RXbj8Avw/Cvvcf0l89wmaN6a2byqZfux6o5ju88+LhLtW4DzaHsLOp+iA
f5W1IIqQOg0GpaaFL/h5txPYKrKgzkgP7Pxt/8Ifwl77ZyTXTRrtrN3v/lAUYoeD0ralkx6DgAEg
iOc7B3SVg9YajFZSLC7XeXiTtsvQe/YkKG4KvzOBW0uaPaBIGJthMjXH5VtZ0cHnIPP0Kyvv1Tu8
1NzjuYdLHuectj5Ek/M6ZCmO4tsBgV9kr+2ghRjF556msrdmzsr1BhtIrfav0CS0WU9EYkkM4+Pk
nlvueR/542BiUFZXiyOHs7A0UrG+f02vQfwbcOLse7uznz0JKpg+E6Q4E/C0J3Ckxy6yTPK41s9G
0BpuYv6V+rr2MyF31Wu7Ki2N/KqvcOju10IMmu2GIfwPOPm5m6O7/JzQFLJUXX60MPpn5jSm6uRD
u1vyNkD2Jj/3c+qYRMr5XAg5R1LSrPLvtLdCzQH1gZwXtbKObpjcmKzuNoTqvWX5y6Lzfnbras9j
muVPbnIIXaekSAPxgKzYh14GCf/HgAwvqWl+rZLTY9SRRn7EGue5g5AZiulk4UKxD2+jT6PCHA/E
Ubk+N2MuDbJVp3y6MfihxsHkl7sRwNLR9TuFhoE2+4/EbYVLw1Ui7QmRFiXjVYap1RNthxDjRGrs
fwZxmSclmJJ95NoQmoehcSCm581D+m+T/3zeJREvNo7H4ZsGsURuqLGvUPUMYc0bVqFxE5bkASb+
hNEUYM4MJ79s4LyyzmiB9XSDWc1mkadJqOMh/enqUpkhshr2vQDe9C8fYXKbUym3Lq6OmamqDDkM
GQAdd1hyhfSiI5hP7EQiGdZB3ce3cn/Xulbyzyega5LhWk0gCjtELp9yN1dkxT4PDHcR/qZdKh3H
1xq5HRmBuHVA6+5A/AqOQtD20qRtwqC77aUh8hg3qM3HahXomjtxdfxWbPpbBwKZ7kZHnnGyX43E
6Z/odPBIpVB0ZqiwyY8L+wkQpOaJiGziu6t5eWarLFZVPVIPd4G+VIkL7mQnHCiwo+kJRZbovgMJ
8Vpu5xO4kaq7fK5v4vr+6UtjtkvulFeZHZCo0EdrWhkoaFbNySDOIoD3Dt6QucD0yFxNZNV798bk
nAIJyyJNiOTIQHrALfiRX6lzjZ1neV1/QCn7N8gJtapDqAul+RIxqRDNCoRGJEriZDt92RcreXir
Xo1Peb0b1UZNEjneHzJiXRRzs5H8oyj8dEbp7zjT+Arq6NudcoGzSt9kLlKoX1qrIMe9HvdlNN6O
oJ1U6vYHa1aT+QrWjCIMDDY+vJ2A8GFcbIdHyFFZZl45iCErhqdP6PqRtME2zXp1Gy3S4JU9aXcv
EdLu8/TcZcdWZ6hyTFILXlCwytJ2KIx1fifqnNFlPFTuuT6TeFXmjGmLqP0eq5iIJ1cOCRMwAHkS
VlSsRkGwSiQL1HR+1E/Z+udVhLoXMVA2TEa4YghOSRGjf+YCFr1RvgCPIUFZvntoM21ZDZiPZIww
fUuDPjZVrHwzM/T6FU2vqGr1wL85Ay6OgBk9hU2WckAidapu4gVbyeG2VwAEJmxvFoEINz+fwZRp
rR0f/+EvQNvBJ6ry2rzYcsZa/X5G/ivs/KZYuMw03tQ3ko3WFop8lQEcEASQl4LKzHujs1QG8D2m
ILd37ZkQY8GB6Jl8vDlqh+4uMO5EPWpQhWYTSSlrC8smJRQiNN+Kr7wBrjkCoiI/92XZHPa9agvV
i8ZcgoY4vEsrLlP8qbjSnuqZRl+KwOeo8rVbg0ocf3N8hyHCbCsPUFBoWIvOpsZdFhzV9PFnc7Oq
3mnItWDM/ybuA2zoD5iPR99Sf8+7NaPTEXQWN1AQUC5dS0a6ympBLCgEPgH8BcsZtyekWZXSwVRJ
hagfoYy7TF7IijHhi/nnpLaQXsZl4TLirISop8f2Q2P/I4S9ZFwwG4OXVQidUC149NugtFlLLedG
h1koZkFNGaJoNN7u6adlNaQ/xiXSlXJjv9o1QIoYm1SBr18U9+Znu19/dQ40Eq0BXn1Ey4SYqoAt
t3cYALR2d74BBLmsC3vrIn0gAjvlR+ytuX1L162yh49FeLJDQ7wqyE9BEydPh+wbsSNFgZt/T9uM
77OQDc87dlqU4Tmj+uoWVoPx7ITs4U0JCZsyg2tHRxGVc2zyS0aIZUn+fb/YgbHGqDEu/HWBuezi
EM/RfkWbn8XP+MBMgrgUv/TtTGKV/8FxCgc4bGf+HjGqzMEAjZxi4JT7XOJTAZRLUmmzHHK0CzYk
RRqu6GPT1jdibRQgzTFVMlSk2rwoMc6MZ+1FAarz6P4rAV0Sl135IshzK+oGpMJJsPQij1j2kp/F
6YVsO4rzgSuZUwLXhCaxLezdI8VoPZ7NwipCIe4gBnyzx5FHzIrncFju9qZjaPEwpcCwvnAY0NIi
xrlOTNNrBZK9CsvjhQ+TXtzRePh5Xv34VP4Xwmq5cH8PRwVUjsRDJmzrY9334jhXR0N2O4KSzNd4
cuSp1svLS1j7s3Z0KkF/sCUzvt5CK27xu7Vc1hRtgxXyt647dsXANqHUnyrPhED6pIoOAo46ltA5
O95+8aun9N40brJ/SrshXbx6mqV+v1hBWQEazIyLCEPsrYIsys02C0nRz5CxFzAhZS/4ZZdqyyt+
RfWzIAkHsiPmSxZTwom5Fvgnl0nYKkEcDe7DZsJXEjwwAphSJpm64If2wq15aYKWKr9QGpjWuT+U
9P1fsa2dZoInLKJevC1zjZFbL7Evo+EWT3rIBZ/yq20OVSbg5q3JcMHCqBdsSRcyBg5qIhN3csXQ
HcQqh6v/hr90TprgRg0p4PQwp3g2mQPiTh2nd1RD+161GGYy48UROyd2YbLjuzeb//H8CCl1+bA2
s+IrYDuLF227XZ8llrUWmBqlGFfW/JlFXo9Y7A0EKTr754YWCZMx1AqnbB6I0YuS+AuG0KI1taDE
9l5ssPcckeSunjw/Elvd1d7PhFeNUCF2vr7uXTIo8UmXrLZjMI5glO1eyfOqSYPFEx3otSGEfWgZ
QPXRx08eSseEVsL91SlDPx/uxaYjLtROOOJRVDw1lBrey8i5EP1UP148M7U1fKhzoKS4kLowPTr9
Qlql3eEyTBpZ6NgJdSmF/oHfeEXsEXa5Wo4k5yk/4NK0Qzw2wwJsOK+vxjPfWUDmTJtuOm1UjcuU
mYikLf4vuI+FMR2mmmZtAZ4WO2LjZNxbemDZ8Tp/fYMP+t+FiQjKBupkpM1AgRIM4HxsZvvfTBon
TzA+yDMNpEgPm40Cymu4dWt6f1H321nTbzXWnz5ArhmXe9GI7rEqCKyvY11cooxZ1mrcmdIiwqif
UroPJvphx2kwyZrqjn/CkNuCoe9EFN+UwH6yZOsOYj3IXzQ18OMGkMtXwgS12wAg1lCg3I688YxM
/Z3PgKEG/neg1NysdBegn7lNpqZj3MapEbqksWykvBPvqWlEhrz0EzaTNZuZuYpCNHpW6Wb/rOoE
rR8afsRk/8qtF5+nS29ji8Y5LW3cRN0rgiIvDbyk5wr8Pnq+zqr8ffBYMK+Kd4NTfOVgZHdy/Tt6
CGsP68vsT5J0sdgalZUkMMABvEZSk0TFKIDFO6SFrM8YS2RV//eZ7HZ6TSKlU9vjg+5wQVMbogNB
qHzyUxT/eMp2/Nftwv4QzH3eKvzCbm/ZN57x7J6cDtlsuMLkRyMJ4kjtaplE8IzHAW1Ds6gqGSkX
aianFg4utNWFtuEy+OxFaVcoYUqnB3He4pnvBayuacVSLoA3/mAvidj8TQpoZJ2kawnvHTxiHoGv
7Wp86qs8ANbLLEXs8glJwREAomXn6Go3aE3uzsa7udgkhQvG1wbVwPPRv9vi1QXXK4azWxj8KlKj
5GoFbyQWxStqydqpWbcAZ9ik+s+ULu40mSFXeEbreEf+X8Dp6guPZkHSiVRrOT8weyCPWeO2W2tX
XNZ0QbZx1UVlqEOBI8bBWLuwM60+p/gAzrEmuWmBCGAhqqIPLm6CQY90nHlMnTi3jhUA2RK/D8dq
FXj9QbaURucfac1wvq7+zyXZKkvWszHd5JoWmwkVJ5LiYUIAwkSWgJP8BfsXfx1sjFLM2imYfu2p
4VrmyD/fOTel7ItR2zrsjAaWhE93RRYZbQAq11gzH+rowpPGCYzdpeoHSxq7LJT2R15V0YKZfiog
8F+00QElNwUVdBaCVxAcicm1CsTvMkjwBjumh6fxVUEz3u0KRMXyrnPOHpUcuD2ZOTe4FTUiujlz
s1AvDXQKmPaOens1X4igo+oT1IYG3FjBkEtKLp6+7b9EiI5yiPr01kKgP6p2ELd+yKJlm0cUvhJx
wchipebxk+LxEG6YTQpJDo50f7kvSXa5SQX9IbfpzG6i5YXAfzw5oyh7rSGXbtIEgpbc2wnIcOEI
bNFeM0hKWjxbcyPVT2rG7v4+CLeE8RgIuVCTm0LNo5LCTwH9AgCojeRs4kxjuGn6IbhcHYSLvTxJ
m5xxxfK4qwbxbM8kcNSw8SvsVP/RMjwnOMR+jZsCPJTWLGqnyHjH4USOmZOo3lL4nFVFxtuAnm8T
7Hlej/2lf6bVTP5mBWfgNvEYohJb8Y7S6c4WmmTuPOopX2RUn1i+jBbg1yJysnlFeHQNOdp2CAEt
TtATbeVDB/LHS4zhB8pVWnbxUALoCv0vx1SzSI9PiecFwscM7xj3AssJy+i3kubwaSK5Q1wgr5MY
d+y3W6Ut0x1znughVadWeKn3ltsSpaDMPdG0VKmPe0qABib48WAXEks8iCh9dM8LSDN4Vy3/dblS
BMWggCWKHACykvSpySNjvyVAYArbYisfICbs0Z2WvwP8A8lI3Hj+YMuhxPX45ySpg+DyDJs5jHyg
4rmLiiohxMCt7piA0HIbtxY1NLGj8bO0QNherIgSCjc+4EjXNudh022MluPGiAA5gXFxtZn/Ge6q
wIEqTKIUK/NsG6FX3BLySkr4EFxzMEJ8dxeERIgNBaAQ1PZHxGWe7iqQlQpOLeGGdT/SJc7io/zn
Oo5T5at7eB8KXTnFcPN9C4Ykio7U5mTcCf+8QxZhm52wLCk2mcN9NpRqExc8WwaI+C2ZNm2Zb06F
mR6PKCRz16L2y+mVnx/ufhzO3d1p6ekpHTyiNUnvS1N/R2lIjymbAN9j/G/78Uht7f3yUiWmcpeM
hBlaVaLTRb1vMj/RRyusp4F7dP0hesH/BMuDO5xATX6exxWPatPcS+d8eOq68+0F+WTf0Bxmy6o+
N/CtB9IMSCfNoDkfzv7Gop/8G67Lyh0BBSZ1TfqOkvDUPyIiXgCT4WhjXtag5FMGxu6FLAQVQuXc
fxLB7llOoSl0pKFlH1QQiKupRTRdGV+vD1hQtujizUkl0jiV1Ljucp0UDD7ENchWaloBYJI4qmLS
6gAR0mW0T7V+kubXkWXJ26dlf19YuTa2S5QxiJEGNWgeweTSFuy48AwCoukUQ+7vZPi1RKa5zCAQ
0hkNs36fZOGGyJocjKTlV0ak5CGEdiDXv2/WsuKcQ8oE8AOC5USyOsCYwYg4+aCSjFXEPmE5XnTl
rEWYlad4YFqu17+Tu9nHYFJpEkA3by0hvGka0wzJTaX0LWfMSA+3duWqsXR4V0UyByMSldOzRuQs
u42gI/QTzvH8g3UlPw3mCD2o8hbqZn0ZDQffQUtxOAYg3OHQ2DG5GlSbAXq7qeQKMMOARNHWB5QZ
z4bI11OA52bozjhs2R+oxcc9TCfzP2B0Cs3dhO5/nngUXJDzsDEjBCDa6bcyGKdiQH6s1eiQcjSQ
m+977MSxvt3obu6H2DYgUOyQgnT/InNocCtA1VbaOYV/eZsP3fph6NEGHIBwLmDrkSTIetKD+gF7
sWRL2YMRIjFl2KtVYcwjBvrqhYzf6Q14TitHdHMK7reyGr+l8s94otKZ5vfcJ7pesJUk44kJ4g2J
r/Q+LeJ6X8iVqkWxnoEPCDbs+cIRr4PYdGKtHLR5ZggAU8cKuu+Wee3Gv3vhBvrmrlVqLMNdtvTj
QDqEqRuGJr5LD2Ed3mZ9U10tQQj4bpgPOPTF8vA4XX4xfVGgf6ou26bnJcKDZii9mZdnWWs7EXOH
Nsus2h4r5t0b5lS9e2F6WnvG+fJp0JeZIMhAyt49f1alMdMBtLx1ERWkE4+AyX/E+GCTMyrE/zDc
UEkpLGeEPXlk+jKaZ3YH1rGsMG/ZpqyIpvAqOYxTt7IymjoWVBtWeNBX8wc9l6in0QU0i+JaY/AW
UDyj939xwLNQ6mUh8HdJyYXxURHeI0jfm0MXbB/DK1A+GDE1XsuhUaQvPkXn90TpQRsZsAlkg9mD
xbkYKFFu3PTfx9PnwnJTK1rvNhfCaAUvuPuvA8Haw+OGBYr2zf0DfAhh8ENrPLRYk1EhBNIkh8J2
nKtvHf72dF7MfI6xPX1qe9i3wDwp57W4sDuFNtTsIZJR9aPDq42Cdi1Ux8SseYrtqto3drB0My/w
iEMC1NX4V3ifPlBrQuBo/iKs7V1U66x6/7FA5Z/o6pNhPgZI6b+DGvIIddpxk6w/pz7Kx4X0eHzm
5V4q8XiJgCPZWVk5a5H2Q3YD7AXI/6FCNGLfBA+rtkw4cvK4VqcFAlE5IiqCOJ3bZ+nCIz6n4DAt
5vCw+ZhaY/ei36CODo0dj4kseCSGuCAO77YTt2M6Osf/4rkzuS79P+YrmTuKj629iXwdGwZ4tSyT
9YPlw7izRrtnwjCP72t+XnCDk+GvCo82WbVGdINRQ1WLzrc4Ue6rjuKtoHQ2PLUMGMKT/wd66TUp
XoqRYAHbGTSv9PcVEbE3khL5jmRju9mqHRWcSErJwuxH8xHiCZHRMzzEwEViSoaBsFAhhB/VCvms
K5UoKfqibyc2Zu96uuhfIz8P44ObGKuAs1oiS0rnr2LNF2qDBNz9V0Lb30EoWrdjHF6CtVu0iNWS
YzZN3Vif10v0WPhfCc1H4mCGEOVMO+T66MX5Oqcir3Bnt8uZ51HdvvyHisUJSwKCcleW5M82QU49
BSVQerb3Ka9N4Uqx7sLMqDNZ29Lpl8KSg91v5o4cNTCJesuC2P3GVS57YwRNld2zmpOecvBindvL
ny2OUWf5BT0GgUqeZBf4RWihc8lgE4qFSDy5f/9Utt821dnDbhj1cd13gSbQtSUAJutAr5MiDtD+
pP24gZYe+3Zb7ruOJi8b+vqiSvDVAlq2IMfK0VUP8NIKskd5JGBXwCeEY5tjGTjivh4VaXwx2p0r
yGcqMfY00AjNo2vZewp+uCHPW0V9z/CFVpLzVOPzfyEYGp6gDQlqaEuc39KzLCAnUW9V4yNe/pUh
s0PmQdPjv4WnnsL0y/1c5S7BlJSVbr3RGkJDYziDF1E0jMDpisW2sHZYw9lS3fe0h2ZX9/YKVtIi
vTlNZG0OdcafcrS5v/wOIYnxPPJOhx2ZYP3xsGyZeEUeN1QNwUhb603EprzjndNarXmSZ3Un/+oZ
Lp0gv47RlsUvgJefs9FGkLTmQnRCuX/c1nhxCyuXbjOdnh00732S/Pu3m6BY69b7I62qWtxR9Y2A
7D3q37bFUOuDxZWdYZchK2Fxu29NsxAZR6O+4zTFhT2i3Vh5tj7JtkzXVUf9MbSUXG+AUWujI+ps
/hEld/UUP3pvH580WlHeJuxUW0XmCkdulHuIQnXkSCPOJxevypS29LCya6at37vduK9uW6YTlY+T
SiB8WFgqPHGmD6jH1x5pBULPLbe5/sbiHSXeI9mck8U7QiYFMOLzD5C0r0EQpAgH6xfgNhfxLJOB
4A4jfJC+TALOkP6jptB0XdkBonyBid/Fxdo6w6NICTITdReeELW/OQ8sZeVMsqYi+z6uvuyphs9S
ZT6kjMrGE239KN0kwb6W7r/xQ1cBq4DbA2DLqW7n2SIbopRuYawAT60tWpSe8gVJrZLl0wa1W7CG
we6AhNGHbvSpIXwx0kRJeMTe3UkVYKQSyW1V9hGki1xzk+7TK36m61RJY++SbI/3/rvNhYM3oAR8
3PX0xSzrPaWa+hLTwM791f562AVknYML9O9voo7sHMMC+u9zqXGV0QVZic8CtjxQrOloZNrOGbtp
ZJO14k0Aar4JjuEBbwnVSX+RBGTs3WsR9n+cTPZyej8S7Y8i/xFvD2krLI8q0xpnp0tdoL+4zhFn
jfs6N+Yvd0rKd6OmbAWQp0jriCiDPzKn6TxdK4NOFElECvWie3DBjaPO+qtD8M3spdQYOStT262o
DamfVVgkrZMeo0szp3WG450xTRk/vJSoKrg27y+mo2cY8fO6gJb2np/q0Lsj28PCfiyTcYOOwRFj
5c+4DFvvi3Z0jTHdxLr03OI6wUvK9eIsnwm1S+LzlDWPN9vbaLcZq/27fYC/hcbnzYEEt7RNcbSW
7UatCweMaF2+tllmC/nRNyjSmj4OLocOyenKhvn7FJxTMDuxsD46JA3FIsc6Ro5W3aTW53WiOkhI
uWhXIMV1ulcKpY/2UDcMgZow8javkUB5cc7603fcuD0KIaAfCjxCy053/VSdObU0rjAW+IfjJpER
1zcqx/SWqQVpmxy2kS7xFVWsCG9mjPLGXum13f39jVZIen+5Vk4ruRGn63n/qH1M/rx0n6nlcZHT
AWINmyP1tl9g85Ar0/hpfW+pzRKRgFFmzLe6PijBnlEADNoHkSnhNduTPAAc3C8YSeaom1xGTGSj
PDu2AjdBSkpQLLJlhOl1H8HW5vYOk8g7CZZIv0yrawIALNqhbf52lrKeP9oPy7XeKC/18vRK8Yii
nijB7Y4KGNfN19ge2vKPlQ+MHSLW9Yp0ssZHM5Zn+TCb++tn4dgq1FoRHHUJCFIuhNSYefOaWozD
VD2mhb84pbvcsNdissEBJ5VNsvLjXqwB+6vjLrdLB46GmqpVLeeDNJjBrCNikYRfMu4rB05NdmrV
4GBC3X5MmHcag9K2ItWAGAvE+X6i3lmqJLgaT+eo7hD85cXns1DX/KJVbOrTNa8W61iWcYwakMUE
0xux0msL158Xx0EbthQqaou3BLAl0UViShS5LluPLWCuydvRevXB1C4zm5NmZd3jpowSaz1N7VL1
gCjGw/zjAy39d8ej/4NnZJRD3UKqdgWqgnQDiSNRrJ5vIoieeh95WdNYgJxFPO3HZWrmGt6loKSu
022zALox46wxZxnCpGuATWELsbS21KU48tAKQY5efmELeQQn+PZWnd06Rc4bf+nC2OixNTYxqxWd
/iUGtMQQFrKh6pQdIL0jNxWuQRga1190eN2c6aYTtrKZkl//GGcd1ZPHY7JpvF3ygZ51RIFwY5ta
U4pZPgZxFqg4lsldecs4GlQLNCcpdL7Fy3uNypsLjR3mVnjQDruNMhM0hl8O6GWxGBc9GuR8XjP3
Zu8q1Gad4sNxdJOTbzlFh+eKOsN0B1BP0vOQJ3QvKwSeLWEFyXqt/vwfPT11+7fHqgj+TI8nut3w
OLSYNHQZ2zFA3SRGytcHDrwULFECa4UjOr7O6UclFpuDwisSdhhnvWg6vl7XImT/gSlx4huYEYfk
CfQAVNUbojfqlPZI4WraID8QAI8pTUcMlt6GRFYMisI/B1mhbk84t0C/mCDtG3JsjMZBt+sG+oAf
x8igUfHOFwo2kWfbppqgO8FOuhwdjXdUyiaSCCl4+SACwwr5O+ctd3ICgdPfi66QzB9QWGz9HBhz
kNIV0wgSVnMW0WMD4W0y2o55SIxxor7nlEMj86pQfizpgVmTdVww+86l8Xgrgo8orBp5ciPk0PmG
hLK1TGKMQfWMk/FtP8EmXx6HunzOHhtxWN2lwTYMJfsDRtqojpWMkvEjhNpafAC4h8qeez8pb3c9
Mp4QYRbVH0l9v6n4QiRls2ayfV0BOgxZWkQs9iOESsIhJPyGxokzbv3fu02Scc5kNL4khMShxFHs
EHtO6WbqaYrKXCOibS58c4NvVuXY2HxAapSQmDLt/uI1pzF23R031PX6iBrF+DKXskIW3fVYWTN3
X3lrjZZqky9kxYXjuOOQ4o4tUKvfNd2VFmg5yaJH5prGrYuliRjU2CxyWn6EY2EXIddzp5Pb6quv
ac+49U0klYULCYB1BMloA/GRpRwxLPn9kt+nH4iMUeEwbPdR+tQ4WoBofyUDflUhf3bkJdLFyOUi
Q3Le5LSR+OfliJFgUyy6NLhNHVU7Hm12JRAy05W7qkQq4OF2JJPy3gyybkKjOtGS3iE9pLZzQ7P9
/OWcPKSFc+E4P9YHkdrklwbzXFNC9j1k5arSr+4LA6U8O3qM18WLGxjt8oY3yGH5kvZc7KPRlMXK
e7lVsJxQctGYmRFMPeFGqB8URUndFSHiRK0m6eavrZKr/V9+rM9KX1JWE6G3tMm+yEoOp9o0xBZe
W3fCeUWstUobW7b+F8urOl8/3Dx023T4tx9USGhBW+vErpInZDtU9ih/xUSs7Rix3fGsoT0pdw3L
HzyQIJPyFvF02RKfU5EQxgDB/Nhrepe6w4qY6uSqmprsQre7xgQJt7LPlCrlBc4IqoPkBf3S02nc
gDX0FJynDxWzPK8Z4nQVg8zlTZJERyENFpE2ZS9wkxQn2KLZ8W98YedU0CVQNYKw2BbPzswoyf8P
cfdDahG6MX+enYL6pwTAD6ljHvoUvYrXIvFyrwVyoswM2dzkolPT4ciH1NarT5/9szKgW/p/jD7m
SHo4NW1eG989eYX0yfXB59fc1Jyrw7nLLyAIErsbftLdTcsBlxmIWGrQRlhu/WxQKT1nOB718wHK
nZwRxPeS74GmhIJvMZTfZVrjdtcz5VchC/WsluhnGVsFuEU+RIGQ76cntERlsP8n5t4N49UyM68+
Kd27nfWxwGbF1VbQ/9OknG60lLI/akOLwQCEA7cfZVz5IXYCb2OMkkfIvoGiWdbMwD0BNSNu9jqQ
GOt0vjLDNal3ArdoSHPaYdRjoZQOmDevvBApWK41ZnqaalcutPKuFXQ7+gFo4mVZmnbMjBjNJFB+
QY0gMhSMMLK3U7HU8vIMgGX5K8RgZe8hnuQFyP8/gb28c2wAhl6oKg9KJzjcF5DKeQhyj4dGQZba
eEMxNqlvzut3UTehFb2usFHiH7vqz9EbKjx1hP1JOnzAJS9w6pQuFvRp6M/nNVsILGkjsK+8Z48m
1B+nhQdXMxiggSbqyjE9/pjOuzRyun5/4lvA1F5Qg1dNtLUxR8b9p746rT+l3gQfz9+giOZXio4C
BqLjvK2RHdpALkUPvRkxVledpM4XnyfYHHrxeMyK2kuCf42GwlmQF+ynzmVT0IlQXYNBEpLu3hih
BDj+4mn2tA6QV4mpT6xPNSSNYVxdk0KMvy29ROGuEeZFYegnhbP+mFhcK2ca1+NQysJglJCyBmzg
kzdT8tmOWiDYlQEHCDOatufVqmJA+5VZkVBJQ5szIVz6YiVRhmcq7ImlfqTCGyKIWYZc3d15vAga
qM3IVxMwraCcj+z/kqtWuCq6aU6hZGRmWrfUsfY+1WzXQSF9ZZmx6rOTDLuMEUw17G6oKht90dA4
YyxfuPs7giejtj5QkuFLF9I6CLA28stv8bLUlruEyiR1Wwl3+8qLgSICxbWK7bTw/iAdtO/JFfSK
79ZL05W2xL0lpTRnyIUt3fpXcT8aGjRuH5itbrB3ZCxlhDZie5P1IloEiH8fNT8pyCm8sldAQlOt
02jTxynjAojypM5gCBGzHv9p5g6XCHQOFSiaVwNJUF9D/aQuHa3JaLAjzjVgVon7ts7C2kwQF9EZ
sCNfkUC3I9YFZ5EqmXHY5czON1DINxAqJ15UoW1/2CfWuWvjBAOwGpC64Da5sg4z/Srm27nvy7vo
gkz9HU0bXIhwzmELqZo0E8/W1tuzCKgsUz1uWKcnZXEXjYyCRDGAf0mPC/thwbRzPPojW63c0AeQ
Rc0ijiNgtrvX7TEqkvG+5b73Ak7ytpAzcANGEp2zcJLLFAdCui8t8I5nGxhRtW0n/9yQPt2hvhez
CvwkFL48tfy7ie8QDqmfH64C9yDB1NZ69EE34iEjrMFxBSqPmLEi02E4ciCMGjRV8dX1gLKo4Fht
fldGaihKqGJD5sbYMo4M4XK8FXSb3rFJR07TAE0QjEzsvzwndbfUwLP91KObS5yCDll5oRhaA2OE
VJmlHhbV0bA44wVZyLEb5aByzLSU3BISRxGn5H/ahzpU72NZJ6hLFh4QCetX6LbOMDqXqB0DPBoz
m+F9L1NcagT8bl0Nf4iGkOBO24fbe2STVrzfhzzC6f8f7NA0zONZnNEVUq7GWINIwM1ubwwQPOEl
cfgofJuZwSKWDVUzrHK2+QocQIrnCICsDBbks8Akk0TTBC6niDEplngRx+xJxmle3GpeJU8iPhNu
m/0ndmv0fddymRlCsNJ/CuVYC3pSS8dPQF17eBHBnDf+jW/rw4HjWRQbsjEC1sxrH9RA3JJXqNer
cubfMjvDtrv1x0biSccumKEbma4wvFQMfQgYZe8IC4oSM6Cyz8vUs8R6bDJl4c51iZDwd6GrzCu1
F1uOxwJqhz4H8tLDqm5FQV3s6PoJ/225fo8t19saPpoK9vl20yv+3yVF4Sw4u56WDjEMn/82RWOH
PJtWYMhAonCWm3SX1EpQch2uwUZH/NKHK/VN4UfbYLAGTbu9q6CGJkP0OHoPMOpgP8zO1APiSp6H
75fArMmH/FAAsOWnSdlOyIjoTyN+MjZIHLdC7fnZCZ0ZaEdS6fF7oXZsNMs6CTV7o1nUgqL+IQdr
5cbP7hKYuEC/Xo+Bofbr+HIu/vP+STac24t7tsCfXx0iBUL37J8sJNJdqhotTbE+qXPvaIfwvsvL
syHJhRyG0Zh1RHMDX2xEi6tv++XSl+sFDkj/O+KtXKXjfAikyM73UKPdIPzVWoH3Q7j63O3+f3Hr
NJ9yRQNW9C2Uf7AjXGu/Us3GJWT0qaaydgekCZb7HNa+hoi+gg2pcAqEfS4pNl+Ymo3ybbtVJQ6C
e2yTCpY+neAjQocLfgx6o7lKScwY/vBW4GKpEuOfP9o9pq0NhRfFuez1b4MEUSxcvVVfJnr81bko
zDSkWQKZRcR4koS2KZi5b9CFXl2a6tqSiqYZzTzBdlVESqbUwNZidwnClT3OYxfjyK6OSjhuCE6r
Jbg1hLzDHOmDnH27F3UwWfqKZWR7+GQBzXzyL2WxLE0QchXJhpk0IQBhlZH8HPCCCl87Mg2xMg0T
J96iNI1yrfR4LzBizG46kzi431jcJ9cKiNDzrLPEstYa0QxBUaqlSTzzpVqrv9qrJ+TDEbB0QwI+
C2tQSz7zZ9n6XRmDgwgVFUzrWYy5E0VJEUOkCzovpQlgoVRyCIVvF0F47LyHEftdwjXYwfqOCtbQ
mxK3lfATxElUUO/PYjJR8UCqu4hsKIDBuvs6oHZfKQM9YZD+hfWJi1hGcAEXRyxuBFD7S8Dr4C06
o0tYFzGfXnm+qEAstIXs+pUnbhptmDq0kIMQz/053jeT1sFngSs5VF+J9CJWsZRZi7a4YWvP3W6K
ma7mzZFsfL0BcwjTmMxsDq1IE7YoQ1ccTItqn/ejHgIcYcAq/tMMd5FXFKmV3C+3p5CAPjQbb7Ub
pGx8xUftDhNZNiKGyt5/HkIPDOq/3gYIhRRAXOeZaJ/6y91w3KsnAXyU/7Jg/+wmsKTLe9mumtNA
+q8XMuiRnGUi+x18SWo05S7WQBfhri0yHN7UqtVGnf0VyJPXLT2YXZYWh4jVe2OIUGPFtZfhZ4kL
vUhZMnbZnTKg2uDGJTf0vtMmZvbtLvXXkeDON9YcPDb2bCDy4ysE3KOYpw4ZhGmfFtHPFuYjDJa3
dwrcql8LKs1I4YIMlNd1SBrKHqCh54OONjMCJ13qZ+xhYjI3VCaIF9wu2e3nN2hUQsPkg+v+e7D+
xbxfOK4+KI55ClB4DF78L9cuVQKWGVr0M3RlC5qLliTXPar5nNN3oHq42usP6jyxiUYvVH3AkBQf
wyIOEduJI5VcQqeqKzIGomR7yFbpHyIgQfgTYE6ez3Uv62qvY7+iYbh78fuqe6Q1dOzIstPH3x1w
QQjgoxVmqbGIcoHqy9iBPgj3IwrYE+2+2Lo5tLmnQpaQxzIbY8XIroBNu9E5Ee+fUMFrZ2AeuyXP
BwAJ1447W+hixUbnDafMdNcO8fAJQvEK1uwRE1ZKZgiTEWWlBK6OXtXtEttQ/4/RPHEik7RFI8q3
sTRqiHvkhcs3nE/QpoTErhVOBysds3OGU+L1Zz9vw7QOqTG5gzdaquJBqoZBaofWtjfsQfEBi1FA
mBPpS3vKYAb0vtdsyEyLhbTTOVle98cTstH7clyBFNTNpFTLp939hgha8fKpjGYtoEnksDCAkjNJ
f4zLR0W1mNSYNNPrC6shKZz5rVpDRHodApoFwefbGyLd1hpsIuAepag3cnCMo6gGq7cyOkY/GO73
yZUO9SYcAqX1TWZ6HgndNbRIu5li/TMsw6Nb/MC70VqJ3AdaBHDhSM8qY/O4/WlTP7Tms5NZzJ+w
lKnOUiGCYhpvWEJPNVjDVMcsytA03PFrc1bhicJV6jHMYZpv4a0G+gGwGVdKfpbyYz7/wttkeVz0
qHYEQHQnmq5JXrVeago2pOqRVq3uZcDn/MEJU+OQLP5rgUVYki/AySBMtHBsQ06mRs0CJhlWghD+
Fnp6ufW7EZF1XXwW0Jf9REehv/LwuowLBjwY4Vb1Ft5vpuVukXeihgnfegWFPiEv5p56Kybu8yqA
bUQ7ADgWVq4WcQOFtNmXaQSa3eAxnNcJedEBZAWi2se8tYQBEJUmhnQuD4VJdIGbDhDZNM+aycSv
F4hrFncAE8aN6D6t3VbERlI/GZgpezUEvL7qXnGUt4QK2lhUpnb8dEbi5e/TdJqlkslZHdw5MEgz
NFpeTztUe1QEweIUyxWGnnQZbjrxCMZFP4SDwHPBBly7PNSah20QiZ/ZMeWrgVZOz4e9OPdOmfNU
GIVnQzwbBkT/Ng2EYMpiOJgJr3HkvfNqzJiF3Po56nL/y1yRMoibNsTubGzO4+9ObxSE7x1vfSBi
5BMHxCPM5xCJZvL/Lmq/itvWHmOaJiOtNWfjQ94YAEkaPqjTx1H+69buM0h1WKfY8SD2cO3B8+uU
hlsuq0xY76AOoCPl7+eFYK6O/ROmpRnFwrNO7B2/tEnFg7ApUg2MSo5MqfGr7CVn4kpLBi3/wlup
M4OkMHW9mykXDE30zl6ua/8bgre69BStuxLtEuOaQQAMbQX33V+SIMBAdmRM8dqWrbT3PfvJ1MMt
rN1XdgHwH30EkBZhxkhV6+n2l9t0E6LD9uiFqAkFYcXczMjUKvJqre4FTg4lQwViOfSXOPMvtYfR
UG8jkLzoImhB207aZyPWDPzWVepKAzfnMYxWwNb6/crBH1W05M4SCtrKg+BSBs6e+S8hM/zfH3Qo
SH229uE+a3+UlRoycuXgSpltNymSjl3TwopIOO/cX/bd8hGPwtpOK5/hh2K0C5X4w7ipNdcXVTFu
VMu9n7KNrmKL/My7gs/ynOA8gQN69R6H9aJaAAjOnWAF40kdTjwEZ7LNIhXeLmEEyJH1AGIAzl0d
a1kLDBl187JtmqO0QIR868uo4ROGN58j6dvNo8mhC8HkBDTAq++mMppd70LMQFNZO+aWV0v2k7c8
ft6zJMfs5aTETEUCm8a880x64eraPmJcaYpGdEP7Dmud7pBfohmouaVFQ3HOzppiB+qGklkT12iM
btyZrwQ/33uzcj8Lv1FK8Kt6RiAlC0vkccGe+eYmVtEMltFbaqndTU/pVHRUmFlBrn1bGOWkc9WJ
JaV+WgEmnfKN65p6Ck4MGQTRcldtkebC2l1c03LPEMNjOqPqX8l7wsKQQ/3iEyJ7EsqCS95KCKg+
PnTOPWAYEIjqNUIYrBoUyCFjQurgcubMhkI0ASI6020r52wg6zIsJC88q1Z3MYmzlMRVQ8ZLTYGL
zJnZePPj1XVgfcGlnBh2KvBj72M7IfVw90EwEnurZ2bzDHx0pi4xviE50f7O1kRV/K/gUOdF8Q19
rAHQmx8iLDj7hPhpV9F/89HMWNh3QWgN6jZctShSrQ5omlKc/XsfbqBpKuLxFzVySYL9dvweW4gP
LODN19Vs5KGvusDBRcftVorhBfOXHBqvWxYY9lIURpNeAlR8qPnZFwgtcxzY6sb3DWn+BH8Tc/nt
/JynXVnba/0RRlwvkX/tYafKyIAjQF/6V32ls5t55/1V91fgOyAZYeFWxo9dxG9g6qgW/N39RSKI
gf6nmLHofWUzncrSiL+FIwhVbjDwxE111H6X6FNBmR5cuhES4dZHpX2yTkADArNcCKCSeffV5rsE
5WjtlZ5vk7cNXbIVJIPaDfizKP79wdHgQSTvISAm/zGQf+pg+z/cxBjQDyfcmNihG124wv+uhEsd
aUYLyhITn2M6xNmjLYN7gdyAUdmgalow8zDjYeYUDuxcuIIhUKx8wpETlkw8SYG3ZahD7wp/dWRh
BG9H/rqBZcFhRMLFyE3d6syQT5jNeD+iZ1HBcZzkdx1xuq+jO9p+HZUtDF+mf4a30qvpX/mgcip/
kFFO6wBvd7pGSYcyEUg8S3K7o0tF2UOxT6YwE6iK+o0mjU41a+tOI3YSF+Nt3AMORF+YfwK2wd/o
sVqYEgkU9J/2WPwHjbhZr0n2ACjU7/Am3YWTIi9XXPeCofsIRlYGpTBtKukBaP2t1oUfdPAiO456
j98tQBlouDq/Q5BG/01v04FBehf25TjojBxs7xKZxSNG7MpNOtOhYi+E7GvdFhf8lOA8gK7nS6aC
2vvD+hKqTfE1NrFF+kxIvLnFh5lIpCrr/+uI+XUs2xV7QzQDx2ZZDPZRotTmZTQe+zwY3TUtSrCB
ia5bw6nM9k1jHkjtSSPDZ9st2SAdPtq+ntrVyBd3CCRUAVpnAW/2WAVtR9w9QBsNm8nS52lCltLt
udv9P1EcNGmN1GTV7IdDTxCIDskPLJfjQZ0GJxrXKCal5AD3UT6V3z3oc3kqyF1zXc4KpDsishiT
c/myrKIKh00eCbQTOVFfRCg4dm7EP/r9WVp8VzntGFs+IGte11uNmZ0ZZZ62Hoak8ShbnjmgbgK9
7Yuq8j1hiV3Cv3yLjzmLQl0WBFuT6Fy+fgROmOhi2h2S4FiqvlLHi27eioZ7BkoZfQtUlltcukPz
APT/oxc6vOK7ZgQnvEwtVF0QuYSjtk2MyYq4d5hFXWSPdXGqD5rf2VNesfl2X6bgnflagmUAxiB6
TLKO2cNTyeG8AFwd42hXBzJHMsHCG2GLuVbPyXQMztAspu3IXYXNBo5eUiGi5/e+89ZD1tU1E4/m
x6lSVhlZnNRJHAgXqnAPFXcRLXs4NM2JOVYN3tDcNQEGRozCyHIQiuYYlT5DJWlmYKYwCDhaROPn
7endX8AP9f14V7tNbFtmrSigo7AvqH1W1PIJs+i+Ag9VIdMeead4NnA2WJUnWxsjwWuv1Of9B68w
UtjupDEUqna93HcIxTdCoYcCmdjTg2jcvQWLc/PjnXAQUxCvkwxAKZbsmCJo+ULVRMoNO5RHGvv3
5euUPzsR9LQ4YTuoHe6wwCkYRgEPnhuh4QBM2oOKUaNYVhxbKe6vU3sTCHwl1qw1++aVAaKnIn4H
C6Np5EjUFsVcsRubSrkmNYaprm/I1sJhv1eT7m3iG8RuAlJJlXpslw/BapsyYMdd2erb3X1RFBQG
5TvyrmiT0C0Gz661ae1vUqq6i47LeJwRZRKPcDgtduSiX4oB3c2tEdYNSnz5Cg4avRJITen0PURC
X/hruZ9eOy4bQAYLGCQwjRSvjXnYfGIssk5Mg0tn2A+kq5tGZOX3jGELiyDcWAU0h3eQh4tPpv75
K7hnRfZrA1V941nihJUgtbH1+dA5DjBL2jYf/eAKPVg9n/xD9J8Qw/FhYU93sfuS17ofyKucEPuY
r5hjSyA4IUNCAzqRzQLNrMmleDa4yhlUNGJuqW/zQLrSGUP3sURBOtiP++RN8ec2knK/pTrh8Niy
hP36TJPVnvJjRumO/TRnvu2+1kw4kzltyF4MBBwy9Neotr5tViMwddvXhhMpP9xtajE+U2WDVrnk
Kkb077pO2n8qC3q8d8REHcQzuQgEj3CKO42kLTHcj1RVoC6eF+ynRMsLoebHsv+PIte5hNB7Cl/0
Ta6PvHZwgpIWRF3GPILb8HY/XAfGigjnu30mM4v/YY94eXnrOlxrHjH8MhK3NEBP6qaTM8zg5BaE
m0y7WAhAyE2YCKNZjqQ2Jmkml4yMCWmU1oFnlhGiUukUBncWNMCXvZaLcG/Obtq75nRhLkHj+N5J
RfBgjO93/rmJcBUnb9N89ma+0B+G5UJSjAPxQrdOp0jBbgZwGZYUx5SMNSAhKrunaSGQns8qKKDe
QBHu3a7z+sBs/ykkzt2iq9PsZFCpNvb60qhA1tu9bNXhf4B3fA7L0b+OtM+RvxL+fFtzIG06gXRD
IWLeDN1u27ZVzA8VjjYEyop9EAS6z6P7vc9rDN6zcepW+0lBHVNcd+iekQIIEzu2dYPKpZGuVls0
j2qvAYt8iI/v0vDV4MZupLiN+LI9f0zENsDyxo9Cetkv0SHMtoAadum5WektngA1s7SLZ0KfP07k
H3sYPNfELKst7Z10leHWvsADT+DBDGj/EoF7rqPPoEPeGVaFwKlEPkez/6n4zsf2DexogQw/XmtM
RGy5v59L2RO3varvUL4VNcM36DNitYMw4mdnerizjvZh50FzQ8AnYwWrXgWpb0Gr0opBEeVuArUT
+xNJxxorzx3fnX/5eljybeyZu38W3/5E6HDVOJ/y9NQ5/6cus2Iwpzm1We3QZ93hwqTt6d+xBGjm
BNUUQpLxeqUccHX9gih9gxw19e/AKcpqBpobLDeDd44IeAkfnIE7tx/VeVN8S/1I9+r0s+koVqNN
Fn/PzcB/yztYl+JQOAseb4vwr9lHOwJSQ5QpTOd2Wo2X6gkWQyJfkr74vLpLbCQA/6zrXio4nXYP
rur2oSoa1DTa2GMzWlN2xEKVEoGB6Feb1DxEBlpYuvobZCPMe9yfdysGrj4WAURFzoUg9SITq6I1
I1FbR2OIvfqzw44X8CLPUr5sUvWjqFMK+Al+qwG1cbbymf74fTdjfKp7fFtmBrjxpda1OHUAvcEN
4JecvHx0JDL5Go31cz5tarcGkAqL2ECYY6Ekhl1QCO3FzDK3dZWMUKgeka3x3WGMk0YxPEIijiCe
IyhxT75m/j6YrJmmvNtsR3ia0ifV/L8Y+0JMZsIOkgFWCgN4uLp/gtZ6hpdJsTrVE0TaEVKdMrlD
PAEfg280PCxEXRr0gh52IrEVS+ikyXkXgwTuxR8r/IMfRh5JZg5gZ/OlaH4AF28BHbQq4BT2TDW4
m+w1UuvXFzMq1c48X56ep9Lw1PuMd3j1C88Zdf0d32CCWrQPVTmePqQ0xW5xH434uqwrfyqt54v2
fw8jkOrinxQ8iy5vdTHEaINLvJbLA7my4HszHVLNdvYdeFyEv59v9nzS0/AJWLkhD820CgHPxC7L
6BKdWVDC9S0SjIPAzaCpnE2Z1IWpDcl8xGP54x7WgMOusCAmoXu7Iq8th5tNSdSbPvpPiAMgSUkf
UJvNh46YkbtejeoBfBXiDhKk68gdT+g2vYkk1XUmsMVV9kZj+7Bqrv6FsN/V7BX7pJMw4kgFP5Q0
gFLO8MLv5qV6pOz4nepTirXX6YZCbnKT5RC2sufPKNIOhcstXtKU2UFqPv36KSLtnpC7huoD7fzr
UjK5b+Vezt2ubuewYMY8PAFPOggXPejez9yZzcjgs4CiNKWWICP3qQbZ9nRju0e0w3qe5fDi3IOH
iPaWZaVUgGCFtp77MMPELMchHgT1CTlPDdKHpVy8OUQiviXK7so9iTxjpVq6xirC6THNMH7crMm4
VbmH0qTvsJfFkZj+/a6NKqBnVDRWdP3D2HNZ27PFrIYnHN/4P2PlluamJSfGQt66xfkSFCNd0+/j
WcPpK1e4OrTnUp89t2mf/9mxwXM2lHp141Du7/KHvmTTAFuWM4mExzVemmTaKOXRxxaGakVjxgrQ
EbUzbuv3TuenEv9pGweSSP8xD2t+/MVUNCu4xBPNfEkznoc5Kukz97gzUYPF1Rq94J1Hs7TLEgXR
0mMEz37IoCm/HNOxjzm+kVZIiqkunBmIPosoJzCLZ07KYoQL+vu359aZ2C+A+VOMqJahIQ+w4qYE
iZcif3sSGZ1elBwHGb+fOTY0WZzwNdZzCUyVD/1v9Ek9C8o2/+ZhozU14q3zuHhRb2g4CdoHLHj/
BFBGZEQqpOras3oCt1/QTIvrI+pLmo3Zll+Q46pdpqQ04/ejfY88PKHYue5OhosO0ft6yGdKwAbE
1dFM8d/ovQXwS/S8ijrc2x1hMeDlZSTT/6NsmY1CoY6n/+s9zTnrcwsczrff8ehqTRGdmWq8eKsz
d5ViiFTmR+3/ztxvIzRtYaaKe/UIoxQCW5QEEcMB/XLU/TttKeF+YhubjySEDRrEwPd41wVH42LF
l6kKNdS16eOUE4S8+AwHmqQZ+yk0eY2klrz9CaCU51eyEGVFvLLCpXcXdVjeKhEOmpE+W1jBTWMn
T93FrlZsF13vBtUYa41J5h1FboGf7MrIdAOVfl2QX0r2sVdwR+nHu+FDXCAVZu3lukJn/UrMLrnT
zPn/9c7qhFHJWKOFPIRiL8A1NGC6XqkAASZFqda0vNqyfWkqjNZa7tsygZNEIOXdzYSDBDRPXQYG
ZOOU5PiG82l/wxr+yEdkYCaMtlY15eQkNXZBuqSWpgY52AM+QoVNQRwGkabfBnHznxEJGgoZlSWE
G08XqqidwFIqdWOxm3t9wBjmo/JPMM3FxG7JEjW/Gt4iqwqRHBFrKVQ4eQEK+Rx2bQLockJdIzx4
Nu16S97HCrhPDRx35eJtp3+0exO7AGGxsd8KXye5+MHdiSGzWkvrjwLyDfFX0mYQqLSG16x0kGEj
Ri85NCsfLN3/CJz8wNFdamR/aDOYrVPnIuXvzJBjpXXiXxRahWlC+9ov0PqFgwEyHgqHOeOlhk83
9YiUDUFpH5wimqTxIQtja13wuXeCiLvehNHaamBLMaAQa1p05rVzVsRruG7vwEetghJadPUVSzjo
HzY6BEivlKXrcRcWJYZAnJYtmoFtT7VGPohEXIasg9Z5AZBIWdkrigYP+u3iaQXH38yJuASl9Dcu
DPA/iFqbHsRYU6FvdTvdExAXp68HNNrqxyuc+F85pnmPPLDJ7jBvRiwnoYnMKo9ZD0E9txoBZNHp
TXYFyCvW0mMRxKCkaNcG1Kca0uGQA0PDcMI5ySvFxgbaRsXA7v4i6ozGzlFU9k3fljZZBbRtYZEe
JAgqkjuJagyU5wElAX9vbOk7wnhibnLZua1wn+A7e6Tj9tZ3jApn6n5DU5MMC6chVSU0GwLwhcd4
K4pymL+IiVuWZ+w8rVXcHmZfS0qEtbucd5HhVE+qkF05FMnobdlyg3kajsz/9khW7g8XBTtYZeeG
anlkM/jclzuBwtRzT4kPvVbGPxtKgRuhdRO3Ak17Rds2FwERuNJX+BCXK3JlDi0bQv8O6UO925XD
+6AyOR1DRlR8m53FzngZRBLYfgFhtLhgWePlZ6PaFL66zOQdK82vUhn/FecQyPJzsA0It4yHwmlN
XxI2BmxgQnxvJAY8BBQAxbCaQsOmHyjWxRQd+U5+TVtRTvNGqtEEeORr2Tr5MOfORgMplIq5SvMI
Z7xZgCcmEhByxIKqcO1LOD43p1hszwCxZpzjWwozXezI105VCqGwbjFBs/NSIjlby4h/GS+X7gjb
rKDkwM+r/45BvTkMQ6vReMbSvCzgvESwMtHIcYVi32K3jrISemTSMh9L/53giFtfLmijYD+Dp87n
16ocEZkponRUfSOTzO0kobWTdiblgNnD+kICR1mwk+UXaW7f2Tn+0w7KW7T0Gva3wCJg/C+iOESH
h9wg27ZFkh/X0vq4U1W6KATSxWElfJZhFPhezeay2znECRaYk+oHOl+/tvqb+zU2KFjL9OX5ODsk
wJpFefSRr0fCzoWalpIX2Az4yHO+sT/PvXYpr8DXZjVOsENCVrYjuUycVhvckpONavMGu52Jv37T
FuOwkW/JG7ahiFgr0zxXH0DnJVkdxOPppckeLMSS03uLpJgTxtbZMFY1joIFpNCjyFQBlJLzLNW5
fj73lefkdvN9J07F+F5Uwb/arXS0QWSaKX0zVE3AQ7EAoBHMvkzzk692S3dFEfZgvBuu22MCMCuP
HdZ1vS4Wuc/HH62/hYhhcKEOpt7GNB/xX2GPgCyasVTa4MbdzBrHNeCXphxQqP+DURWghYVjgOhu
+vTQJLJmjqa5TAjuLA4FGzcy3JG8UK8gp8PDxo5yv7u8uluP7Pjl7RJRqzIAeCKeheTt/bBtKMlQ
WpQtunD7+UtAkbk2Qcso+/WvX/KmjREtuhyeLe4hyVf0gV0Sg8AwxQmEPk2igcjnMktCesAyno6A
qKS9Wr47ze3jgZJly5KdETl7UvucBRr+ACtXqPey5r3glEDNW8HdC8oWo+2FNkuZESnIK58hW4fG
N+YvvEXtgtCPJQpjp9xrj/JhlnKEbpCL8ofvqJlDxPTyEYi5RjV4q4m2YGcic3pCyxw8kBavaa5h
YFB9+Xt2n74Ll6hVyDTt4zKk0uGcM+AQNRx7/VqrckrcKPjnh+6baWjVNYvL9JS9ksW6RdD1tPtL
LS86COsYNX+DFCEc+USJOtCWSNbIeDYvstWVJvTRasVPrflUTR7SjLbaZQUXieVHVG/rqNq7tRO4
qt2MFLcepjm8Z659GKOXU2Ik0AES+VXrk3L+Nh1cyicxZjYuXAlrlZxyMC5BYOvZ61oQrrYTpkp9
HOEAy+Q3D590oWOpBtCyolNdH4MMIkryutXefHybHZ6+N2+c1BTQgl72k6BHuLe4jNXnl1SZAkWy
RyY5qq0zwvgsGEue4F3NRucu33DOITbdubyI3jW82se+kqH5vK5bCJOtTG3e6ddVkAMpaK1B7D2I
krrh9yQAhqNH+pdqoY+G6ere+Yoer670DywIJ4U/ML4qiPo5C5syy04f76X1suVLLZUQo3wnCFKl
wB4VKsXnPfGsaPSPX8iPDkSWYnDcMyFlFDPbg8Duf/xz5cS1KtYGod6cSRzSZ1Zf5wT0UQawYoLT
cldmKLIneVlZ9yW8xLqGGRNtvH3gMHxwkY2bwMcW+/1oypoubyKwbrHVo+lkFZRru83tSEw13q1/
y+KhUK1FhQ8BlZjppt6u/xFjgPz7yTGlNlU8a1XK4zRJUHbqff8i3SeCqWrifS5P4Dxf8FZ12r33
pqJhzE92sgfXen7FH29AGAfdhVti5of/ZfDkxgjMBbVkMiPywCe1wXZ3Vwq/d563X3DAFhT58IvP
9JsUABnPyFJHY9AcwWrFpaNTIbVgeJbBf9Dnzb4BfsS310UheHkc7b/mo523rbGSZVr60QwejRmE
L11YgWpHYnNHWDyWxnf7dSgrdDAqwAQ4zGEdnQa2tegQ+ahzlFnzpNoCbwkM9dvMKfAM3eoU+8OU
wO1kGRn/WPPqkw5fw/e5zGyuqLNEKMGsGKE/x23SfFrGzy9c8u7cM5ft8BSxJYYsc9yqckPQKyR4
PsLtCR9t4PfMUYXXoYsmMF2+kdw5ZsZs3YBBDxu68vqgJMQfGe6+KGMYPLXvvUOPAGz5cUU0Qovr
xpgsdkq+Z2Rqd/AcTRXzt5HlaFf67DK7caRuBNqsTuZfxNCCyotlif615PKxCWKPQKbcwGdE09Mf
MwmHCxOTP4YxDBOMY+u+ksjzFOEHaXKEAFp/RU2zpXSmjvskLY9TtQAzjsOnLvtSQ0fZ/dXPAx2a
tI8smdw4xP1atfghJVaV1xlWi2KhsBephiqeIg53txpd+onusA7pmErpAU9Eqrd/9yeeFjw1x/ji
sOzhUbF6T7SOspTfm8NkrOMwMemmfEpqpRPis3rLlIBblIsaTiQBA2okaFLQZfqhjh3CqP+xJOPH
geu1YkQbX3DrgEr0duC12LCKfaT1o4osgOSsrfsc6hwHK7qyxioVy5Man3Bch8DPaYIi0L3nUusC
Cq1Cc7Dwni11c0615Qk0yKufURc+R7dJ0+j5V/aNBmNA9Y1ZmtopDEs4se5h4is7LDojHz6LLeST
CDzc1dhZK9wtzE/WE5FIf+Lry6ZAjKe2SC5OFrvIY1y/OSVGf2SWUXNcFt/FiAino8rGhJsZ9aFe
f+FQJNVoiiaUhWyYEomZFsAHeMmNaKJjQFEezQBfZ/Ffuqvauw3F2tXPINYldAGpyHsnE8rIwsqS
IWDua6K01uXeK2Np/7aJxBtR4dxOcNwE5t3mLlGcpEEUjGri86OvArsoESPZaPi3yM9HXv5U46GJ
L+mYh6qIMRDso72mRjNQbjQNhInIL9ob2+wunHrTdrXXShtTTClHX2rsnMEvRsbPTVD9yHOZfnME
ItwSjSPFnZLUAjjQEjjZOkgKANZLlNeQS0/UkJR+Iu63MF58wfMhcjRVST5FyvbjGcxNivm+T1dj
QlAIoMEpy6/PwzJz0terKDvGDsZT0kwsSte72043znWYgvA5JHlALbFfkg0SXvV/wr0oyOSnyEv/
6GyC1Kb+QpWcrh4vDsH1OOpelDhKR9Cy9QkkJGJHWij6aJIqmKDvRHx84kxJq0N5I9CRTbaNuPfc
/ZzgJ6NtemlEzrNFs2J9+j6szJXBoGrn4qOaRk7yWh7JaU9sqQvGtgp41fwKSNuK9xyVXHsXLt4j
83o3YfpjThlNsg4ESf2tE5vK7XQ12iEFi6f6PMUdDATFCvljWAx1sDlYA/E8fnEbih21by/AxO0D
62taT0a/qDYb/0JsjVQk+Ki1vDJT0TAd194uLQuGnftsaHNnjEq+43CmJ6D1Ycs4biYtdOyolWeb
Sq7TTIDZ/F0yRQYc9feXjpp8h2rL87OKzpF2I8dD4gJT8ivjUzYQonLCfznhzFhfWmOW42MMxM5U
nL5RcvpL+qcqYyGiuyfTwp8VMhaucjGMcyhEg/CSU1v1T0UbeVgoMqcM32kR8AmByytK2AnHDP8y
Pk46WbAKHwly9aKAXMsB0RGkewmyAWgYJ1qTBkUD7skErbz5duHclUTAel/H51212Anv1tApVcxb
JwUlP8AoDgUdb4Mem1VKzs7gYSvO9SnAhX7G113Z8CQwGMfIYjBwctLbJ8RmjUdfn3wVfx2mFECL
Ik5RLbdhSM5KkHsB+c1fUGF4Dga1Zj0fJ5caRh53BxxNHCb3b61rhd5duWSFaDrkOiIDV3F09mvR
vnePaRMkAXHnZlKE9NaE5awEh4wC9GHcWzwvMDIhAhDFeD89IE+ZMfXkZbUgYsxf32p1AuuFDB4R
UEp8lRv8N4Hmf6vi5ZtNOfsoDoM77GSGYCByhvT0o3T6917sP+eRcJiIbrU5ZzAi4UgQETGCQVgw
JKnno0yMKol0xaAnxBsVIGlz0df2SATs/pxxpu7scCznQt32o3DVXY6Eka68MqRIhbXeiUctvs01
gdImuxrkfto8olpprbeTWaq9nLbFngJxjNbnp1pkeNsERIt7tY4N1/zhTMnC2rnBXL+5HdgUEo4N
ka0nRZ2gihmSLLaGV3LrbqeKlkLe2G4X6i9WzDmW6TJQCyvD96hisZDG/ggxfwLPQVQNKRlOvx3V
dDt5xu1GTfqbXfLcxiYwtjHq6ysA1i7xYAA9ZMHvIX2aBpBoztyF5WX5okhmsjn6b9MN9la28dLS
Q8eH+c/g+QK26TW41Qq3swbPyRr5SXTCwHG69/i9kWdpgWnBtbnJd9PI6Jk9EFYDIpWYGqDEO9+/
qzpM30zJd487LinZD5/cU91qIbFLKiI+3iavQ2wQM1x2danN/SdUN4NS5Lh7gxZgifhroZIEYCjL
2cB3Bxv5E3P1dmk6XQG5mF84fQUCMVl1YWXIPUM5O+miQSmj0nOdoqPVOtygKzPY5M3wG6YNCFsj
GuInTvsoL/xK396xXiIh2OQOEQAcv8TGgg7MtnvO7HjYj9f1/Th6AIAszIaSuy3TcvYG89SM7Yay
1hXwZyRPYRpFme8+6tTbjIIdbMFtSpIFAmOeSUh/TzK2KgELkc8ShuUe6W4PtrLJjy32ZbqvAzda
yimqBn5IUNxGFGC6NbjX13lFjI5s15dKWlJ/OqJEjIdaIWKakO6/fjEr6frCkwTc8mGstKVrI/yE
oM6LAl0CEAAxujcPGpl4UPdJPKMzU4Lv5/TQ1XieeanOt/zMPmjILAFIYWiROlJNoQ1YfN0Dm5L8
wNa6dEw9ddM/ExfB04A3rhixgioosbMFkvP6uVi62mvbovAG/9hKGVryT0OMURxEseByazZBgQNf
Sh0hkh0g3A67fUAwE+RUvVAB0z1VipHQt/1TgYyk8zBQPfmTCo2mzytPJWjAzDLABfYMr2rxLfwf
rG9Yzw0/5P4DV4Spa9Dmo+KHDcE/w/OUalQVtFszyeiEOK+9q+qWYmWSUf/qidyU2EYKytt3mye7
7Zl1SJj4G0MuFZQoQSQ5pUvQJYnSfVk5aSpQSIMpJY2KWtDcBuQh26VWmSUrWQqj4UrDxOZvlURc
PzBunBPZoIc4t7UnQ0PXR0rJsn1JfuW/GXXADNhExy3MGt03Ezvmw3s7M/3y9pujPPD/kHdQ0xtp
a18SwrWvyszU/FOBnofOfpFvFd/UhS3TUmPnQ56azxX0bAo3wC9jnAAQtUlTNyOIAdc7OOdbHe5V
keFonFouD4RtE6appeXA4Z5nwHLhr/r6lm2hmkd7BVcH1nRB5TjDKUhiAPZsXkHmbOUgJIS792Xq
CZcuCsDCf9KXuuaTE6iuP+L8wuFxYmZbZWxVMMOBhNF1s0q69B56bX0mNfNMd3QPMBGhQ0ao6Pgj
avLskF5e5j06e8o5ZFowVlVdq+HDJmcSmFSKQReXE2/bN4TgwWzUZsob6UYSw1r7uB41Q9ILCJWI
CseRAOCB9a8fTPiEN0617Zf4bMRWVPjs8phnIb8L8imicJOHltlsgPAt17U8Vdo0699oV3aKbobk
H51GbcL8pdUQCrwsUGQqcZGK2ZnqchQWfxsuCsCZz2BFSxHLN9c3vRCyaWPAhe54l2C7u5Cun0VN
Cr00zewEpxYLgT1mRbgg2UlkQDCtg3RdrObxDdcbErys1wmaJySH03Zz/F0so+XMP6YOFuaIonY0
aa69SZ1jaXQuuWli8Cz+gqL4dAp2hzdmz2d6Y99Hj52jgXB30BVQqOvbOhmQwRUAe1F5el3rwxBj
owmBNaI2kWNmbmTOlc9ELOlsV3zo8JAzdhy4WetzJzXNmcDs1x4U7inPLR+k6u99jmPQsGnQLTss
r0tQg5V9n3XYwtqfae5mKKnSUKvBtTHW5WlJaFefUZY2uVTSzLSdndEoyAfV+4PkbsVyo9HM0ho2
XlcFDLup7RAUeTcXOtmb2hyMhYUDt3Gkc8giKtr9L5Ct+8ekJATTcPRrmV4aqcfcfJYtQu28hBvK
v3OfAu4r8L7Q9dO9ZkW89wX22pzkQj84fo4XEvFrJSDyMQxD5VYukqXdOmdot+g3vy8QSYQn20cw
78vp8TrINTo6f/cBotkp4TmmRkyNkItUTnPKmuvmpzjXauLsmG2pfUBcJCGN/XQqqXkdR/raXYv6
ItNCYJoutm69F1BesqS1WYCBxudkX5urt1xrRne4uPvU9Ez8FO2fpsunhwiwXeW4ETWxQqU7mupB
c8MpGtxyZ/Ld8HN07SQUgXD0561/rZ35YxhwCI39x/9xIvPLrkS6/FDyrPCKWJ4Zxu1EPgUxNX3I
T9FcQqE5531xH5UCfyWBx6n4RcznPLtJCSdmi1G8FQlObKpxkjJqV1cQNZeFh/6FJ1OzQEoc9RMD
KQOO6PC23UDtRtxMYKlwboDoMz+0/Gd5Ml+XlvItg7jZCCkXoZ3Y14LsUuHICCun+WHOg/koaSex
NjH9oDxoFDzmvXCg8DekVuC0BIhqVgQsocLwEzMlICcTj2RL6G70pWu83r1RKQ37n6wHlo6e38nP
m4mH41n2dTrhEMmIH2v2HnZZEXFKTWo8y6z1NqCxxQ8iVXwTsL0d0SVK0u1iKKA5GN0pudnXAOe0
UYTB2QNjLMBG1r0kgAoqmomoVnt3K3927gaklmRV3/hQLAeiliV9WeVn95ypkMUlmeAYit7Vzkp2
XSFHPZgoEeWuv6SIK4wVH3iqlM/ewoNfEOCRq/2l/eGenYjxFRRzfz9BAdcHRQ9qmbpgT5uTGCYz
wqb+gp5RN2zgoL6odLMDrKLON5v7TavgbigctwIQLu/n34X24AHTjm3KvxnWP4kKbQN7DxCUZwYE
U3UHL1QlPr7iKXmrp+cTQU4yi/IIacY8vrjYQch4Bl8YtfkhOlj3mBTVm51zrJQpyhMgmS2dxhCJ
lzQDmtAG0Guzm5xHmttKiFaGeBKvVrpdm3cpYOCsOjfpy8Q1cY06o8mKDrAaLl7r7LHQtuxqMJvs
FyYG1X6y1eqUoYpb16Ii3fqXgjxhBqlF5L+S2zH2WspVe0Ic9uvPyumdUpqoIT+p7LX+/xyxNpzZ
IycMmMXnQL5EMntJB6V20DzDse6i7G7wuINEF5qMJap+4F223Kl0aaeWZzs9T0GzNJW2N8J2ZBRv
VXWxBOqP+uEDIIV0N7nyqAuy+pAasizHS7Yg7k3HqLQd3Lo+zXFkR2sE/Y8WXe1z6rDwNJJOLq5l
VEm89/x+ubtZ2mDV0ZLTk6vRf9yEws058bADa75q4BJdvdxMdeIWzrdf9r5OLsXaV1STHk+++p87
Gkzc+HNlqhr70LSAbr2y+7O8ktw+WHYDalkke7QXQwDcFx2eQax4TOhosQepB/JqUIwmCL7zi6cD
dKU7Ms/mVmXIFxI01n5NhdtohRuYPRQKscqkSa/86CjFafO8w4UNSuGszh3027uNzYWRbnRQ4DkF
9WBSdeliX4lz4YirN1Q98yFvR+VCt7Vvf2J/JTR4hRq44z2C/dWBIV0WeihQu2u0w/2yVDijk6Ys
RYuu9yNDpZu/yNIkJBF6d/R7P5wUNUmTV+fvGFIeoZstrMhHPiQsvsO6tcg3ZVu7Kn7hMJPiTMxZ
fcMSkkJKGqZO8GWczKcsEPygwr+GAsKl0M4DcmgRbslp/0b7YTNUF5Ky1lAXInyyHV2AB0czOBfW
TsbJVFfhbIP4qdxE1/l90mYMQI1RPgoS+74Fzh66PvM+lMh2bDmMbAglhu2SRv+2BOMP32MZFcD5
13t/N9MOV1smTnuUoSKOa8WMFevig0swm1Z7v6F3Kxjxij/AwNNErQ85mzWLP2Tw0dAtYw+TQFS0
ha4KhazHOAj5BzVnnZWZA+D7MANKyR0+6uoVI1T0JUTN8VKtW0HZDr7WKF1dJQU3YmWM4iLCruPE
KKmCgK05lteV0JEFEJjrZec5+xRLFsxaTXt21RmgxtjlFD2ejfvQl1WDIZjcbAsuMYOMY08DmjeU
6ABhnlM0KBvm5MERxCOEyABpT+j84m6CGCIZVpAww/0/pgI3WzSvJGRXYR7YDAcOmv12qjxWUK4s
1IVedWTxm2YYUJbIgUNgxpkHolxrwOYwYPG7dfTPqrj6qTgerL/wVxYAdY9Q+ejpdVsmNsgTDUNm
3GWL7Z0M0/Ft+cT8dJS5dY44cXzaxDflMiJZD3GoT+pWngp74ZTBIe2+TcAgT8bxPWc8OB8iH3xi
3wjVJiq7sgYBcbGFbcTylX+LoXfy+v5WK+ryAEGcnc/zvkaO24AyyzMd00jrkTop7q7BdgvAgLDm
kG0HaS7wRxYtkxEb6DiS6zijK/4mKVGKEjWntOsgnULHa0M/E2pRtstueCy9/Fgmpq7+dE213xSo
9zUBb2QrM31ZjjbshPpEU/1z7GIrNlWrgx6H1VrdCZ8L+gkelfwSLqOxOs8+vl7wB19kcx8Zsh7Z
u0lNbi5f1DvEWm/OYXRcRh5i3Z+SOazHiea4VtLkAF3ntqLdw7E/nwd3d4k8jnVdWIewcO9VA07Y
tiYUBUNtWf70g0+CQnwbodzfnqMx0I4Qp/we0WW/PVnm/GKdZvlEwT8lIb0dhLgZjqDISBB5FyYR
EOn00FDnbhx7rH08DAs/AnLBx69YB5II3RqfIaWd9lTbTtinNzZfhYJGoty0gqli6KFPUabzWB9B
nkpMt2iTjebI44SMKhStDf869rPmOfP9XJ1Lb204B42aR1F6rPvS1PXMaEXg/XdaPqcSx3H/1oNi
1SWnyokeSidL4VKzo5k4Sevh+FMtv1SF87sPQKit4JgtadOUv6/MtSg1vmVYhL86gK+wiVg9NjTx
oKoaWxL6SKXx7GQeVeMNyP+L2Zzl/OvXkO6WaZBOIG/Ze53IZDx5e9O5WVt9ZqCX5V+gPShPhHT7
BZj/+g8IKjZlFFfZWCxHJ70Ce0wQ90RAeV1WAoLyaMOvN0RmeDQz/jQBrdo0XsqOCx9fTFMb5iIh
yG1YQLOoMrGjWCe7Oytul3azmBHxZa3el6CR2ifYKBlLUPT5Gt7Onv4uoyXt/usjNExQKwskAkaS
+Mnv1tGHzpGB2nubJquAKEWoE4fCFY1KVt26fC3PSDBfRg9/52u3rJ7LlI+TsCQoixU+hIUI78Ge
OxAu+3mbgkVyUcOTHGO8He0bYYFD8Jshblz0YJTDZFOerGzDVPsWJWSZRG8m8sxwzoMewyxMXcv9
u9sWkCZp1HDCupCE2aQg2XdmvfzNFfXRQXX7FuN3btJEmVlNchorgMQklSLtLIvRy5zQpbkUCmTB
I9iim6oPI4GDkdgOLflee2olqPyDOfWCV6KNsbopELLxLUW3t7mtXpE5Q0qJrHOUsjR2jH24w/dI
+yy4SEaOnC+QiuZ3k1t+zgUPT5Z1boOODbSBJUfRWgEEnwokV87Wk+cV6TY75QIg+T9olZuVP5+y
ugQcm73fqCMBNilSNzb0rrJnGmJ2rjWSrH5j7cO08Qnu/MyFJx5J6HVpez+pNJlbYtfWpxzldg8Y
uvHcEC7C1pYfuJ2aY9n0kvBjmJBdpByfWc7102CQDEruQc7AgQgs/V9s/aS8/mTcI9n57F835nJf
5+mrz4oD+d03BlKATcWMn3hsQmashSlVEjKI/+P/uV6cHPvJ/aE7S2ZnSmL56aZRQW+FdLCp9tpG
+99Au8Ax8PpgoG3wb6eqgr98W7AJIHRedbjQAgVdwN5wSwm3AgR9Wmb0+LguLB3VZCfL1+yBqmm1
yW4BNpMqB33uxNi4QaKZB2gqx0jDBfrXC/HUpCaYMKCcCrBQ4IJMBGCAkYfmlutVMSWVSaRKHl8w
xhuJVncNL+HJHS4+VVYJuLJwsaRdJ3W7eUpO/CTWyI+mfuxS0EPookfJlMLjF7ty9wMRX/RTGuPq
0dvWOpzrJTucveOVwsLAr20NDvhBrOSUo8Af6EOWyO51ZWpZ2XgOGglgHId57dsU6OMw3IXgJumS
N3nfuaibRPcxHMs3H2MxYtfFxU8ui8l1Db/cy6FnkGvCx1RzArZS4tFaeGXH0nIjHYKEKr4uwKlD
0DeJjHvImQLqhUFtzGOWR2yY1H5yJp4Wl3RoVmieAJX2pH6OH5E4oOU/TZ1s70xkf27MK9fhusxW
9FZYP+xpLp8bTEs99jeQGmIrc/phPNv9FOtXWMj3vOBXRxBPCEMaFPbLQPjuuzYh8FBzOUrbNbfH
JDoGxW8iwZSQq179ocyvg1Fb+nhkiO9gU5JjAXb/KsiKiM1cPe2imRmAaKd7JfVRrfhfS0in68H8
Sz4RKB35gmEiJuLsish9zXC1zcqMmoclHj60kajwWXxCd1ZnBf+KTFyCWJvhxFQ4JFh5/+LK0oXx
JzgcbX+Rhaumk7+O19UOooo9fYENQicEESzWHY0w2IE21z0laAR/ughQvUbY6PBzvO1Dx3TiU5Ji
/dvIlOiWHhzZeM9KqniLtE7EzKVaAEpTbXcL9P4YpIyZ60a9fXLQXE977tgy6QPifQPwi9W7RPFz
uj0llX5EsFk+sfA92WEnUAi+EQEep01hizqlmvIb9x8NgwkA+uEHb4GNVjlckStROT5BnC/BskkO
KDSi9OeNe1GUiK2sbNTAtivzzlDkyvu4j1UcWd5GRhNdynM894DTbOkqjcN3F/KbOHmIC3OhFB8V
3H88Sf2xgs9dv8zllscH3d+e6ewDQg8V2hGHobe+rCKjcYj0Q2xYxWMIfGaOKH4CW7X9j0FU22Lx
qMrjZYP7YMyr2NtPaV0GIdslwudLNC+2BfCqvt4O6mz/aNf86ro/KlQgEJibPrQwZm8BNFA04NyT
g/K6BjGVhR6AOFzXBplhFqTYvOepCmQdPk1ppnG2Cd8SVR2me8DMhcIvFPoa+x4IwGKcINiTndXk
ttupqhwtxFv8X+IuQmkDhwe0hxM3JC8gi4Mp4Wm1/NxoSpj03tQOneLOnDVOWT2dTsTWunTZ4LZM
GDpJg3s+LxUee85ADDN7I+daTmjkKqp+7bdEk+yWSI2RtR2dUnuN0a6ZJJ0B9NdSX7+jmmjUdSd9
TVI3AU4UyTxQBWeT2Jf/IjuFZb4OBdN40YroakbkQ9DngxV+LTFMUqi5AH4UsRlbB90Z5UTihoRc
m8o6CTn9kH7+R6OeqNp+Ya5G8FwPEN8iDAz34aiWrWNacffI0XKQcbqMQmYYPmynJPBx7YO2ThTm
JYeY5BCHqS3YgzIPiln0mdVqGJX7fLDFJ0Ud/6NXLLgtDidkgkWUckKxh5TO0Vi+SKwNruRBgGLZ
NAm+y4CnV8QovvSQNbJ9WQQGputiy32VGV0RvZgAZopuATj16KMDYK+AUIxbwB5DJMGkRIf49Gl/
WN0ipYMbTNMhQ8niWFGiBaJ7OliRGAc3GUdjBU0OrTx6t7riHacOd/4hp7oet8n088HuP5LDgH/6
8cwY7YEgjOkSFM86Eu6jnW0ipBjoY8LHZGuxGAtrzjBf1Wn8m6OodOR1VHJZ5B+IKWZ+BAMHj7eQ
oTQ+CU01cCiWBr0TOW6N/JuO66XsiQfAqtMk5VZT7/cXNHM4FR8e/iKFo6iyJFsB7BVjEa11n/o6
1y2PNmWlWksVMBUfJct6AAOQqjbtNwitsYeSgOb6GU14ayTFiBme1YFxjA2/1VRxcqIDX3rgATjY
gww9+9DpRwB36Y13h/NM+I25q8nrG8tIhNsRWC3ytXGJY5lRbz2CtBQUrKbrxUomkkbPEDFuWnXM
uAfkpKDS5Fr1fTev2iFIZI7mK1rKGIH0QCv8/f8KvrxCh45E+ro2n7ON2s+Bckh8a98KBbMctY6W
rreZyqOwIyH3WoCu32Hrdr3MTlP6jbv2n53OpLau4lRk1F2aH3Ui77W6B6Nk7CaNpxhEMzVOgbMJ
wWXDzF+C/FdS4gHuOclTHyKVjb8AnMr0MNIxICQ4GhxiIRz7obhFTiNSjplEOwcyLaH8AARtU7Ak
aZQYEe5X0PL8nzJU9jhqInsWybpGs1VXZx97GM7N6RBiXi5/cvrbE0fOCevx4F/OlbTzMY5fUbhZ
1hiM9SNF5wxyOJ4d/E3jRqeYO2ZjFwhBkR8TH0cYth8GM89xqerMsRRLd8DgbUuKo0Vbjh/Saqc8
Ja0oB9r3+oZkCMDgcRFDxXjXNYSWlmMQDPqmJO7Ydd7HD/ng9zdyOMOeJx8MczzQVN4eL1MA1kPm
VqwExY8yZbNeIDukEfzmjZyNEMTzkwr6Zci8xBwXBwWxONdDce4g8RWO3FrjAxFeKtmYkBlVqYbP
M/y6FAEEIICAv423EeVm88F8micZS8+ThtakMs7T/nMenDlZkNK1pDeZ8AkponIMZbrRB2CL2v7O
aNdeqbscxZ81CVOmScMNEmQnkLPo/d2UYqr6N9i/EbJAKGEG38tx5DRogxsqo4jAcHiNK3vWiHMn
VHXrER6CTiayTvZYXc10+jHORzycYgyC7UL/MEjbIw2d2DVSIHNTnN9yx0yj8GtorPbmtRGl7VOQ
J5ujEtvyZMl/laRzDU9i/pUVzzJ9vgnxyGMWbxghgzBC0/WsigwCXwxvKLv9CcaOVokqv4AsEg8t
pXO/e52fQ2OC2cR0CThDv74Euh7EWNaFzYZyM6zmfdP20QV0tM+QmsAETevfYf1tmMSW6qYZxUf2
U6UzLkJR0kJs8WztX9MoF3csxQP503M8Xy8VxvKNk9hxGBRpPy4/OsuNFoGYwjmsPygiEeI34F7M
mRsQs0+O1hSzwP7UVxPpeZE/Vm2lvCrhn+OWMUAt/bC14uJPa+lXA6rZ1znZUlSJPLmHxSnW50yP
Zo3cup216iO1oxJXXyvOEv3ii+Wv9pi5yRiy7n2S8JHjO/jQaS50Nt3EioT3RWtND2Pejt5VhaMj
lHRZIp8wgEUJswKVfVZZjwPThOO4Hg1XUw1kKasRPYXMiNFwYRM5LzUuwFyjj8NHsICE+d5lKv2i
ae5Ay+Z+iEeStMHqvHQwGYHeQoWAkuuOIg5h0b3+7N12FGKGsdNvnO6l7po3YIEHwHDWY9zRju48
bdvL/qvXctJNhrrGwmzbt+Fie87j4Y0ykC57g8rLqujPtUzqf6mDSnMGxcQsp1xAggF3+1V/c307
DQprpJSW6aqEhpRTQcTpxvgmJ4ArTMqaNLBF9/PnfVOdvl8gX3ignWHUjdMB5708aSwTsFsogkSG
lQS7GjpEkCAQY7N++KRLk07WK10KQbvPMIRZrXY63FBHEcKlWQCiHd34ZcGmNCIIjIztPZIm5Hx0
pqBUkUkaGi/BjdTMJQVFKyY8oVfzTFMVts253UZ6F/8Sflbp1tp2ZCsIS1vMucj6yxK05BOGF2F2
1bcFY6nf6LYsZczNog1Sebe5h0cRPjCLHpOtWY5UxbNSnz6aCRpZpCtSNzd5EWYSnla4dGy5fou0
W6bdQR8CiMi3lT4luBJdcmooSETO1ed0I7dV6+eyftVn22KyL6pgXFIz/14LGm5fPYm2DjDuv8m4
vxpe0n3ugJR8lUGPnyutMtwU1sPEDidUqH8crI8KI/rVVkpPlEV8WsKtpBv6KqUsfBoNS/iqbvt2
X3grKAwnNtUZunN88k72POaWh9QcMXFh57yWRmT8hNVwOaJDY6TGPXojC1yG5fbgy8qmmbydMiaj
9du6SAOx2Vm+ozJ86YIHmsbkIh3Kn49gtVGeSy3/nYBMi6UPxFJb1CL9/ZI+MaXOn1C5jB7Su40R
AcxWJyRRnwZAk0DAhpOAsgISgERyJQDZv+8Qug5pJQZM5v1bo6hCekiZ0tqidg/Wau0bv1pG9Oys
uDmuTMIh+GLhNClRJTHtmHnZyK8KzxiDL3k1cTMF5tBK3lOP6ckeR2vEVT/BEtHYR8/W0iw1sMD+
1r0LmSGjSkJs3YHj3kbHwpz/wkeiNWZ8zyOi6xJuFWxaxqsJud1fvPlzBCfDHWtHHg6gPLl+8Pph
xdk+jDhw2lJO+u0GzTzWvvrOgkeRc3D337i/r210rSiaLBCl7Y14DJfycOYH/rtAb5uf4zTqXtee
IHuxb8CW2EbRxucuvvOyjd3dtoSgpZpwD4MqMH4gwrdoWafOydNYoGvzUYtlTsQ1Sm7ceXmMx2s8
93pP9+IReoH2VbESXWwvHlNchFp1thmMP03ZzwMHnfBDBFbzJdL1p9EYKE2iRx/rglygbLv1ZEjn
aQKWwBYEopuudmGaQh7eQuCUmJVh2O7zJgqpO6EC0CM5VTca7L5vHDvGKBFc0CtWtTWdZAHAqrin
dhbfv6MH9vDVNaEK4scC9pIxrYv6gG7u51XltDwHb/54UMHgAgj034iaPaYwU8l7sn/+0CNOjJEF
r+PnrPudd3KU5tn7Y8izk70UI38fRNqHPZ9pNQIyaJAOKWwpdd/Ojjg7KrDck0DNKcQaYK1o70oJ
XPlgVqonq7xGGRH/DinIA8PMI4ke9W9TjozExtVcWO5gGHJt0/Q4vBIC6GFNWe+W7VhjDNct5R3F
xT2GZuiTzXs0UhAILxha/cGGi/a+EKCGbPbT2f8KZv4Hb1EF0Tcl5xt1K3P5waAv+yAHFG7uET9r
kMEbr/ZpLLWJIeeNukNI8a0gCVLQZYhDqYo/mlOdnMfajgexMpaW5OuQBGuv27/ZK7LVStECfFSr
sZpCAM6ZjoU/Ezw9gPsAmExPfvQAHAC7t2HF07Jrb6/joUGzSpPFcTK+gds1+xkptkqSq1wu0pBW
3QHTxmKWVf0PRtqW/VKHrUe/Ne6L/rqGt+04TyoEFD1gm7H5iVl8YuEMurKbWlzgPQvRGBdBOMxe
iz+NrCq/v+Ap4LlzOEjti37dt+8ShpEugf1QJ6/YMieDW+SKbxiYFPy51zYyXVwEiyWMqFuc7QmA
SlwrVlvgPWAvyyoXyDGVyB2JUExJV/8P6A3zfMIe4qf76hMGjs6da7lbeITUCW0xpDuXsl9GWNgn
w1d5OsQgXx8SNJ15CRkCO5QYBJrpBwxYruqkiW7KeS4cWxBH2YgM0ckFhAevZz35zAMpNlrskz4B
syTxTgNj5Ad9RlWhuIQfKaKmbd7Np4YJXjw8tEskqVLZS/FII2RFIh4zQXXbLhUeuqHvvowWz7pP
tgNCj7hQweEYesxfF3kYd0d0QaSl7T6TfIYaU+Xtt7Qgi1MYQS1zosQAmFjknn17djm0W6QP8SzX
VxynEji26KfJEoNIh8UnihuCfK1nrf8Vf1er8ThN6s09pxhiaq2AdI9fiUEs+eDpMEG7Ieoh7yIJ
Fnd3Ar+xFufLy6ssW8R848bbZF/zjsK5eZbcl7Fy6rqH60uk8dMJY5LJH/EDxgWluF6Vy/0qTY1M
JwUnqhN169CxWCAL21YK+oW0hFGgxlkaYudlYg8LTm4QbB25bv+Bp4gRxe0Wm6vJMpSPJaK7scNN
6ddo545goh46d71POCOaUcZDI82OHNvThMVsKK2aC2QDnYFH4zlukcSSq8HS6lgHJAEHYGOR7+2L
NLyy/xrFREae58jmNhwn+/Z+5IRbWlzho9PcMl/Kw0lNnXbDEKqoNTNxGkU+kHtEzE1TouS94IXO
EIRJpWenyZ4lH1/0heBTslMIUCI0DjEgCUh6FMbnbRsGmJWF3NSQOsTPI8iM23E4lDXGQ3MiJWX0
/RpSYlocY/lymEPz4XNO+jCWR4XrK17bTFm9w3Ej613WEhWivoawEPu++R3soWauvSlI5/iH+RaV
aj1AQ7XK5a5jG0rirne1IngWV8OrkA5IAfAcKi0jaRX9Xzm/E5t28HcZkq+3vhdhd1YoqkG03Tkn
Tbr/bTmGQME4wf38T5wMD0R9/CZLm7K7W2d04gbXkfD6bw6uQC5A1ft2Yy80LtRv8y/rEikI2trF
sSFvn6yaSKHD3weCSyIFX1KgzaftmnJAI+JnG3nJ3Zomryp/G7tzB4Ok44NeApM8ha3Es3qVBu5s
z4O+nPgrblbA/3KsU+y1K/AbLWgAfRkWxGctx1hgesTLwL4m2Md9Rqh2kuS1zcrJn0YVe1S4pfgP
R9QkEBhBJ9FkoL8V7z1AIy8nJ718RzYyX3T45nXPMq+ZlOF7c3j9S4a8ZEegkzdETujWg3szpL+Y
Bu+Mebd9W28QPslWX5DaYSHeD/vF4dU7y3yRvjwJiVaFmtSemulxcWXWvIrpL4kADcGa37EmmNex
f3iEZ32/vnzEzQE9mQyqkysJp0tNPlUS9cOV4YVV2Uir1aBogxLy6aiP/e3q0R2jDsYexxIABTX4
VT9OOhnypLSBC/HEO76tgTnAXuC3v1/KVFx3m8jkPLFJDVbOTdPcCdevH7HCxAE2zPJeeCRJjCsw
cyk5AfJaCItjkcnkibDU6M3/G5XuEjaVtEr/Ek7+v1rz8qZ0Qbh8kjR+gXzUNoZAaIcGN+4p91p5
pCy5QlgkCE8HWpexSTDG2V3sxvshQxr8W0+2sXNe+AdXdrLMwEshcgd40lKYaDZEQpcPFCuXAwKH
LZ7serQ2O0eo/6hoMg+9ek34id9CTtzczfrZkrVNpKzILlKL9p8NNyRn1IMsyVBETOl0K8p70qSF
2YrzHcpPNNW+W45fLqYBmhUY8trufuCOFjWp27V72KpXVbp03bJjNPIs9/wv1dt4xgwQ7XEEc+yl
DboFTmzsdcIzIuxAltHYWKrEaqG6RNUgQwWFPMwhxc3fslE8lEnZZ7P6iaFrrsyPsPTRq/xAflKX
A5i1n0kh45jPxpq7VwvIRnzqNFZKVLBct85AvNaG0PWilsEnz2HWV3HmSZmJLew/Pt9nAc7qTKMZ
rcTDnrlhtVvQdtm417eai4NGYy1IyLecw/BAWA4ShN34euZsP1vzpcKBPlpuWcc/0h00C5mjvlCt
mS0V4wSWKHV7JQ/b3BZgAq9CU9E2pZcMIeGyuGXj2hR8PduouaKBMF/Y1+U/1AWoXbq+eU9INBFT
S7R9sPEGGiCSNhwA703YY5+oBm73rsrLVN0sqIf0c8IaRPxZGi5F7PY9+3daGlLOxRFqz7c4xgGe
U339Y9E969SiMGlAOMepzXc/GspBw4xNYBnKtWpxNguLFMASpfIMIoT9M4NNOy85MQt69A7AeRxH
+cfjL9KYFNgzNtFtNRxp5iQNjmFQBW1qeX9fCNmcv1yKdG8yAXdaXMTt7zsVqeCmJ6j1fP0GLD91
QHK4z8rzWBGWM4hiPo+TRzs/OYsWi1vSsQ54W5mzbpWpEX4xjhDSuxef2AGFp34KLL9VT7F5RrSw
Q5rcunH6SpZb+R8ijfY4COhyBRwNQBR/o4oYKhWI0qiSIgwH/nj14L0lLAHxCDP7276Db5S9SBOB
aDejOlxK2H3wQgJG55BlkWz1w59eZkjDTddsW355g/KNe1WLz+xrSO5Za28b4vAt9BjqdcBamcIt
e4/XL/YK6IZr+2qCMBZ7anZDAwF70GZVv4PuJc/A18udoS2aXLkpERSaIFyGn2dl9mD7XlXMf0TO
0ugkgNtwo5g7A9ARKJ4oiUGmrIeU9UHXbSaeg4Z47OjpNxu2vkbefMCo1gJNhRds2njvW/bFm5W5
yLXpmvoopjCY5Yq18i09Q3bjNALCCYfNGtfJ6YFMQdONna8BI0a8HCsxaQkC30hlAZhskX0HYLTm
O+9oHSXxFFafM/MWUyk0Sg1dB1wdVsXG6jsGW4gHXZKhuM2Xqd4DwrPhYNn8iLPhu+T6YGF4C2zR
aZTyE7/AOC55Wlxn18uIiPH8ZQezR4vRxUvTPQqPKXBSlkBb0CZCw8A6cElHufval7cIGMYEuQ8t
Xmxm3a5kSoqpT+SLj0WsJgHam7o0yCpCxo3za5HPLJFK5UAR79t80b9DjPrSPczEuijEo6zOJwaB
y0xC5HzylSMjoQe4uk8tuCS7oec1CE2xWIHZIS8v0tfMV7WIwEWiMIPNamp3KfZl865sFgT1uHe3
sdLHgrG3wcI7L9sr5o8f2C/rJmkzS+/sj1SxhqlBgH1UtpvZG22Djy0ERMAzTchf0Dewh26nzbFm
H5cDWPFnYseTQPBDdMo4zi4xOnr7m8Ipe5XAIWo3wtHSPZKDIGqrvC4uU6PozTQa+s5F6STNtP9P
YnxN9FyKk2OQTUM/EpYn0jSwg3a4a5uraEsFJ0j4EPm7rxoIeBABcvCOu5zEKqyw73Ny0T5wYioc
6IeTUsrbNcqsB2pw3jdxTHCjXAadsQyz3iL+ffNl2WgTH4JM6UKrkmmuM4nfoRnLYxnbi1va2gBE
rijXuvonZzAOPV77QreJRIL7c9xJV/ZfuLcT46/R37JMQf7KrGPvpeoi5a+OBVIWWFVjsLg3IH5K
ZbmYGhzAvTF8+MAgdCERe6g53oDUu0Knl88KCP1JFWB3GqKyXRGoTfKs1KiXz4L9w/QPz5UmYtfc
CJ2oHtaynqY4t3KN2l/qHDoiuSY4ONA1zg0vfzgzDk2i5KotN/dkvopFcjNk9jf5iJOtxNj8OS1D
TWGws+CophiU78mxWO2CGeyeT/kxgNXDKWtb/JRUefrpUyIhcACSfF3RrWnzwNQIP5ro5/3tL8dB
SK1kuOOhEyiq1euTRCTLysbGs2mS8A/AShLnf4xLbveTHgGohBv+Wk4NqXJPjvILa4z5oc3frMVz
Daoewtq3I95BjNoolLLCvRqMEKYVT5dCCmq8OfoX+vRr9+9vNPhr2vCmQscRKsqNTUatWY+q40eJ
TAxgLMbWLmCMP/H5mxQdYUTTbcMwXvzLoWOio2BwC5WJkB8MBFQUfRnhNKjy6UsqJD17Ujg+8jMF
mxQunmD18nC4V8h5PgXs7mS8Au5ntYffq3cxoSb5rZJgjQT2np296kgY/0Zy4iqvEaKUXWZXjRTr
4BPIfzgLPEetcePs3aX2p2J4k8uBo22OcUgMkNkKvz7M2RPxPc20bVOaLO86FC4snrPtWWflZEZh
debJfm7d8lqCd9D+vBu3ueOTkcQT7WiAt2628xokEOFnJWsl7xdXWAa+vooEX3Ydd/Cb9N0voFgO
H3/1OYHZLW6dyUVIliVTxGrPZ0/bdW0xyF2V15zUaBMTsEYyRM0/n0L6fUZMEQOHCg00q7px/eAf
UfIF03pkQ87JggA3dlwKos+Hbk8T2dnOrs62nShnUP1pVZrMiUDuWfD/Oi5bO6UYkUxyCNcGuRug
pGYyuc8mgzIVkxiHDd7x20er9FG8OmED+3xhBlL9M5D+XE2b4vm4Odu1IxiuLHIL++uwpGWQ3Jg8
oGHN18RP6XeEG7DJwWrwNl0FuZzknZCTQEEVT2ha4bQuLd77ZuAUjh78mOdsfZ5m+ytN/wVAvPG/
Da5l96zs+gahxZrBrFoCw6kppm/WTORLoeidMsCgtoii9iemGqYLhZj5QsWBV/P7KfNzTdl6d/lO
fRIYgnaQpwc5Xjvgr/qbYCEtRW6f5NwqHoWO6At3kt9C5HNIXotxeTj5RUm7F1xJpCpF3md0cVdX
Y1Zf+w3lvyEUAOBrMCbHXUMMA0WcCc5KEV8miRs2/0h8bTuYIx8xrYzOgtluChNgnnmqGvVb0uti
T5eRC0hXuuZyeKuk+nM8NEmNvvPrErlUP3wwme5mW/cE4e2LIQyOZuD1j2ug87nmpZQN+ejebLsE
Lcg8llhBeDBwkeGdPzfCjFAhK/9N1QHQEqUWvrGacrEoLDZJMexCS2WmBdflBHJx+2ldn8JzMumF
ewgiOVSqUbJh6C9xXM1iDlWWfyZKslxdH1Z1ZAuZject/8dLEbSlRaekmGSLklEIvWMA6MwDz+D4
+v39at+t0Vl+6bo+Sd5U8l/bzLSMiC3Tq0jpqRkRw8tdnctbzAlhiMwHhwWm46QS/2lMthAXDjEV
OyUE1ibER73Pshl31TK5ou20K+w6L6qb6j+AWS2xctvCfXCIXHSlW1zAu1JPEMO6W6cncv60sQy7
gbW94Z289xo6OqqF4JhyEQIo1el8kVnxwn6x8Y3qOzyYQXiZtKdPLG1AVwGBLYUWQG7SMgn/O/Vr
6UU9UC27n5eabBXsj0csghQRiv86zrcEZrqTzWBgvhsDEODa5LJfTyh19n7YyK0id/rN+qRLDhld
0m23xd5FGX+8IeFzZfmTDwKTiEsde5gSp3PScMkXWtSMw7MUbV+Pa9E77/n9My9XUiZYwZcWbwLZ
TWZKvx4oCWAFU6LzBehIhkrQn7x6kesaHT8QGNmBDDgOIoqS8kSCY2JiTSabuufLkib2ccOHVRDt
Gxttw5ollTyH/8DFcEGFKoTScYUaGI/NlewRneQ6AGUNQuipwdZe9Ey3snx0ksVg+Yozfv21bNOt
XSXMtmgJ4SXgUJiLcK/dFQ207ZZTMjyGpUHE0ZzY/z4t8GmHDYSPUWmfzOzxD2Dl0iFbefP7YMM9
eiCwPNsoC5RGliSQCaMqlKlspVUTe5N/iY8wa6DIYYmwSWf5jINEhqUZazPG9ZGGCtQ7pDonzbME
9lhdDzv2WKP271FgtMU0YrItqjtqZ1ZAZCbZHzIiC8vI0kxHi4vc0iscwn1FgLiak19aSNKH5XkR
1T+wIhDDFgjM74zSzzUYU2vSk3nLgo8lwcFLDjEZ+k+TDuYdzK6qZa69zeB/eWAYKqF5fD80lDuB
hWW0WiX4TYX6SNMvqeScDkJ+5T1YmQPlLid7/OWshaUc7RT78p7vunTc37ktjzoT4H+Ik5NgvJpm
NSQIWZjGmhDJ6rRP+qu5K5bxOyqTb3vb2+zB20SZQOKQpAMxse6VG6LEEMQ3z7yezn6JDlqgQ/KP
T2xVI+VEEisvJU5tTORQo972afVXkhLgUpvMU2208oluoYTY6F2emA3eFipiQsArzdKXZ2Fce5dQ
eMoBCy5VodxiUrAVKaxKdRwHSjAZxX6AGEuvvwy/NU2mdBU2OLzvMDAsWyYlHD0yb3rwi7cKGOE8
vfLIMphYKUb5jEpbISFZzLYDKjcLw6swEf2LJE8rNKhEDMtqrcpTVeCMU9+gJsQ8MfNotosACosd
C99yhFm+hQkqMgLDRuCX5HQ41myRdYnYxyR4AqdfzkzBGRoHzd3Z5cIqThiXFgU+emSqu5Ccegln
0S5NIXwOZ7HTasrS1sV5Giz+cT5k2qDZ2VNxVEbhxZbTDQEgQg4vIAzkzGAsTkv4Iu6gGjVVnAMK
AocnDGSf/bwfpq6h8Qa97IYwRd9cRoQE5HP5EjsSHEki892Tw0QwyH88Y3DqfKRlbJfFTSoe65sJ
d8Hu3MARM6KQ569w0neKYX5czebAzyvf50L3bGDukcEcIIrhpc+rpwCphLKJNHvfJklrxXojJCaU
5siLMF3KZ4Lro2cVsXSzip9zEje1LbMHWJY3j7o9l2ZQVmve9OMPhVaRripelVhtfzyoScxPGRbx
xl3Bf1cw250W4lrVtunDCNfxabdb+5KJyHyWTybT83fplOT1KnB/NrQwwoa+RTtc3mrl7iYR3BLl
mZvqoIBLOTBkFjMQiPeet5XuP2qUAlYn49fH0DUU9+ugw6akrqA/wD+bg/YIHVZfHLf6GyBvFthq
LWkBUnZ98z0zBJsYslo9hfXXBEe+A93ZUSWy7nsqV++VWJLzSIhi+8lPQrOmNlbAoksgdg5kwt0Y
01rMh70vPAv0bHrtZZCzJ2dc3z9TSAlfJ+T5ATZHC13uoPtcQ8WrzKUbks4KJuIIFwsqx4pMa3Oe
mYycKvK3iZiZCwKf/XJpFIkj31RkvyjKXJV+5tkknHSHNZ4etf7PYnGPVW0R2ucuB5sRihah1t1b
2KgltmpRfsFzztv/K+AJfHgOxfUuK9HdWNdGTeBrIOVI8gzWA/lJaZNdLzwPf9KSARBe+m9nTU7G
2w+gs8ElvZyyc5wVCLcpqjVzcgh2ntsdhNfH8Gy52UY1AumaztOpr096RQ6yVFJ0hYQi673GSgHf
4Q0b+goGUt/CBdZfpoBVrj+VCgdCLeKUFvRbL2tWn3aDnRdB0bEFXRK5EUOgbBkDYPh1THZb45Dt
hY2TwT8ZURUjOJ3Ux20JJEtJ+lRASZ/8PjKnWk788jix+TdVm7yUrGUAB+DdxKpgmSuHw9I7XN5P
h9x+jLGopDMG0hEdqEzzQtvH130PR1ovmianGS52LkuaETzj3N8gc6xzTWQLZmLhqp+I9w1YAx5M
b7XZtQbJH8nEU4qey/zkZ1WMUFNm1cnSU4mPgJUUkxyQgrfKixuyaO6hkRawd2+UBO5DP9zoLQPF
kTJmFZU7FQK5wETMENItE89u8V9E8xKkPTgXiWj/2PeDaht22/W63Mx2xJlzlSoLwsDk+vuO4Ug9
IhhX/g7MVxbTQ/z8IcfN55Aqy8J1uRuJiXic2Fbw+RPpmr1G/UL2glGAxcUy56fzAUJrSqGGKG+0
9AK4mvOKWZyWGuQ5KKBhDyzPsj/21lRK4aHkuHGDQh+18BX5IVh2TncMCYPKq5SobNfZ1O207hQf
F6pSip4e7GfoxkZmw5x0vfHW77tghngNZHfT+ca8Q9ZxWRKTzoWMtC2gbhtp7rYh1hYDPiWAcXwz
DpCJRlfyAZR7BOraVBiOieBe51VSVkbAvhTS3WEGYA4I7PJ0HEJyDcCvZ3JThz4BHouPwrOSygNH
W41hC27lGjEd1C+6PTsq4GlSO9eW4udXlHJD3B1vhB8iAkyT9zsk7GEq8Ny9395YaZMxpdDMTTf0
blks0wh5RypbR8+BvUtHiWpWA3LbBJmctdyuP9SG74JVRVN+1qqUyZbdjYHR2Z3f9luqRsY6Tol/
10CXYy5GIHttS+5LDgd6g9cK2uCD+gTTkedl0yBfVlNaQnwRoT+3ScvFA5jLp+NnR6Ji+UgAeHVQ
LnBo0PVrKVDGZ5KwoLJ0cIycChGvwXOHdoLSR44OVDHUUNwexb67FcG3eEY1HxLiArXA9GhB379t
DoJFG39z0zUIT3hcUAw6/AmqYF7zjK/xvz404YfWsvXbjrEZ3APX60670gyZn7IT8HYiJIKU5P3r
RK5DvXv213kjM1dYYfM+eE2grMWIdQ24Z3vgEQc7MRmVItNU1G/6gmqDAeVTCQxHIF/RlXo2UE7v
ZPLx+wKk5hE3FKU1HWn5LYZf0UKY7CRUDXfCIfLMgtB7yHZBhSlX9icG/jp8/shmnJANtSodavuM
qqJvIiYCMBftEqxSfSx7JTiqdQ0syeDatLVpzcLLOvgzbs2z0L/zPcEzypZmLQHJhqBiTi2Hlcwa
fBD2e4qWQKRJ+jISnfKmxxv77Ohvz92cY+LVMBp+T9ervKD00r91CyaPLxqbnCNDOY+DUvmCVFPj
zETZzWN64QXAVzt655Sy11qcfc5ai/bu/+fpA65ox/iWGSmZn9etsFxoXOyl9HjXtPekBD8zFnuf
M3aQFtvR4Kfu3cYKSt6QvVWgxsbTHoWrWXb5dHb3/f54ZWpjepWRvExgNkvjQ5L+vFF32hsnEwH6
MT+51WihROWgXsPywcf/gQFSwJ5RPPbIsrfaZOhB27vaVgi6eXAcG75w2ZemY/bKGM7L4CKQMg1r
baf0n2y3D28+vQjk6sryMEW7IdzeJPdEZLZYG+38BK3Gw5uX7tMCoIkKPkDRDQZ6np5mC088ppYJ
yVvZ+2k9lBL80INQ/YJ80zLBuRv1mWPq4XdfeO2daYSFAtL2pyHQBlwQNjxdb0uDS3MtW9/Hbf/C
gO5LAp+83hHfMzSRdZ5LKg9jvezbKoLR0cWEoh7RNF2r2rs0d83/lt5YvBgQcLWDrrHa+QQUwy4Q
CcZm2oagHEn7jLhDbMCalaV+k6dF355Ul/mwCmOfUwfqPgQVZy7pc41qi8LdTEEpFbZ3JN556sP3
vcTekEHgOtdOIeUKclXQwh2TgkuJ/TbOrTwV+uFeQq+WlcCHzvprUydvKL+TvnEJboFjGckyrpQb
f+Agdtm+qgZs8KUUCiR6hqI9L5EDrr/GHFmHagIHX5n+XGV0EpFEgnL2jGM0D70kKvQFp/CM/EVB
kY3tW/Gedubns7oELTsrEjvxPJ64vEjD2IeUCUmK+P3ZxpZ0Q/iMvPnZOMr78e8SG37vaj4auaKx
54D43lzx2jJoFqKh3BywiS70HDn2xtdFO3PkA0tKiUWSshGCaeVmXY5hf5TbN6QbsJUjMuKN8d1o
mbL6uNpo0yRIyIZMMmlyAaCFa2XXH4370GFpdxnznO01SI9L7UyMB/RSePwmp1uNAh9m5zBit1dR
c/nn+ptE+HIxJUkL37gz1x4D9Z6l7pMlNhF2puXps7sUdsVtY9s0bNZHjJyo46uYRoO3ROoomLCe
avcvnfgpJ3uUE4BWwNa3HrsFazi1F0h0h5sczOpwnl3V2QuHc2EH0spaNohty8lbN1fVs9o9rw2g
Ci27flEFJiwR6dvvbVTO+LbzTC4Zib7DZsITk6Btk80HuvSkiXm8AL7052Wq00yRcOWu1ObcNqUr
XnBI0SmU7A3MsLlDyllgsvyQzHK9rbwrv+c55vRhbLWJJaLTbVPjfGuj2RI3aaAMfhN+Fbnk/gdb
pqOim8IJt0fcoifLgJ0+hqTgrobnc/ALeZ7D1pEOQe4+nQCqblJHEQ0fZ3sM+R61tvLKrrxyatia
smrcU42pdlCubkGXX07GDtFoQPjC2Z/OtZ9usaeIWNzmNqqSFtHc99Bb55TGZnuBCUzbEEc1/9f6
vNRyKDgCzh/MIbZRWVhGYy5DrI8uFYPqbn+5cFnXO81T73Zsh1KiWPP/Vtdl5opVJ/rgfr1KXk22
ucYYm3qP4Sz62U7oD/iJETWaffnPxliR/auTsiCWzyvJkc/rgFh/bPguIu+UfRR8oS/uUT+BRyhv
uaZrVvFmOAUif3aRHhnByKmcHLxfp2bHvlcwrvv/cptufDC0hosasU9MGHGJui5B5JRoKYa7W3Wo
+xmWS09cY7pTqXv4Ex4u6ldLONzwmu3c3f6yicsAjOvMiH5RcgyLuAd1uSURU8qflQ2ZA6gXAuDM
gD+qC5q0R/hX8T9beqOboAPztTpfAzA5dIswTho7Mt36gI+pwKJrIEpvQfw1E87ypmNAfUUw51EO
CVhbSL8pSG3huOclrFBxyIjkvcW9uBRruWqDYcHWlDD4EDW98o8fd2/rwIY99OWUwt7ywo0Or9qq
pDSfNWwnA6T+cBXy0Mlw52Ob52oCBrEgXe4t5v0htKaxC54oxucNERuLkLSo7dIduOviRLDsAzjN
3DQ92bnqpyo3lC99aaGUsginHAR4y88v9Qk7w/uklHn183vGk85IVKqu8gwTwoxZxwcOCJLLJwt1
zUuviVRtSVnMifsuDXZJmgYF2PGddWM4h5jFlmSHwiohlnerbvPesHFARvEyAyHqnjhF7Z9Gy6Dt
oD3BOCi+mn0p85iGbyk4rkqR6WUVsAKHaSUiuOq1rfkcy9H2n9HHsRij/aDB0ok7vMCyhDaX3GuC
HuGZRn0RNArFs0WXlfrZnuYZ7zzJn89yYuhoCx/D0WHM9fJk+K3yco9Kz9aXUhQ6/A07Fj38w/hz
KE3m5a3bPfZJP2RVS7TJyAPRtZ/cCzqjZPRey0s0PRCuVGkj9tplHdKo85A+vyJFNrRwRISewYA5
dNHHfRnFaXkEPbAvWwN2d+CayOJCe/LUA6HE2xmWd+uoC1pnS8byuqy5WRzp1QrJDrdQFz4p3OFl
wubr1RhO2ZTNBK/OBGlwFqM406+M8w/obGglBddrpBvVFP4Vc2/MhxLdEjmoxgnjq0JWH7p10cRk
DPqtBpOGr0sRz2Z7G+ykLaWT9v1+wPZ0MIfYKwPGyeDDqIBhCSUdLr1UYGy8fbOlLNtLEB8wxfMq
7gmRCBEvt/aHInAfU4hFkLO9+Oqa4W+bRRinsjUbHUBNnDDDgHr1Z/DhSJpTVsHNnbAzzNbk9WiB
B8O0N/b9ZsTaNSFHhSCkBRYMJLUhmzWlMpqpelXvcO/hH/mvw59lk+UET60NvFk4BvBKEC1bKSOe
55A9oFG3g2a0t2ECNYthzJgtbFYi67hQ4AbT43NQiXBluCj5qtHa6m/Y4PSz3EuqV868NHuz59j9
1jjV1jhlwtiMFBVvj3r0PMAoMPGzPO2bk4QYyPT82ShkEu0g5puVh3fnTeHxDYbD1iIBYWlhTfSQ
JKZ57zB9uEhiELNl8idUjwOlqG9nODG6baG6UYsM3zwV3VRz4lBqVyte0M9YmwQ5gj/S0RtyiSNf
ZSFtyvqgX8aAd8KGgIHYK8Ao8WQukl8qK6pEvl0mUyYX/NaU5IlnlK9RLic1hh0wiQQJ8evN2p0K
kSD3CI5J9Sq9ZFLmC/uWnPAeeK2GaeD+6UQkqnVRRiw88I4dkehu8iYVe4JaMaKDqo/moEPd9yPV
SQzumNfxR8wRsj6+veLdNTgThy0/t1cj/Phr+Js551bEQR8TeFouvptm5UTdVT5aVXOFw1xXvYeX
5PBt/YxCKCgYP7+a1IhiHPdKrh/H/G+qa/2il38G1D+pO5fdx50QOKSdDLgnd9uWcSZ04iD4gwkZ
t57/sPx1p2y3/LvsRy6l2mACrXIjHIcoF/FWBVRupS5ftLRbxKAhgIKSqTIlbUUvBHk/TTCjy0Dq
lDfCiem+hEsbZ58Y5+/DWd/lNN6+WoC5Ct6henrMgT0vMEfzMG9lkgxTH9uiA9hsQRpswNYM8y5/
vbfBmbBTBtIIEuzrMVihN4l/1z/OTMon+OCFEnUmjo1QProXNvEpW9cyuRXdvtEbRiNqGhkj+jtU
tCJR2iCth0j+UDM+vc709URjUaEbUbXahZ97/J/6/qrC2xGoxYhI4cW/NcVFPlxnjmRb9xOdbBeR
D+m0yP2ErdzQwjj+jNFoPGHFyeaPceFmjzeExJBZF4S+GTo8gr4n1FVGVPHu8IV3xDfnbAlIY3m9
UqQCtKFVw76bALLz5xPpYkqGcmCJ9BYUJLKcFC6cY3wdQFs5j9XwdgMob1rdCBlmVjwx4VDK9PWT
A7ihesbOS9JLNeb4k1FiePC4yvZ8qOW0Caz5lAAamjiURxkHf5i1WAO5OLE1kHvoH6CMwYXXYnVa
mCjylL9/Pc3amgE9LDnZJDKqYD3fOT/ncdN9AIIz4NdWyKtIYeTMn1fGKnCRzT3DNXq6edXehCMZ
pwUI5VhcBfNCxfvkL9qt26rAKJx8JakuKyFGBS86+PFUxUmEbN9hrW1XlsZ1Dly5qdgX2Oa3ESNi
vp7ZwFfDiUT3W3wyZVHPCMgCXeFzmV1R4HkCAW/JW0y/blMveEvk2QefeM4lsCyR+Abf3dOCVKT1
/jkDhlakOc+ZWnC6U90p+i0mVqZd6ymd9JgFHm5KK6X+BFXZQ9a27GwVhVj8YDhNuqhfGhN0a1g0
Azx4ZBy5sKuF0H3ObM65q7nQ55Jqxlbn45Zv7wnAHTCHZmgrqaJx72R2Lw4HkD3T2z/D6AtwwIF5
rOl6lJpmbmBJmGeKbrbsn4jOv9S+ooGptbfgJnCnC0M5ae6rz4VZuanHJZ9Nnde3ijcgXUy4JGpf
9n2NJb2R9I8biUUy/ycBL5n6kAhnNHoXpGfHCDbLY9lGBQdcQn4ffVhGOGgs82/UCALOI4Ilw/dZ
YVXSwaKPoqpE0v1LkoDYyfL3yvVkGExCIrlMV046Q50b+pkkf7K75j6wlM+ccVzdCou9kV0L4HIV
xpCndN+K+giZg+G79+rsKg25dItxTZRiJeJ8r+I9DJyUT5NWUygBv5cSpu19N9s+32hz1SiFJ/VY
UNGKwVXamUi+uXX7Wy9ZYux6HCZ932tSJBEA0p3qJvLv2sIEsOV4904WnptM+/VIfpq9BAYfcbhC
FQ1KzXYb/naLMgRmpDEs5zB0v3UyU4oEZutV1/vl10Eqec2Y4nqI1oHp4szZV5riw22ZrdiJbgdn
Ks/dNfXrzWitI6xhwyZyOYZCuIix0H1PAjTzwpSNthv9Tna2bBrNXjCP53hfPUzdjUlZIdAA93Lu
EJbv5aJZDzmdTmOTgFYP0S7Ib34YYCLy4nvbdJA40HXnriU791zSqLfWlCc15oI2STVSb74oLC10
qUMitIhbQJEdIXF4Qx5YiCI7NaKBQhLTrMWkSnzm9hyUbUqPOt+aa/ThbQISfTI4cxYTjLMbXKQH
5sbIl0lVr5dnxA7gcoM7hkqGjU35Rw6rLb4zayuOXpc3nx9gFYzmNKhfasEv8ahU5DPkNGTZbQFA
dHN+zSZD56Dprti4F7rgZYG+snamdg+nLsODCiYVyM98EDAYyhxI/FuaCeZvoaOqllZmzm2O66K2
WOUnwIhddAnQzdJwoqlra1sLbls3pHJpRAkPNogDgdKwkYUjXnXMMmZn+0dTMYngRwxQ5hANeivY
Zs3cdbM0G4mAv9srfF+aIYAKyQ58OLhvRAEhOirsqNsSO/H5YPNpUcnqvNIo04tgocpWlzQaFfaY
zyxsnA9mFd3irDWgt13rgiagPxhUknq7k189erQLwLmtM4AnDwg3Rt9mgnkIhxu0NYO4Z80GvbLm
nELfDzCodXsT1FvozD03o9Y/0vEjF9kPG4xzKymBglSZpJjaxN92wIVHS9gwKRk6MhUtAbujrI7r
PDeo/Sm4/vXKokKJ437DvDUQBMPtFdDahol0Egf0N/LKjynK8w11FpiW9c+m6cvFf8f+OSb6zjxi
jXbK3B/jabRmaXEubKNtj394uRT8G/fmM2OSo1lYD+6tl08sTKNWP9bLYg5E7V5UfKkI8qoxay3f
nM2nmBCCWlR9MHHgmh1ZMXkjGX8QoCkMXqskXnpQVqjngSY4v96Xp+ip8J+fTtwMehM/2RTt/CO6
kXKed8uV6YFcEfJjCz7SdzZfl+9bDpfvggwseN2xItoZjYhRIGR6Deavu2Zx5fomT83Mon2J02rd
SCdyVn5xiKySxZTE90VF28O+r+zxopr305yvbSj4X9Y02a1OjjUWM15sflpQMsf6UJbgm4prvhdi
Jrdv1771f8h8ecxFc9rN+Odfjnwstwn/+2vTWVGN9/E5gaxwQYTQzdm2glUyO6I2DhkW+v5uaG1x
5vXKM3IbhnRndCm6teqz4uszyTziII0OEGlynzMsLz0SieE4v7IvcMsqdv/0C4W1+Afj8b7PAUu2
nWZ6HdN5xNMSDd/yjnXtmUVYeT0nO26tjQwdVDtNEY3S1pjwo/u5VR3EaI6FJe0IU0cSkDTntN4o
+Q7MKNFmhzoH5Ttm0WsNH6ORXHektGvve49rekUkDSCSKiyUl43wwWRnQ20uvFVslZFOOIs5uutK
ClCizRkonHMnZylTgK5KLUlN2MYBP0A4cU4zlgJF7R/rVC4CovrIZxyUc6p9B3f2f8uJ3VaRkKDU
I9UFVeBHLTnDqqG6banAap7DcN52UqpmDRuKyLVJx//HHUKLI2KO5VFMTd3QXNBSpgAuDR6AgF4j
p1Ygn/1+J1a5oihv3tnxrbeTpjwdni0M8DgRIPRBADm+t22c7R50htDMeAqVIJi4o89FVAyNvlAD
Y3HtZKVZeWp8tYd3jiJkio8weJW5hSMr3Pk3q2MNdJ9i7ZXyokos0cqmJCNsv5WOhEkDc4oeaGPi
5Pb4HC9ZtgQY1pkNH9y0CjjCotuXdkN/tnJSYO6L6o8VzdAJqTBwGUCvvSzcGYVEKvRF7/G//BTV
q5nPE4yiIefqh4iKVp96mZ17FuVlbLDHtNg85STgZbnfkdge8hI159HT9LjxHAAwcC9Z9HtgKRO0
MSvV6l4lCsDyheGHPsuh9HnmvWo9F2WA6yVuNUOrkUXYHlXgqwP0yI1khlEB871fH1XIPm+haCEk
QyfGrREQfSh1Y/8vEDjV0JXZamFXZ6z8wSpnziaPLL8Hwmyv0JuexPQVku0SQ8QyspF/JzMFmheb
AYE4djYLNHcHAoRkjmR6R2F3yQ6oYKlxPWeZyjJMslUTIa1JJn7CFE4vIkSVCRLi7jJ5WKZ1HifW
YalctdDvUu5KcnIoPGHvjAutQRKWQhbBguQFxdLWgfh0RqLvYb27LShV5CA7wYXfMs3ye0Gmnt4Z
hPw4TTaWhm9gsIWoGZZ7VfG/2oBx3M31hItwjPLOo/X/2GDDlPmCsBoJR/4VdyZZIOoV2sJFCX3+
tDcHU6mMmS0oeLwtJKyZQVqA4wPu/WlwiJZrd5wVPme6HGk2SdHpP6SQxCwP5qkTbYFaSQK73v+C
tioHEzPE3ObqEZkmgiZS6L7ico3MrzW9gF2JZjVvcVPAE+gxj+s324nX0eJ2OtXl3fqyHbf8gbbB
OdO7gCV794MVkcptz/NVxuAwxzKsV19rdGrTCoJ89I+m8jWrzN725qWtJCmczMMMoVPEVh5/e2ST
513jedzMBQtNhh637s/zCI8xDkAUb3Qyz+iDSiCuviYowxky8N7ANP+w/dodj19FUYR9agPnVoA9
zVQlOQm/NnKrCzkyxSFogQC6Y6owZ4pxCU22tZV/ABA0aLgqGB02V70Hgm6EnvjACbgJt5NQpa1e
6Rg+657s/tUpH9BXiDfRiJCJytBWLs5VnUlJV8biMKcsopRnvW+4P+kduRkeRdWkZ84eSMOGjypX
huhcJ2oCNV8zcncXbOqSS31jlipTY9Ar/nRb87OS/H5ozktXdZ7pxmisWqpF5gjS1dQmlDzpsnTo
7pJ3/RQatILi2WmbiCK6VXzL0zRTVPTH+v3xG8B/eDCXsyZ5VfWfzbkjylv5DNnRmLQPlFgMr3Ay
//jRTv8JoI2nPkjfrGCFa/mG1Wj41xhOOhKCpUmmKN6gpekI6sItOPV0hYky2zviCgkMNLHjIa4B
ZD8p5Tp8DW/AHGw0mVFpnw9ITGftcGTjNbRHUWrSu9pQvqP8UV+6UPziyBdtX0nW1N6n/S9J9MZW
+nrxLorBtf9tC+4KcCQ6dy3Pc5EYBstoOc4OgG7/8HlMlLx/v1cPIoIkOQirEUHmnMWlUmdidn6B
e8+M6xkEh7lGbgVOv1fxQIxUGfBP6E85uvFltbqTrgVbB3/N7boEVUss3K35kObegKaOZbWPkWjY
zfuyhN7n20ZewpK6yVRELuLA65Y6ZZgiYzwaT+uhGBQo+lT2KnPdiX4ZYOUGyl84szqyHO8TW485
Z94cYtYtWv2K6I/e/goRhcwvl7Ox3KNbnmulLlKaW1IY8zz2QrZxMAAj9ssOMFcE3wVuuvQyWGcK
ijJRZujowzEgScbi/ZVB02juldL6Ic7hp5HR86aSlsAIjEla69CoOh0E7/Hk5tJQh8WIFT0+RxUR
bJxlHv+AkPpaE0C5kqd4TQpGHsnMM0Y4AdhiVYiSbfHKKtvH/MDbbQzgmYUpcV3AsIRjt9tQvrUj
sWGnUB5jBVsAjZmQtn6xy9cZ+QQhFkvKkl9neS7xtYEXdg6jpc7V8B461OplzgQAi8qsdJYyfjKe
7hvlVwfRZrDLakb3x2UmIR0L7GQB0yj2of/5im/GuX+yNDcMr1Ttu0r40Wmg6GppgihxTHDig263
nukPSoJuWdVBf0OhDqY3prcmxWVbeOctczSRX2O9nEmLU8LBp1JoD2JlDeiCnI/DlCd3XgHF4xmU
TrRRlIv9FhhDMI9RE4BE/BsvHA90uuXpx759EnLSLYg6IjxjM2X7sTm/XegAGdl/1fPmik3n+JH4
nuQQAUNir/997LNoNhyYWtuZ53XN/bP1gzrxJL2P2b8SRjkcN4MyskBgP53OanY+hZa62YcHkPBZ
7wSQm5fWqLIKJC+ByjOKaeKtArEE2J8anEPvjSHSjkSW7xp3lOSjFIONSpVVeItx2MnCAU/ULORg
0cZAFfSQzWcP1N+lKaXmcXDo/tlkzNphwPEKTmy1gdJvTk5ixHDfUF2GsIco4aSW1wTtkShHmfs1
RfoyWDgJvWOT/iWxT5NP/U0KWlFq0dHIv48Onv19Hvc/p0lNNl2CBpKmImNLQVd0AgmZ6HHa53ud
HUA40heqFt5nlxkPOO89b1zbMp1Lb9XVwfluHoH04OEjjO/ibeHoce1Sn7RAYLY+CMY2jni5e66o
QMbQAOnkhoOQ/YAFPBGrrTY5r7R4gVwbLnI/drW2ZhgIuUzg6oJwPad+gb3NkVi35xBS0Ha3tQ7T
CCltFWXAM8RChmjG7Ix6V8UwrBM+KkIV3JiFzT3GPz51Y4YThZseTAuZtQTQOHaZidytqtulhd6n
hVHgN8z5ucTUW+wBS8E6XEksj3Z3tky68bYktNr8QFG+l6kHqW1TjZSsWPJFmcsMmq0ROH8rJzC1
qIx/3xY+CQ+FiyMgpn+vm1TmvfI1NfA6Wl/7f5jt5amhKnZyAR1NGGI43XCVcOEmXOzlFeHmkDaa
JbBCrY+EtH90F1OzMQQsNPONMRdAeofju70wweaQ5xRHbz3Mahvvn8PZfbcWEoAEv7gJ4XFWj+gY
Tuu/6uMDW28LNU5KatBEqJWcSjncoEOoEDFPnasDkI5VObaJEp38GVssmz7ejEFFUbphBje0w28r
qQFYmU/PBx6v14zpgEyqhwS6b5rkIW6WMNuvzTobhcNlI01e0l8wXNzvEGYrIUBRNn1+uvqQquZi
przGFxT9nZTwy4Tsc2IqRvOKsLyDZExjEZJ0mdi3EozFuvZ/sebSUVSrKqdgriTCguNywnD3KG2e
zDZ6OrdRgKVlbuvh1Nl3tHlx3AUotJDKF5jeYRSKHfBMV5HuH6h/iVijIhEUTyzEPgHN9Stbu7jf
c6uVemjGX87s1T3eXxcYmmUkhh/lUUPATeeqS1ImTTy4loi6XkeJF4cBDAqsfTvwsZI72xH7RXqM
D1zfbcXrHzR8917zH4qgcUfcmOfVCbF1qMcXQO7B1UZhc2Lfz2lFUMH5S6g7KB3XzDtdDqYXgqRL
JIfoM/kA1Q+gdsRbcnMDfcQLKlgP5vSc7Ig2FGHp5f2eqAvNTjMqD+0+HcY9+jAMORnDwHVrXrTE
MQyTQEzw4cnTZvwkPnqjvGNNPMdIC9wEL1mVZch+nn3aqVFQfcKcZnJJBpBdW6u4FXH1tyPCrQVX
BnQh5DIPHfrH3D9vGQRfm0SrdaYrY9titjqz4TWhwIWMHc3ICdCWagG1wwU49shPfemebOuvwa2c
rFSUSX9kkeavnyw19ape5AyUbd0EriUw8bcb7xSStmXCVsHpfN5LjHdrjK9rbHm5uxvkKuI2mcA7
Ixfgk7uGQWYYcN4w25j2r2en7vNrw+Ln/jrqeeytu8zh3x/tcR4peFNBfekR2X6eJmSvwIoNlTRv
eAC51YXH37XAZTFUVAN2aG6kcPaCxdfS1JF5Qfv00OjXHSW2e3QczsNksPysTxeV8/nffBb9fBVY
DpAsg3YHSyQbCQXQgBvN6c9n4xt1EmeaAyl1htNWSU0gnxvkvUTbiLXEEC7UoKteJ5Ap5I/5/jmr
nKDtz1FKukIKxj9Eu/Y9611kt5fzvcMwNo9PY5iPjJ1pYu6+tXH7h7SlmMJGfQc9cqE5RuND0FWx
a1Sbh0uUU7nGNJUYWFjStaHaRykKZxktFC7t4mKqb6FDdjerkcHnBXoNdQKYnSGCFKiEdWnF6hZ0
PFTl32gGjTQCNLDiLiK1Z+vCCCjMAtcqoply+ZcSxIVi6gcLTJu7jYx6TplTR6oNVaFNStnnSr8d
HrPAlDE44GICkKAwwwWfWaKdtjstXsDZ0gAHh38XGg+lrdcQUGA8hW97Iy3WUHzNTAHxyc0/oPh2
1qiPsI10IWVnGwhrwvy5lJnolNML+lvmYvujJjEDmvXyqfPdmKpumEBul7gaN50MKvd8iYgJIZKh
QbjIqJQjK5PgAO/k1yW3Fs6eShCYJSWo7/Sdji3NBzlAwnOqjUHSxv0zX7qRo64MInfA0kk36Yt6
9a0VHe2t/eXP19FDuYXHuC6gOkkvUpgBy0KVGfUtP/P2c33KnBx4djg2rz+4m6AU7ePkw2S62n0Q
iR/03DvuE8/3dkE20Fpjc2GSpDP+xe/6fFcXY7BhaQViZd1H3GQCOOB7UbE+a4OV7zQiO+22+0iR
v5vVlN3rEAgjmwKiTj6vhUhDwcvnHQHjcYPtxe4gOQFCix77PxZghebH0m1BO8u6RUpz+Oy0TC1b
Y5rDa4Frry3qBA823tIX5VFypZeIUVKeh78nByUHc82oaFXc3URifWmpwwXUM+GiT3yD2ryd4UNP
EAZXf5KI1/8aku5vlPf7N35TaFhJmjgr0gIBwZm+GSuci21LBd8khl1AgBLk0YuLEMcj8uXq3kxU
8nXZuZhxYH1QOEXaMFFJ8x8Y+Ib22PgXYyjUeWQE5TDW1oZrXbt9/eg/btrXIgLG0cSrm1PZRbu+
hYu5fxGY+pWWYZiUh7/BqQHJ3zD7BLwYdG2B1drsrUIZcSPl0+hWSLybWmyupoFlFEHaNdlZIkTh
VYFK002icAbQli7R1MOn+pyVtRIEQDWEWyP3jEIWCLpQDpb2nbfBTEhbt+tGkCfs6pQb3HW5KtFj
qA8fdJlsfycapoGYd4CrBWaVhBtQgYm6Ib8BSWJsJIChfu7SJNnFJhhCIRqqLY2/E+YqbyyhTpNv
AdKAmltqefgZ/I1XO1AU1I9/Iih6r1YhpqzNqypJf1Uj7N7PxDc6YaLEE6IlVFt/tJIMD86FWxd6
wRUye7T9SnSwb4ay4rtevGKt7oZ2nLKOKwAUQVsjmoUgZ1gFiFIvzMwDPzwoyMIvundBGCiHIRMp
ECmUwK1WFKiaEC74LCYnAnds5/JsDh/O1TGtfDlf4vtGeHt2L3Cg0zGiVfrmu5HDIcUrhc0D+1Ek
7usAFo/yWVi7eGf1mFA7CmeDWsSdbQvptoN7Z/OfrKZT1t2axYczVmEGwD8TDMYdohiBkeaSQzuF
ZOKcBFVehzGoqzPsGqIKzVX73QNVHx58VIaJaFcNsjI5ju4mSVt3rpJJY/JLsCRPyWotK8ChFJz8
RmMcZMT8wrEscy0F5lJkv4YNWLi6Ve/8DLdWxOP7fKWrEPte9Iqp20+POvjsq/CrHXVNdgfyW97c
PunWXHCvCILIGO3IYzL5I1mYfKJdR5DA8BxdHa92tFbeyEySnmnAAY1ZK3r7sjnTedx/+TcjduoA
M+3FTt8Lsfu6At1LbPU5rNO0AJNYohDxXcaFoPhyMHztX5jKtfN1PHNcyqLEocWwFrurBrmpXN86
lzMRGKjJHY/EUQoghs0bzmlLgkvGlK5uS5Kw3vtW+uJufHDGYVA6hoU/YW3LQtwuvSwNBWzqz8kQ
WHzKq8rVORwlKn8RVGY0KO4E+NKHGCC1pgL1n02a/8PjdkOoc9xKj9os88thriFy1om0ch2CB4K5
VNw3gOC/VST51M/SobmC7nHk7yEY68XJ/ewku66oWQLczISLOw5jQAW26jURu2+zIB5m0g9z0Tuj
0jWB4o3gPnqfioKRnvq36hFi7t7ntXqApmegBkx+Q91xQTbQUG862RM83mnx1frwR7qc/r/dJlyP
lrzpxjeh4ffVlsTklNTaih6ZxXDpKSYzlQTMS+GZKumvgWNF4kT8363Y5avNcJhblrA0DSI/AlXE
yG/aqNsr7p+VBA8EzDZA7iI0RjiImgY7Jyx8uxvngKQtoHgujIfSzJ22lsL+3vEzjRYQGhk5O2ea
OQ3G/aL8ZKRsukLHNcMVC2BHxvL1jZlvu90/0cHkv1OtujK7ojuEV8smrfpCLV3IwSeliCiZ+6tp
BuvTw9Besymh/4BaXObpggD7v6ggiAsQ64rcioSq3WK0dn4sqanxTHQ3q/yo+EF8+V2qgs7pomLp
LUM6tLrLilMChAdcctbBOAVJ7ujQAMaAJ01Ytjg4W0o3y8K7y0NnV2odnzyX/xUYeQs+m7yHHdan
U67O0EtQYYD8Oil+jQXLGiT36C3Tymf3G58ea51yOYI31QUNP0BWMqRx7cGrevRh3h82t6telppv
MU0RRtzonI5exBOLbGQ5+uS3mkFAQmgNE+BBjCxo5SZpMIGTyjEDdr6r/+1LRY403fhkJjX6zncQ
ynMhRQ9tZzrzYp7pK0hODaL8Qoo/WFeIiI6MatOH+pFyiqyE9An2IN6N6VA+Xw/xIFLSeK+dPyFI
+pXWY6M0D66C/qhxr38QFKogZnsEFW5O2a8uqhXFwJ89dgkdV1vPhtXKakVRLVeqox7bcOotAm3n
m0R+U5irnldz56WtoJYiuPw4b+/5Z/voKlHSqJLsSDnaeR8Ro1UJxHxzLNoxAwxHXzOb3JK8WNzJ
ltdrX7FrbpfaordGP0tS7pSXres0D5HoggZBoLxboz2cenPUuj80xsOY6/4zSmhTgbCCGW6QwtT1
6DJYXjqC8fi/0+8stjAwvmrkEFj/hgH1vItLL6s5uztSXWp8mKLvswn9p6+qqsvA5GofdpPNiQNB
VgEyeqdW9ydLUKu8KQaLGjTsxD1vyNzfw0FY+dYh0bp2XAXa6/ydL2f/iPjSNUmmchwAxABeX1xi
bxUadLR3MzBsz/e0IXugPYDPrS6B/GSfM4FrxIA78asJHGodVcRtcVdTs9jSqcM0m0X7OMCFGDyh
qgp2f98hCv8rBX7VnySUwECDN/QANf0n892i1XtcyEw7SOpGVIPzzGvAysu0WH+wCLCZSwNKH3Ff
GQQ9cZm4SKruej77kyvpIaFn0Wc4QXeI0fA/ACcoacdROEKfDS1gJt0R1U3ClQBzJLCXO7rshbk6
NsfUErizwjkLFfTYKb35ck/huopffksxR/AEQrIyu333WUBxzxMHWREplGghgnLQJtEzD3gItn08
mgATzneD12g1umpbSpKN5aTAeT4D4lKE1PsO5nJdcBMok5gRoesZLUbNua5lCjaxcGZEzceBBptL
8nvl5Ie8CZffgZRql6SJp7xk+m2s+EogfbcQIFb4oLEpCJZDizYZ8GVQWJm5jRJA+mFZ/B1BmO//
6yacVidc4q6EwfFwnBNfJKxQIzfrAhjDuDgbea/eHzqCKLHsAmHPBnTWax1SVkzjcbHGcyEAHGVk
xuTJxoFumlIlvbyUA+xT1mY0DDCjiBcbJJ/PRI6SlSLe1nCJHav6lKcFVCyV35AvdemahXLQsvHV
xrkUmlDF0cahjqN7nGUJ+HS0wvjzPg5KE7Inpshq016JlD7mPt0yNub/DF2KwKpg6nHEiu9Sr6He
YPqy6iF8owaYmS928FhoQKkAizPY+hRS0ejvNhIWhDddv58RcMMOQIo1mcYm2jfcNZR83xQa1AIi
tm49CA6tu7WkXiw2o49MxEyPMRyCBMNAY6bwT/pr8Gpcbh8fKpvrI6OKPtMuRFFQ67wXtkcqP61g
srvffLvMS/eiifoCyNeVHPUIDTftMGW0uAq/HbayLL4f4BSAT8LJaV08Hcj1i3CSzwV+7mcH0qxM
lgwg30Dyv0Y8q4DUU0Y/OdYvICwZxrHTKg5FEP8F5HdINzNzLOMtZmNmBFZkR4JU6j6JDr0jnluA
/g4gq2roEUh/HeOjdOUPZncQx34ss6+eMIEvhn4T/UZTukK/r+gDUSb7C5gFxSCknrHI8iSp+XMm
0A68YaKixbJxHUSzzfKEMjG8LhQ3kCcBqdwLTIbmFK+03KlnKcWIRUMmos7DjU+1WnEEZxnHOZBn
+odz46VhCqjrhg9Lp7N/pW333wbaBwv4sUOpAvzEA1EOCqkDPdIz5MHw1KGRyT3WJkMLX+aS4uef
5dvf+y23nXM8upoBDBrWjPV4+nvE/8qMNbfH88UuaT15Q2yB9DQEBUjEswhIDpbZUnA/H7WLhCPr
oHJSex+Q7zExZm1IfAhcuQUFGy9QuFq04M4Fq0LTr9bGthIgAC/b3SwIM95jYSz4EUnO+2lWp+Xk
5rjmA4V/IC1f9zpLv+qtlP1nkYWywCZMToJ+3zffged7/nZd161MCVUcpIoKWDaTaJVq4RFVKN4H
46qg6NjPOm+XUKhYqvA7XXmqpDB3E86ir3UwmjhuvInhlj4RrPde1QWZzlSR0WemgJylLf3t9M6l
b4CiELLYaTfeh4/wzQQySVYwrZrXuW94+xpXnNQg2ssQ4biUQKRwHRxVFaDSv6JXhFtZBeQvcKJn
U+TquVskRlCCnUABTyQZW6fW2KLl/5me24ce2gNOM18kdgJIhp8U9/rqQM1TpQaGKSQXUtjkL4Yw
1c380oAubR99hcDEZ3rCTvKuL8JIqG7fueAcOPoKwH/qCimbJS82EexfpxZpq4vbEEEFt/5Ad+y0
Pu/pUWLtVJmRoSoPdhNIhQ4DLVEZlNu1t/sqySN0C0RtYzZkdsgO/Fa+5ZoL6ay+mM1GEnU+nhcJ
pSuMI1UT8qTifSalXjSGENCgpYPbixdYiQaye3Vgav8BdSn92w9aY/nT0SNmUQrayG1wso1xSUYs
f1zL5dZvISkuu1/O27F8OsFb49F1DssWCg5COyG5ykfPoBkCCEGWpvDRf0MnqvNtjcmPYY9qqlp6
tWnKGmDxFPFx/cDSmcyIHaCcseIhpHU79iXVfBiIfy92BFAso2Y1+NDTNZPc60/NgMOkNJ35PtZ4
kevMD9Ft7ufZaA9iD3ZcZvtUIxNcO5NbkeEyaI+KPlzmqCCAjeq2n0Je2rdCyAPCP08MhbBpD22o
Sqzm2msFVVOHS0kltmlk027w1+ZHpECst2sLDIDYWE9Sg7++AOclpB626WaIBKg1zM7wt38ofxcL
mvmOANDFjSNeH2qqc3rTkY5m6hTZIbNK9FEhaWtjns2aI9KU+Le67rxnJpt70qHP4SYJ7I2UrP4y
U4Y31ZyjP09uB7hIVXFQ//3/jtah7O1lrgT7CQ8sl1yg9Tz+CehV3ydq6Yfh3KYJ/cgycax17sVp
aExFWA23LFX5ad/G/05Ae48nEUVtudBbXywPZyNJXDXTZ3qGvZ2oiC0/5J/EvXYbUbAW0vw6UxjF
E7apGgSei3BH3/R0MZOKZee1T4QJ4tVNIsFxtW5rLTob7G0O55C6Nhlvzk2lpQrTROhqGTGu1e6g
1PCeB/L4mOW9G263zy7GqmBfqCmOnLgsBf2vqtyTlwxNFqipCHfaoa9grgNkKJE57Ml3NLEok+Lq
F+WRex4H65Pi1iN7DnPlL4SiLd2ha6FkF2c5bSUvOOEDSUL4mT91w7sMSVptJDjXlPUJtKNnNo2i
SlrXUo6G43VMxTfT3D8XsbGk6iWqo9nXKuvIPfOXPCzo6bL7uAnwXUiDrtkZ/fjZe4s5LGJB2TpE
GrfZj/Ki4dxV5vsOXF4TXN4oHMEA1uGWQWfKzI6nqJtO3EUnXSpOUWH7PYtw9qnLe+U0f6LzE2aE
vwtQFyiHmYmAUez3x0oW1zGIJhFnizQV0Ckx7EsrG6uXfVJhd2Ju2yd54Zi0/obAFgReeCyWyGVI
HkTjRrOtxepBsycfjmWnW9oDe4oKjPKVrUxTbUJo4MtHeLNRVHA24SZ7lo3ywpNDgBci7Z1oXUIc
wXORvnQxN+4gsUjHh44uiClePmaC89l+AqwAP0yDCLTpiQKFmQmcK80reSMRRgHvTm2UgMGQphnI
zqi+8J59Urv7IFfhMz8ZGOIxBao/AN6rOiSDVpITxSgVs5K7lRPRfGl75QgT0G731ovNd1MEoyh0
0a8/zemJvhKwNGRxt9Ap94VoPqmTIW1KpYsCQKw5zDNdDgalvjaKR1CRLSosSm5dFayS2cEjsO9c
dso+rSI2eINt1ZuxqQjjER6jQoYTAQF45wWUXPzFDYTL8Dq6+EsRr3LL0sEM04xL/5PrIg8apetf
KqbH/SNAlrJRQYyBOL9x0iQQEmQgiSJTK3rFKfH7dL6E2YeGIrYB6yiF0PUfeYR2n441T9TnF3mE
zkvbYzoCpsNaTwLH6SplrKR/gnsu0sjtn5tn+1X7ydboADu3Lbfx2cCimy2oh7MTeHXL6bl6GEQg
D4YVWRGx07YrDHT0OfcKXlZ0e19QDEOCjkoprA9oPMXO0cNLVvcXsdaLrjfhwjPXCQLryGg6NCB4
O7R/bmiRg+bn+xD6hnCmiaac5iahd00VnLtPA38LhPRSeGGhHAehemiUckpvybJKtLge1d3yakSZ
WWAzqaGhJMmB6VL0TjwQSKCcA35c4LScMRUvcXdjuziZCchPRw3CJANx+JNTOMTvL8U7X9Ek0Njm
/aCwgcSMM3EtFIoD0KVaolOqEoZXf0KP+O4vwtSSPPeCjN8uaUTO3IUEkLIeNprjnGnNxZbgCRXS
xALKxwJhvRxQakIPKt/Vee5+O4Hp7bPYbrtN5AGH3TzJrr5EC8euETL3OvObGrXN8T1eABrLt0TQ
o3eJPaBXnWi9VCkOc2qt3Fc8GVSXPq3XtP8eYJccNdFZCE0fzpYi8bok+WtEvRzNB4mS4UmVwxYG
BUp49ptXWgq4lMwlwsu77WRyHAur1kCvjFvR74SGr9N6d53a5Bh4gAdtow+xAWRtBvxwNLDOC/nb
uwtw1mgTZPLycO1/6Vg/QKr8Bmdpu99QWn7GuwLMKGcG4w6XL1yftXoROIEavLgjLvQE0GnSP2oi
HQ3vpbVFG4zAsqrCaNynrZ+6uyguvXJk9HGGcV4v80DzBYLm6w4DpdREYepiOOrP+16iLBsb+FR2
rV23EMgWgezESN+b/EZsrngZtHfGlOCl/WL6FUujOcN+uGoDZ7e8tuANSSMquvwgl35C9bOiHSiC
HqlqVoqrB0IJ5jqEcVSSqoXn/ZPZFSXWSfJHUXEGsfdk13al3leELngX6fRVMmzHT6+emn1zeChr
ZqBTbPiLaPUca2KoL+OJDFwnbIscjd35gtdwnslXMdH0BcJCThaL3qWtX9cuINodxJPLqt94XyGb
3oJu9q6ametY91eBHF9VW3TcaeV5q1mWTYb5N/ncy5iyRtZKyCfx/0b9eYA53btOz3ilVwyj8TFg
DIJ74KRkZ5DtMT9x1bYFZ4HMU8lcb5jcTtgJT5HSptmdA11RqQFMAbCFuc8zs4eZfudfxegCyWWb
ZUlPPb2Ka2cb2vRge0zWszV15yDgz4gW7rkSN5XEqM3vPBeaXvL/iXYEGNawUEJqTyVCSrXv3VnI
AvjEh0NxMwvpTZ6fmX8R9EB0aEyyFrmoCBUEzKl1iRcMxFDHHoHV3B8+y2vawNRitRejkqJgEzqD
ePnVTreWVbOpS76f0OAXoImkD/krqJ9W+l9jElEQjmiIwcqMWV+0iGahjpu3gl3iXIAjLJXUApSu
4bTaTpvmVUdDcZchQfKiL1mcNbznCe8FzPRvKgLmeD+2vQSI6l9BIf/LIF4jF1S5YZvvXmgrCAJv
bMS63939a4UqqNpQaU9NMShc5dXrHab0ZDmzdhJsYxVhHsUUfIdtfqz1eYDhJ2IxqHo1wlJGTgbx
r5aG/uQVePNedTJSjZi9tphODMggY9UzyWVEjuLvccXimKE53jH+JT2VD2vwxuaOgS7cEa4SjgHA
PWRPwJJq/YujHuoCiJzjVObMiCfNFq2UOovDGpJ+5NenQ7ndKa3lGfxSobo4GNfQjkjiAxA3z2N5
4BICZbgFuacGFNuQO8j+iGLFrGr10V8p5/8WUBbFNLiosOxZnZFXEbIma6mtSRpBwTvKjPGvHicS
hVQ+wvJ+RiwVKE1d+MDHSMcMPT6eVb8TFYoZm2mGQ6y1ccWRp+E/9KkKyjoQLjd3cWSfXrf4v+zS
m41RlsUgmpxLLIHQiQCeyeEkKevSOfHBEDOfbUKS+Y9Q5qQ0xKFkJTiK0isadG00bI0fAjpXfLst
BIBbZOeSgZgZUq/3IjJ62O58M7RFHhEMQQZgEzE0L5xgkBswUiRoEJezT6ly3m/j867TFoOgqt9E
upo9O8/nOdl1SE8qKkkDG/HXwX8cmwenPga/00BN/6H83oVnb29tPwro4k6ayzRsjmOJRymcq3B/
O0nXxIrdc0nRUmqSGnu5MMWcNxnL+kSaWqao5+nq8ei1krcCVc1W/r9bmxCS+/s0g0IELLImyI7B
HsB5k3clh5QsFcX4QM88h8V04mIsriDtoszlykkzm41JwkKYwgW9EKbOoF/8pgSSUQH0QSjmFM2H
w1vSaPCJFU3aOKPAuE0u68ZfuPnYyHN8zos6PQkcYIwzE7ccSYoQJfs6fiaC+ivJc73SDFktcyNC
3ec6ieyOKvVnvM3WRSOQZs3nLJf/daRs0BW8XFdQ2d3YzScByBCSYcsypMTVTmMlS8+wiv3uDGwk
+t8xEVdOzkkLxdF0rUVF7UsY85zOo3Qmtnz3BykfKwTZ7Egi2XVZRliCPoz3+PQ9JKG/s/vj2d2P
Hwu9XI3zn6x2hRAxMo+UY2zxRFLSyUZnavBAjOeJrZ1+VufEN0pOiNkzHfWbQHBHEkvQ2JrUlIWb
zB2mW2sWGdG/KsOmt1vzmMYpkVtBzYiOamLMGiTiPsojg23xNvjda/paHL9zgt0j2OZ4wqfLz667
Of9jIydQisRzjsKrJOgKMazqIKagpz7cyX28bywys6zRmojwIbTlD3LB5xpQdafzHRCk8LdZMc7j
EENVpxZgDCN8j53nn+qTlEehJrtWriCyiFFFLVPIAMm2b2JE3oH8ApJjZyxdX0GnbnMquCevqsWO
z0dPcYgDxYrcOjGZr8T4Vzz9q7svZCfP+d4UcnyRQCsRl8rzXvv+zaPpM0Ay3nkpjt17lslwpojU
D1clJouyAPq6eNtbVdT+1h/QnPSHTo1hvT7WtQfgEJSNn3kOVY2YBg5nBCj/Kfahc90S/ooE4J1K
hYlnaTUcEVspS7vkFvymkQ9UCT6bVBG1rxWansSuvyUiwXs7Gz0A+pEH4DTQ7U8YLbFEnGBUyOFH
v7rTMe4L2xOoIWnnDU1mzcQMdeGODjarl5U7lu4VdkjJIJhFOZ9wnbUPSWu/wN9972y5vc8/ZpDr
Efz7bMlxtJrdgCUclEgyhNlsj1NP8P64CrSsB6pOmd/mMB2PJoJmNauLJOX05hWdR94fLSrwfHy+
POvkmiEII/LU+aQYlKciSubcx/6K32J4DFLCk6DkX4zDHrg10vEHl3tBTGEDl84TH95FKqvczZA5
cAaeyWfhCAOl6UO8g0n7DL/9TjbRB6SjbondMY/ZQxP6Vai0z9ekEqQup8Lj0ZBG4WQlDk2Cajvo
JEdw5GGNza6OEBz4OCMU6HTTW+gCdQskEvLv8dN1j06Ychz8wjLAwqN7matuUJFDxsoA7ZkaFYB2
0h72BNirX7JpPOT3nsqP/HwCDotkU91MsRI/51ihi+nfxJXBPeenfkx0YVujIm0QPg1vn3fWNBoC
N3HXhaZbVsPxHJ1JftsHoYGRAGC6q+cIH47s2EC8sQ7+HqjxMaFLLHDEyc7uEd37QSDEQvbYKNbh
f3e47iWE4dHy3dS31cOfTVAA2D679AF3J5C/5RUlHRzjwlHu5CRowud5Gw4n0ffFZ+Wtae3S9IXr
5Kx2JiSEFGbaGh2AW6LQtS4BhNygfVZahTiEmvMhqhsi9ALhXgxs0zYYiDeb+au04aas3zZQegbR
Qi5jdTOLYjtvdqjasF10JOlFkn0pN+Lv31w2qlxe3Vr4liCKcmTgX7pLZVl6SJcQ0mmtndfeZd6e
2W+LqYmMJfhvn3suFlc+OZheEjUfaJado+86z0cxHDgx1Pp8uqA7IwVEocpwxCrjb42Yc6xNB9IR
0wjkuB7HBPLPFTQdxOHkzYQeMPIRBHZ7d9ZxuOy+uMrEWlLUKHnMgStm4BAiW0CJntqehV5vrR9a
hOpiN8cNTGeYLW6OTb7QD1qRp51jummxmhhl63r+BEV2y7ES42XJbhyUUkB4cml75RwloZKjRUMN
ivX+OxfxPVyne5bvg8KT6apKOWmcmR456ltnT/qjFyYhqOHY795Yksvunij9QO0kJLVSYD85bfjA
m3TZP16Ucw4HxS3TW+lt7qe2vAexuG071952cDJ3v6wGVrrary+4P3GzKpyburNVoRHu8pqKmJ7x
hqdGRJPiT/BNoAPgIZ4ReJlFpETc0agZtt6yXdUlh054SR0uRX3aTtZTrBLMx190D2Bgal6D3hUS
fEMloAEXtATi27ezJ1dhgkJMFlB27YgsojjYuXzCII6Rq2NJOI3fEwasdcJimTvkHU5BSpdVctcF
qkMacTlBw3ajv9k1W03DE2GKfYF7AlRyYdZy7b5EsMx+06V2zJlf5T51WCawIRhDH0Z58vwXJVFl
xfkxs0+5xboTU36gYenrFpsYF0xzJN9Jv+vsCXP49+LKSgQLcOXg9Si0JIaWCqmGAfLeBjsonYoo
yVI6Ptd9bWHCXIAoaJ2QMJXuv63u5M2ZMqt21sGpq9B5OoM+qWiZfXZe/LIYLHfPFnGTy8v89Jk2
m1spUFTYsssViBU4EePUao8b0AMv/eEqIpumvD/TspsSVh4YBfZAtyf5uvsB07QKdBbw6RRXDqR7
WOIGh6rU/T7fDyesWOnJuO+gbFa+0e3iXcPWHKiOMp07HQaFSDs0VUXurH90EPkI9i4H86paYqEf
9GJGLITuNUsM0ILqQwa2GZFK1DD7Wl/LrUWsqvGG7O96JdWgqMnDdb7ibJ3Oos6ff7z+BL0ta+7X
lM+1S25QoPc+0iq4H/HAGcFaKEpRGkQrIrnvzEx4c6DNcREUwbxL0IhQcTRrvSONlEhGlBD0EW6S
zAZ8D/ARGMmyjyxFSufcdY8XDV4HAlF/d9GTStT8v1lgZvFtsQb1F31i9i5XZqHLS0R8fbUszS7e
+kuC6dj1wSImDsIrizYOrJCIPKN0B1oIHkxQGU26vZxQosPb7W05U5L2r7TQLE2U71IuJmXVBt4p
WKKEeQucH4T/C4W0vkGd7ne4SBK9+gjLRKMNEG0znb0diTkiPdFTIAOAdEitv6xoDFokeHizgNN8
naRe+CFV457zEtS5veZ3Vj/0L3ZFWzu3kCYTXWBM57A06FBW1hVA9HPA99AQ4I3x9fl6FG5SNW7g
fpJAx5lIBOtKorJBDv3PE9PIA7bW/Mq2zOCqz9PGNoNrV+s1mvTC9s9DIh8mpYgAgGLKQUstc4M6
SSXK3wnNPb1BUBzuA8vaLZYC8JmiB4PNqy4KedoI5E6mf1+k88Xj+kxEMxVP5prO7CF1yxe62m9C
kSktNaNKmrAHkyOupWMbS+F9EX7X6ccGIgMQPmjQgUgULKQgL/HKH/TbW3QNGjA481x5d6fB3ReY
ofbMYToBPqKHPfX53eH4C5X/CHThUmeN3VBzGDUafxRt7be5SmmVYIJdY4lx7vDepeN9dLdg+VqF
bl7IcvxKc5k32t5vszJrdcV7xE4kwQ5HqUbT3x7FAxj0eDF49C0Mj+L8A0Mj4K+qPu2u/yWKoT6T
WPx15X46IgIhEbwwsXbxCmk5krI8jBPEmGC/fAp4Y2WAOoNTxudMQ7kPU6BLpJGsAXNmbxZaXO6h
JyMpUThBB/azqmTw/bqrbWnz+IUErk0AoIGb0XyH3ZIjn0V4u0EfliCAUmj9g6xYa6MiJEPhMuSK
rXjnmBXvtKjEtqYflkPJfJlI5XkxDgqvr248kCqeohfuNhQOd4GDH5x2xVG2pr2NvUOlIcZsT4Wx
NaNHtbIIOclAgL7vAHZC9FK3EcWxUYU7UOhZiLjMqSnlMGrXHuGrUbTobdxl933rN2lPvbw7md3V
T5iYaL3BHqVppnRPRODfTHBOtcfgCSFgGvScT9T3DYY3VSSnfUA2MR8lohzNyaHzEax0ATOF6N6X
ak9UHr46g1Y56nBzXpJ1LvLvW1zaDLpWIk2mc8mkaEp1mvDJ3RHtWsfL6r0s7DksN7xOz/qqxksb
6gI1kRkdJcQ3+dMKM2yPh3xdWjQD/++kyi1hPiDRidV6UfaEVIkxdHKbFpIZbuDmbGYkLGVnt3dN
DaCCOO3LTOBasYLIshwsGrwyrFiGsJx4vFEwyqS4pqTgxlR/MANNT5CTM7QhATrHGpemyTCGoHuU
pYllP8cPydUrIOagj8TzlY3JZxQyBQwXevhEPyhkvIf6NlunuW1lRNQ+FD/NGt5VqoWfJbSZInFK
SsNYaFbQ4fqiN+GQFQ6Edes4kAvURDW+e9x1Zen7mcA89srdhJCZ3GOd+VNAQy7Kgyj7zdPMx+pT
3YtshaW2oavN+2ZLPkYSq8OR/CGKK3CSAUgiU5inWH53Ca+HdLU7akTykpQcj6K5ECRsG8gD+Eo3
22BidPB2GZLU7nBSRt+XwzBvQS/QldH+cE4ajFl4XcI3p0NNlMY+u3x58XN1DGlLCD8lZsX0Q20M
tTooj/U6e5sbT+r817V1VGkInQB6XvT6i5qelbrrxZQ0+sVgdcnbRQq3sVv+Ji8Dc0Zotc4jIpYp
CzR19+Y8CvRHV1GZBFTpqBQX3/SSuHRzoN9SNm7eZAnePiZAtyDc8+VrVlAjFawIGvOGkQSxLdG+
tRlQsHcCLjIwBRBNWvUVZVpSmG/D7LFnYnLdYW4szWBtTQhyfKuvgELz5ieun3aUcG8pGKgiqC2E
mwbfPLSGWokF013BHqlTMxEIDiYEv2ejMzwHzsTOG0/6PpLQiTiuPvn6BpkuOXXKUMhbd2U4x/Q1
rAFOToOXpEh1CQnTnyKiXUwbRG5lMFmpq/NyIh3iZ5/vt69ZhUaGgZk0fKPgcKPyIoXjYE73Jioo
6shI69oQ3iV4y+v1LSP8wyf9FS0Tren2Atc4qSrgo0G34yp9KYlZui6wcn6eFTx6jm/a+P3Enx1g
lpGzg2i32gDpw6wzNknVjtdod8Adws/hXKIj0VgaPx7oIWNDnjJKClbjSDmFWyNrozQ7gtWg5jsz
CVEE9hGqN3AjyZlPj+JWmDZEMRkmjtzSamLxtmxFPkKPTRvlU22wYWswjcUE/dE/zfDc8LjIA3JK
Vmf4R7YTBQ55un3Hh1YdcZEXaQZJ9lIF1JgIbWozGDM05Umkc3P3S+s9qehRZ1l0OGzOoFWkEr14
6XZajnq3APtq2TEccCytgzV4IsrXLe54SLME0tWqYFtmxDP9wyjlGQuuE1jo55MuIB2RTSaZDX4P
XkQ7Qr2HUGwAKdmNDqDe4DuVlFZc31xh/LQWLYTjw4/CpgvvHLO9QCa06auL3jxAtylCusfzGEO5
vF1kEhMtp2+RJxSuPpGkPgXtoMtw8FBjvWA/vQQiTWt2K3qgbSp13pc+0SeLj23zeS14Na9wsEMt
RY0Wk1oTF3InYoDlihs6R0noxWPfQTN4S6cAr1VlsQKbsIcvV6XqH4/P7HWVpO0w1ZItcXG/PdL5
4OLDwQ3bKJiVSvzjMvp7SCjXXIoKMaHl2ujdHsPvJ6Qp4NhGiTEUo+//LNLFA8S93IvFWvfxR5W1
3lgM5nT7VC1vetGVzh5KIXwE6ig3Q3jaCK/e6rfE/+dJoDagaYi5tyqvK6DsGKQuv0lMkcN6PVH+
2Gbp+uBPd0T1C3LTYYUIMC9XXC8/hT15EoLh48UYkGkIOMo+6E3QinAr4dAyoFdesRboAZ59EjGW
c4b9zTN9KsmqDCXZ0ymgYqNHOxsjOG+a+vBgtMgEtgH3S9fMRQW2RIYhD/PgBePF720QHviQDFWV
k/moRU3S7vwKe/CtyvGssuboYEWRhdODXzjxXNXhR+Z+8JCPVTb59/IeidwrFYRT5JwUgdFchTmA
LwhuWw3MoLleAG6mAddVyYpbL90/2S+n0zqEmYyml4kQsS5xof86D3tGvE72mVZswyWSRxtqxNCS
OeHLpQgTK56BpQxQ9ydvR/cPfMTs8FRA3YlpM/AIVQkaFmE9UeQO2ZqF6nBXJDy+hm730uaPW7NT
sfWctzrAPWhSyZESR72N+dwvIPKeGD4v4h9bzkhBuRBwoNi7hx4vAdVK2JkgcpzbXiz5dnspGIz6
my7pVRHzAaRjFRRe0Msx9/4BlularuAAuv2soRDE6t7sVNz8l6BgZ2/6CpQ0cN+66UgKrpzjUHxx
/3tE6fCIKDJkEZ3zklRBPAB0XTnPK4e+SoPcvuV06cDW7vAXTo2omoNTgsH7fflWsjd3QWnD/9el
V4J0gkufG1tGtQ2l/Bl3/5Zw3v2aGapi4YGK9ws0af7lKFNj3F+AmqIWeCc6DRXK1fPrXN1zJahS
bzcS3uaIosEXbuW/o1cjWz5aaGwlZKuS9tzyJOj9aX4oHaiB9XvetiGIz6wfMXNSHbOEVSRtvJV2
KurW+KWITFEBz4rK+cRkWLYlC1MQVgDip13+eHXqII7wRm4YYLWLlAHa7SSm2I83BZoWH0N6iIeC
6OuMSOgxM9B2fkByOksJURIX8NQ2ZE0BMDYI/XcQo+y7xXjjnbcCf2ZecgKJHv4Vkp8u/8alXKun
nyjOH+7VmUe4uvX1MzYc2ikfI/roxeAFtjAgsI7NX2gSSUzh9GWGOkdSqL9SxWaFWpmFNAH13LT3
xQ6withPyOxLdbfycx9Qv4Nu6IK+TSCbeofotBe928yW630t8Ir/h0GbMRhOIFI7JS5JJxCmcV++
rbZh7qNKaFsLRMwC9fYgICqQJBP6SX9ovLpzIh9bCyFJwrpA6LcW8wLuKEAGrxhcjphKxdcDlhSO
jhzSAU6Y9So4x2xkAsVoFlGurtnQbOCDi0d6QIQkS5mc3vFqNrnXJ/nFptg3WowADDG8O0fIddgt
+TNhzPAm2OpQJw2pwjiV+v4Yom4KPCu4rZ+H1c4Zk1gxd6mdaUt148DKED+Z9g/GNDVjJOePJ3Xa
As9g4kNJrSNlFYBpCTSkELsq/nyeI2uZLEE/jA2nPyFYWfJlgoncq2hH3gAw6rSP/TXvDFJn5B8e
vSxAG4kHTBHp1XWSIH+MRjif4r2TvqkzkSkPBESL8I/hKj7wlMiarpLECadpQt11ZZrnBGH9koPL
WlQ7EPCzkpal+MHHQl6HTyUyJSGrahiyDauAfVLsaGYKF1ACLqkfQ7Ap+EoLMccJPwx2scPYQ6ed
vJgyIKZbVLMzl8maZSJoo+nApM8KQ7H13Kh07cKbtvkZnARbxcMO1hVqT9Lahf/lUKZc6eIFTqyT
o2TCHxcMc8Iv+bP7dkdDOa0DEd5w0cb6WL5KLMRubBOX4Pi993Y1b0oLwRTaTYdEfbYk6V8wU0lz
r6ZePqG22Dn95M+UYiSRAeUnOYNKisgSqmbkww5D3eI7UqYnjfKmPvVqmIR1wzyfCxbll9uGpm9n
2MA6hSAOeJFhiFA/BI8ihHQYo2Q3yO0h4z3837FQpEB1qJnBoqRpEgk4lwwG/KYkUVvpLaX/8raD
JsJidCVArjCw8/HgM2SsZKRscYsywsw8MPzw4HJgldeXwB3VlYXI5Uv33NNTHAmJmxD4Wjeo7BdU
b5Yc0CVtNUpg8++EpcV2dDAwm575IvJo0ZFWJPU9U3r8yJfVWBNp0M+lnsDObyKqplBStU5fQock
aYEMd+mqcpmhVYmk+EyU/qotBp38nBPoP/jN9hWaFaHhvPleRcWBCltTCDyFfXbL237Za5cBFl39
daW1CYH5y+G0omDxbZ429mL34u0rSOEih3hFMIE4wtVNZMuUxaCv8Hc5Nnwr1xbyFrDPk+fp9yKW
/SYzZ1AN9iKcMZc5WEj1pPkQbALvZZpomTIILbTD+5k325OHf0xzofHDpmPVfFx5LOm5SzLccNov
X7i/Zz/cr497vV1gL6qLRVbp8Q8MZvKOpleB7m0qlItHzgW+mFUXQ7sekPSIfvJGAFcQSLB44/Lg
0B1EbB8hlJ8jkM7ycb+mhV2P2s8q7tshi0nnhFxitgyrF2oOlpXqGYLWlmRYJerKnPZPjr0gQ+hM
C1Bd61UgNUx6APUFEwwPvH/586pGVzlOSVfVwqRBYecswGnE0B2QWEA8Di+9O5nFFzyhLZjFjUZe
DeaFRwIcPnM8jcCWwsgjJDFaSrG5it+yEzlZLsA8Kq4g1ZUj+l+ucH8SD8GdkdtnP5QynTjpcLwT
/u0HDTYfKf9CbUDYAJ/u0cgcBkuGlbEtG5kT4fMsrspsjeghLL9f9TmO7VtjS1Hhv9I+QDU71q08
0Y0au/7P3jCyp8E6N2sM4SwhrOn1ZoERWZz/rNmmBIDJ9WQ7YPFFJ42I8/fWm+6BF2kufpcCksI1
dWGERcdiu+DEdW4RxxXCAH/2mKQsTRdxCAwMaFKtmWvtZCx/YGVkTu4KhKG5geg5jMPW6OgU4Bpd
yw3iNxG7DIB0jO3tp2dY32EM4nuW76uiaVn1/Qj6MbH1PFLGv8+U796zm3o2Ito5MzLJ3dtUy6r7
aujj18dE+m38y6nhHziTcBV0E9q2wsOjDO823UGttmTlCeQnGmQ+1T4acPn/O6Ovjeeb3uZVnJzq
ThV95tpVwTuah62Ow2cz/5eM1Ow8uTY4mOpQ9Hxqp1GMMEQ2Fg5qQFTonq7IjFZyZziCRk5B6iv6
fRj8oEp3JSjkq/CGwoz+sXXQWk7+m1yTSvaNQ1rLKAw61Yf9Wx7mx76QOx+kEfkCgwvqnCWLdD4m
djjdZK57pdoId4Soy/9i017Epq+idIJGQ2+yeBA4EIyNBIjxH9FeH6VXsueLRdKkL22dyzxUi7Ij
/wKmWuuDEoVfSpwnuREFWq7h1/L2x1m+8JvJCGFo3LYDx9NIZSs8DsayAI2N9opEZE05wYLWRKvN
u8I1IW6O8240beb7nP+rLreqc6dQT6A2Fl3ZUeKu/LtbEVDY/XijSVdBWQT0ZHaFuHhNsjMGpIHp
f6gmfXMkEh3eiBmj/rFLweWvzAI+1RIghvp0j6KY8QNOlQO6L6NzHT4bY51C9nvfZiXcz/288kzA
0NpDLfYgsieRSRqlNhSMzE9nFT9hHUMR8wWwEMpiHCb9Ntcc7m0/2Mb0rQDceTxsZx+wPVG+d+na
lR32l0DAGTKSCbLozI8xPeXYMHHOOkuOPJlhSPsX9pRTa3QnrzXjk94a4pLDkZLrdyb24b8SixkT
tW7wB6+YkSquEEneKaC92fCgarByjJhpHkPkkzU9DsUc19d8K1Nsy+swk8qM0KOlGYQ3gesU+5XF
wM0CvShvkEd6k6X1T5aTbwJPHYD7RnvxEwskPWcftlxYopXmAwaD7hW992nkpuIizc/TVbHYJ4oY
YjFIZ2GciXgucgFENWLiFI8EzBHaXJdhwkWqBT+BjkW4TX+gu4JuUOFccSYrvraW9zmGbtnrgoDw
SWTOrGwbKFK6m6Q4UqKOeivOiynThSyyswDMPKkV4DpJmyLQwvM/U1smpK92ZFZL+gyv91/UDWX0
UqrhVO7aammArSQ3srZyhPcndq9bT92UAx1OibfhNxOOb8N9HQZIpTue2HceUVSZkFUwOZ2vujsT
6xYBDJKGQiq8ePO3i4cvVCV7j52PCc7R77PkXXyEAfHxw0kb8M1qWj7KKVGUevu7Nxu5vW0X7Qsy
WLfr7vDahXENs2BxClnek840s5lUM57E2+ylnRG/fJiXpLho0IBufZSa8TqnK4mU4fpnbMbfMdGL
n3+Do2P7lwhsdniPb5rLLtleoKG35fLRR8jRpW2u1ubphbt4UDIbG2QSpkaMEpUWaydb540fUNDB
hXCYByvAZU2Hhxxgr+glhkPCGDxBgRoU46VNUNKUB8/+Ht56q5VFa1oBwgGiaZCb6D6qR4VpZYM1
eQJUjuA+do0n0E1aJCSZVlwwPTFetQw+ZF0FhT+uXwA3DF29cEwgyeM13rm9wXzYdrV16ewqRLgU
gQin4LBwUkIh9Hjl+zGz0+XuoTaT6JadGWqrx/wHVAtckqGE6MdtQ+JsYPibVsJALK7D+NqwTWFm
rHnn5fjqRiKYu8w126ks0P//msn0Kd5Ls6eYpx7ksI2CiBJi9uELMDLCDG72FtlneWICNl1kX7Cm
YdAOyouY6jegzQyCeFugu0VI+N6+ilb7HTQrPDlhab0uzarjSkmoz7Nrirat3GDFe5R2XnUFDQB+
zKV6+mSOngc3Y0f/YzzwtNwCieKB7jwV9Z/mjlOaTqwdf4xNrQdeJugTmm4kRMmQgnL+3VyEU1ys
6nVjh4isyKTv0/yjAuz7cZColD5PcvaK43PT2TUPQC8EXBckx0XZMq3Rd4sv2QBP3FA5yccbA8Sk
SepFaOKJgGuMfTfh+veFx2J17OnpEo60jZ/T1IQG2rvbwJp+wZ36elZReg1icLgWIr2VnJtysELM
+cJo5fEjkmgL8X5AYzG/xnRf3XOl/cCJIvPfUfpp5jRE3lUgopMXB+CSuhSNjuqRbPxyZnixbEBa
wTYUJJwiwbEz1Opqg8+X0QXIJ6eMeBY8YYLNAQqcvoi5faX1Zhn7qp0LIFRsV9prNtIRPOWvRL32
bzbI7IbvVbJNNEEexz8/mzGAxXS+oNYOLQmLP/uJH99J+L7w4zmuEcUHFsI5mbioQKCB3AaFg4O4
HNVLfd5IkpJmJQ3iCGG0TuMKQ1ZeD309H0TQwR4yloe24UGQ7/u/VeP+wJVQnwdJ3Jyf82h3rsQS
sQE2fTQKtzqELEWI0rW9vc4XQNOI2j5nsMbz10DMjrJ4uZ8qa6SQRRZYXeJ20TO1tbS/QilUfxUB
3uok+W52RLK3ZkL2CSHGynvLbV5R3LBr90f6F7g0aUkEaSkkM3Nk2yC7Q9+zuDFj1xqzR2G477ei
Humc0Wwh5T8OyKYSVXMaTnI9aOqZyDgomAWgin0iIS3znR0SoU5WBBr92fU7agYAMSjHuakFF6a9
ogNxJv9FcPIPIwnzOxjy7HAmI3H9qG4F1Kl56Kk11O4Kr3DCpNhYDtQCa89wT30i5nXoZ3Uxh3sh
+YMvPd2f23pJO57nuQlT2oyT9Z06jerpaxS3HSNljCFUjU7ergJnE8oo+fMI8C+xk91XJ9fQCnWF
6EJdAfhym/ObwleUzSnlYNUjw/aoptSW0FhneVd7CxGCdhH5EAE1AHi9ygz8ffgffYuNrbhLBh+g
JiHBJlDVu7/JpusOgdGpCvAbfwH0va7icswfy0Py0jy1jA4H4GU5AuEkgFfH4puSluvx29yjESw8
KwGgkTNaI2A42BT+MEMpAdmMJ0CMJr3ZaGsA7We/MqiDjAf7NLQFYaz9JFUNW2/gRwQyFh+eyCbG
2y+OyUu3BP9LoFDI4KorD58QgV1yFZWhsTH+n1eNkhIFuqtUcw/p+/6jwJqIXDIiZpm9FoK3mUH4
as2wlntQ/kvOFiEQoias9PKwtPZLWagEXez7J/JOpfyXeRhj2FfK7aIyRxA8GZoDEH0oo0pDPAAo
llyD/n5pWz8ep8Ln4kp4KvqgS5nc9uZckUPZkqJIalTkXR8VsSs0mRX5MhiE/c9ePCmCaeYtOWjX
XtdkWDw3GjQx8MBLq0pxjX4pr1BAz0v0wGiOsMFeXD0Ruosg5auFLsQ1EXmJy2FqiLSs/d1Jt9a9
1mP2wus2T1RhvzyC+gLa+a2qiYbYntzf62mxgV9aZyybrSIETWaaxESgcYOcB23jkqYr2YqYCvAX
BnhmfeA2o4dam5/uwhYWbA+ouS1llEJFQG1EbxPcxbkhtUJdxC5ezc6VdeAtzQjeNLuL7qadveIP
oyNwyCR3XlYzsdTU6zoTDq+7zNVuqSUQJiPCFOm7heJTzBtsC/++h+YuTOUw5sKTWABwQsuWSb4E
zenXOO8aE4szPIzvC7thWAgjc1FmlpeuY17DCEBujdUCR6ccWjMnA+i60WBarx5m+ItAvihjMtbe
ZaYYF6k9z6D0L12KzgsRY4sTF8n9LRxs8n65OKKhvFPEp/lC15NR70XXvaBcQ7Z/348hDvqtL2I/
FY3dE3wk1wGvruQxfVxLklPNFlgdIXs2RizgZY3QW499oNmfxndlZb+gDzRXwXCHNmRqxzTeiSPw
K5ArRpnJQxmCUpRSMWAAaHXoIjF1T2S6Sk8iIgbDCxxEQInioaWyxO0U4uPn+QwyDfXDMNqGlJVh
9fmrIHCD4r+CmffRH7i+DIvihwzAmB8p0Ioz6Yb4GsKAetEbVTFnThd/onRxUFIJMyhQfJnr0jCI
iSykjYyep0LMrtl1x+vn9mP1uhfpumIa6MP1C6o3uabmKrb9aHXN3dHIwAycGjG53vulLr1dAQ1M
TqbAED+k/zoduzR9p2ugS6DLzDZNACvK7Ilr7CSWXfDiLR+ALY45dTaoAjZVD1Hu24yULc/LhIdw
mlYoLXd+QereI7hVJlowe+svN6ixJRc2d2lE9FbECO6QRKKPsHj8EX5ANG6KAg8ruztZTt4timHA
Hg5mnLiHiQ32+HAbH8UZcYllkiynH+14mhp2KxYJb6lMlaNsTVK0ffbURPpFVN56//cNfhhGA764
4031NBbwsCUGbU5CyPPz+41CSxXqX1Gk2mW4I2nZOOubGVQsqXDEgv5ZTaWO1G7IRDpTk5ct4MXS
E2q+SBL+XopNkm0RQa3fP35e6ARQTawJW3D5dc7rnZ7SO1ndOAZ1gVIzTICWAwadRhYg59ll5wxZ
HCB8D++EfiVxf4UOZ9lztI/n/g3d8w/lqn6gM0/jTtWHEgE8OREZia+JCk12xb6P+0OF3GzTguq/
WFuvCVYKnPtG8xNpafAdeKDhaNbm/u++3uzQi1L2jrZr7JZZmL4Caa7TpGC9t3zyxJ38087zJTHT
lHX8L82hfJTfSgmob//NsEM9R1h4PjgdZdcI02zvHGIps64nRRLrMfLzRA19z5cTU0WXK8r500Xt
BksWn4NXc3p/UtspyXQEjcYveU+qNoMQdf0d+9qFF3kfw8lbpq115hPLpzyU1T3/0pPnu+y+jMMO
7Tgik1qGNRegRfZt/Y4zM3Ut8csNx3S+j1NKRLIhkOBSdCYImQn3EQEV1szUB5ONLDFH6SgytKwL
90Q8sK3Guoa9tgvzPpb0RqBaDzj69pSxF7iUF1VCihKgFEZvMEIZxuZ0c2e/L6WawMht80mLQnhy
qLsNy6rc7Javb1MJyIh1DiguDQE7i0kpKkyghwuSuh0vzLneUqJx7JO+azgv2Zv5XDWWNvzvGW1j
LL1f/L9j+imuu0MuDZUWVNOg58DjVGDaBwn35YMVE5qsj3i2SBaWC0idruouaGk6Y1qnLQSZ98+Z
Iu5wc0xl/Vg0EgWLItC5OILBc/auyOWtIzGJAGRtcbBiLeMCXNGPjQr7exrMSxx5ATQxMLYTIz3e
mt0U/kEgRpNp3gCqi9FBGVleIQfwbAvBFhIK2hQiSdUhWbj8+35zvLRnd8LRMsBT06RbqtxtPT2G
AGeQRH7w/yCzOcPoXJFEe35IshW+qvDnbI51nBaMb4Puolq74T4oiFaqwMJhZs+1FVMY/p3k5XYa
sBHBtQPtLxhYuk9K38//tGkuJH+IpxGRlx4sIGdRDNqEOP2MzzumssZ00Dhh33CDRXvQKnyQy822
CANlAs7rsLMlMrR5lzDlblGxKA/DpVMmYuM2/ErzZoBOZtm0m5hhhqyPgyi+68jai10RmAVGu1UQ
PMGJ0/wCVo1hDvK2uhgnrsY+PxoXpcc3iy0KdDlor5MkhCuTkw8GXvIUDDIjXpzgbffOnUE1ofFb
Hflo8ueS4fN1B/MSBDNxCVvjBgdTSaHa55G9/cGuT9MGhM6nNLwLt9mwrmYqZlyz1H5LoizvvBO5
pffaIpN2xGdyWrYqRTNak8RcA9P0qgMxTv9m+GXuVerHDGklJubw5+/FF4qU+4m9mDqzCRHC0CoL
8lvnRbToyTxd0w65M4dJOzM2fJNKkfNJDW+5jSeUw8SZ76kq0qR7W9lpRV7VEwJLm9T6sVZxnfrL
b8YpE0YLTfVxnJ6cLSCTaPKxFV8lSfAoX6BdN4hLorm5mjgphXS+Frukg5H5sLy8ecmBOTFIGWX+
f3btMoVTuP9KOVmlDQBOOZFR6CHTy2AX7ZS1spermz3LXubV0c6P9zxZQZU48mCt1PUpkop2Oz3l
hXU9VhBrJDTfHTle2eutxG0aO+wwqp+UxCZn77I6+83JHeyNjZ6oE1wwqPrVDWHgDynv9QYHv7Kd
lGl2FRcro02B9T9z8DbtASpuOFhLtkfNkOQJeH1rDvZqI9ofCiZboP45ocGGsumg/R6NPxnMUgLr
dFAzNVpVU8M5uAVWjGcEV65FUJyf5ex87UCoJFr5mJj7H45Z6tJSeYB7ZKTGhMzO3BFhCwC0XSOE
WxNrwRbRnI1hxciYmIKB+kZJ6vyU6IbyCDiCMTR3ZOHptnC0sHgDItc7BsP4mCk4DUGVYHELXrb+
btrxewdiHzPiuIAkF66Vo/viLFeyuVWDpvUDbxD07sQJk0Ce738y54Df7W3pxVv1Q9zdqesqSohJ
OM968xg/7wfX1HJrAR8Rck3gU6M/+QCRskSlResrzJ6m4eKfTMg+f4ddzsjIR2gVhP6vyh7/Nlff
PtPyxSRsyrKJx2NYZoF1PnIzbL6c1GPFtyZ/S46wQkg55v4VszK3v8B6dVvgO8qy27k7HbYVqztf
faX4uAWu1a42Yc+PxZZ49rFsk/Gi4Dwlt2eiF28QrE8DiNfFcK+9/WFpHKLuj+Re6i6Jr5tV/BXo
gyP9gSOO3Y1yBDwyNNyMhkm2SQMRtXnEBnfDFbIrGveG3ndrlOXZHJfvyAX76a1ZXCoSWlMfO83p
bxoZSsznp6L7xWFzJDOe+S5u5XgEQEXctgcfM9R+D3wueiSLRPKPfxHP8LVEqZlLUZjOIMsRzMN0
2K+rF7qN4UT6cfAhprk5+9mJ5pwCy8oBSynG1SwFC0iRGGgD/gvGh2oypVik91n5a31Sf6oiGbAK
5t5SqBQm36QaqBAx6TxoKBLsofiN20Rr/87p65hhr0FhjtHN1wzbKUD5Tq9Mjz0rVTFdkxSL57yV
WRhYa0N0zNSrAF9KKYycluzSCqnUGanCFdmtigUqi0hHJiB0EiYaOKJmQUUr7o874jWm2q2rvl/b
D5LjQwGzf/T6wNAIfVuMZXZBO8vp4DTXUX4Tgys+lEZkTO2n6lOljnXv97VJw6pOEsroIRyDPdSk
dfLKjnjAmOvKTNBexHvq2TdlDOZRVyLHuWh9NMzzS+NwRGBG1R0GYB01KMWbM38fUbQU3vwFK29f
zsAfrhLZO5Z22SFQXW6wYogj/h3/vWUgG5xWrsVl1N6ukdDD4fx6JF9KnmVhgWBX0rneAuDMdBjM
kHnEiYPBl3UupnPC5LHGBP1mv5Fu+B8wfjLRqX1NcyDBRxDPxOkBrBFMci55L9tkdvA4cx6HF31o
i9NOhEajIPAZcG5VYAj29vD5+ngxXdQsoNWvIwPjCvRTb42KFDgTAv94lcDKayrrj7Q/DQlYHUmu
kzBKgSnhvPq9938pbK3id7c6/1uYte6+nVlPTazpA8orrxciWiT9Z1uVRYlx00syDcz3dh8pEqJw
KD4hzruY6lu+LaxznWNRSWtqrIRXJY1lY+TQofAI4Qod2gOqEtyGFjfKCuvm8fc4CtLChwPuyMFI
p2Sz3rh8P1R1XvlKapIwKO6k/4OPlttddp+ecF3MQ54CbM09+Kr2AzB6PSbL5j+XZe17fU0k8TU3
IGow2TKqgi8PQ+Pc6f6zZMnybW35gA7gIao7O4VmpE06AbjI7XduhbfgLmCi9QP0mz0BnIQe9jsd
VYsj18KqnGQvbh+BNWYWmRQ0TCKV0gr77MvpblZxqnopsFfPSNKsE/efgav90qsW06nB/HrY/5MI
/UzdsiB2olBzZsQwirqWmRdEzh00nzXwqnS8CfL/XgTcPpVa3MpBmp3g92b+QmlCQ/FOL6SPUBip
C78dLjk/0DiZ0nL5qLhk8pdZuRrUQKKk7eSsumUvdVW3m9d5Dqz7/YIU6fKweHG0PkZjGsGc4Wjj
OspDB+Hrtqt3zD7/6iAi/co2e1dw+AxuNdgd3woTDjIxgESDpMDca0GJW0nQ4iai5CLmcLqgR94E
NfNWDk0SUqQO/V2l5RTiDQt3j96pTkmd1IR6lhjPGGbpfLHNW0tQobffF2h3eAANw8n7bax9XRYa
khHwhLRTCAcws3wVVopXSanNo/e1gKvDEh8rodMxtS2zBTQI2ivdCdSMVz3INxrLTTkvMzDTN4Jo
ymaDFCIuW/Y/e+xXYbzJaUSKfLfTOuYLJ/7qTXsQJbkTDKzf1R0jdE3IsioAwhvXQQbFXqAVr+HQ
KPLXptFhmHEJ3Sn6IR9sTBFVpeLtuEYc+TUVK4JQE2Z/n5imfxAgOxZJzPuiiPPPysmJTtVnYXRe
qZ2KR0eYb+NMpOHqSJmjy5C9bLEX3jeu1vpq31iiTrzRh+Jw9rPmHjbSLUOOPprbGul9ckuDKPrY
xaYFAaYCTlqziQYMTX0MlNfScVj5DjCHQpryKesbgWQbhcbri/AtLJFf96v2E9f18PRgCt5snU5E
ixtcQODLRifhBXtHLKLpgHBWAbb3JXnr+Lt5XrsWA6PU2SNwjgBK2XIOtpH/xCdY4Sea2y1Fbie7
ICBSihiDVhLyhXg9rah2LBpFSmY33gKuZS79fK9vCrAJr4o6AckdSB07P65aBLKNnmWQOKPwvEX3
lyz6hu8wZTt5o/NH2Y17T5muL1uqjEe931KJSDJWKYRaUoznnJ6QJVkWcZuoRRCGJnglBPnilwb3
3OVcZlXhSsCuqjyR635tyRXWuwrSYTOR6O5BPdJusiiGvT/6m2D4tCCHahxKpEAqRDnnTPAUpY3w
V0ZRGF1QfKL7OcTdehWX9wVEpKsscnUjQ20dEmiivE5mxhdESScob9P2C1I7BDibk6/CBmxZHXTX
HQH02WAxomlhip8s9yR9HrN25lcE18M+FBrAzC/KJVubIcvC7EKgCrHhde1OUFeyVIjI5NN5YFuO
4FAKgzDgzJwXIoCpK0Ks/MF60PInzlrjOz/5nFBB/soJ8MxG9ffZYZRJkeYMXRYufQlg2uNJt7XI
jFVzBVYQvTlnBU952p0liptP6tmpXUZL43qsywuE4NtabhhFuvU3fcrn7OkGmiQEWODJ8UU3N1od
DdC3h3zEB9+7saWVofVKnNmPZwcHMFhs+CUOxsQI2WfE4/0180Rq1ZWpqAeXBHpHlYVVt5Az4Lj5
yV3Jk89H6ucbDQ0Bn4rrA8Kyoukmy/Jk0upQm+Nb9fi/Hn//pjMIc2ZbTasOJjeU2skRUZH9i2Vp
UsVM2qGLFjfIi4jKON6yE303OipcV1u/fFtDCLaTzq6lbFphmLfkZc2KqaJpEY7D6THpakJhlrwg
EenmOycejS7IdX8gYOH+S9pF1IS4c6QuI8Brr9GkecIMDosmCC3q9Advdp8NbqELNZKcnOw4OYnp
Y1PYEiDxSTOzH5zDw+PAyyWscraGLK/bbHEHK+sBnReo0ltObCxRZHED7eatdckxVwE7jU4mRbys
dIwnNCSt/S5s/VfQeVpM/m3nssHkskdEvH9xbdsnGzd6Uo8wMXdzFriEuYSDVnb+j6QSRSJSK1md
BVNdUTVQhsDbRC6I7V47bHy0DLtcri50VXqZ+FCdg4ceqpicxWsEGKQxawbuyNQmJKFivTL3t10A
fKjycJDOPTOQLp7G08f25NubE2Pj7pqg6j76aDLnsa1wAhZJ/p5BLxs04PSO0ehnFbar9EN1rRPQ
sQUjBHhvcZgDnWzTatSmO3VPLFgeJ26y5u93KsZ8kXVDthFeJHhgI/O1IzhMABrfkCfIP1Bm2XgK
6YwMlsJoTBwK3YI6bG4gS1k+riiQhDwTDj4BMoCAWJIBA+E3Cdu0eAFvTF5MFjtEBjU79JHP3ERw
JStmrbgLWNiNWf82mJxB+hGQ7OADMEvPw8QDeH6xJctU/kRyfXEO5ALzEIeB+BEFa6ESPcNDMUNQ
UXKZsNWJaTr3WTVFqvzqF69TsUgtKdsBn6m0V/lLGwJIk31Ai8ZJ5pWx4RolteprrjfmjDTjP5UB
VH5MffWFi3hc2ePVTgQueIPY1ZLQsMOsyz2U2aA54lUo/HA8mkk5qOscIu1zgjFxZ4C9zGaYAh9f
Z2hl5yNrB8wiIqxDeqea88O+kMsjzVof+EHIh7oVqruczeRYtFrkrPQCWsAIGh9V02RLz2YgG4pQ
lq+8FEBkOfigmLRwxsiuhmGjBJY2GFdb/HzHMuggxg78i17clNVPyM+j66IUUAHDnlLhLCaEHuxP
USnFIILkVU4EQPCbUoCM8+pE1O4rRRib5ruC3Ge7ouUeLtNa4NMAd5SanWfSp9wPFJGA4tBTFpDv
waNC3sscc3u9oBwxfkxZC/+u+DVWZezKe4Km0jPQbLWT5On9pmw6MnSZoEnqe9aKFlxl0DVa4CrI
Fw538AtEbJpE+NF8OzUBPLZu2w8sBi/wnjx6iUVyll55Q3VvLcX8Nbcdii7OJ0E/u/lPw/FV6Yc7
OtMTosl4MrPPTXz7HEooQJSHOi3ai0EAWuQJXzdErPMSKcOYANFI677mzr0e6qUEXeJSo41Tv2cC
sKUe8S78RF9l9WrZZlVlPFB0YE0vfU1rPSd5/leoNHS3NxD3ypUFEQibDHu8GoXXhThXdisY14W9
0m7YNdDhsZaf583Y8cG22+LVBSQBvqbpJ6j1X8X1lJx97jyCToI/OGUq8ku8R++xvS9xaLNmnbeM
CgQKUzFovHSOMHxC8l8HOdQaRSSrUp/haiVQma0nVOBTK9ZDHo4O8pAWLYON90SwUKDTk/g+pBAC
rK5GpGQJPwm9kVliAdliqg2P3b16mj6Yk+owVdwUImX0tzV3QUehKnid1d9xEalsc66GO3mYwWRQ
nKUpT/u0wPoeiaMstMERqBf9yZYEvk5dJvZYSuW1wfzOyxD2bqGLV3AWyx9JimRqQvFiuhdYrbvm
g0KQWaa03XU39sq8ZLruWXhOe2HFAP6+na0q3TRoba0gFCtTsYahranXzt3btXsS4ddHZ5Y0bjE/
hMJNllWpfX8ezVMkP268YNU+c1HVfWCPA8m4f8B0nhh/y4rK2pXuXPoDnD3wY9XT3GG2vi4cPe+P
g8VJrhfhIlpnQXsN95V6TfbO0ZDRP0Oa2OOPKFAJso65G5iH7EcRhyibkRVW3xdoJLqAmTDiEbfJ
6INKndEwD80pcceWpzINwhNU0uNAGVrsUnJHfMNWRX9ZRTrIK3WoInd/9UzAHe0Kl2U1eMM5UzN5
86OJAMU8kJgKmR7OkJcRzNhLu0RI8CWhF6NCidNHAtiC+rwghdLqnuISMOZ2Y0WqzVNFgTeXGK/w
zLCOFNUFZfo645f0wGllvgngIIZY95MhwkRbKJ6zFWAv/Kom9+Vz+TjovVoRi8mGUjx+pjiULSkw
wM2GagjQyfiE3utwgEB+uaHs+9hKy5Qg0EOMvEhfZ2blYF1cdifuk9bgxzDehdL/mgphBafdq2Eb
aRM3dzhF2Lxt0R/rzTeHApAcHrTxDuuZyrh/LJJQmLTgoqM24XtRQEgaKUKJk3+9tbhI4vwJhDnP
ANmTaQiC2zmhqBJ0KU0tksJZlddwxutTXQSxzk6Anvqq4Cx+0c/NSbxpFsOBdGOBQmigN0miDTxs
V0u2lVRw9AGmP/w1aUkKle+h4omPtPyhKDaJ8gL1q10wZNSHTPFMUlE9wy24QF7noVJvZxOVZwcZ
+muSHNFiYSEWg5pvAoLliRqrSiN7aqUZYA7uGIZ0OoEL1QqhyRDbHcdjYoM17LNsPodke2RGRC1I
lOX61+3le6s0St5mV5Rel7xcwbvI3wwCpsTE0jjol4p2+XY9o8/PE5/hwuAMBo1KbNqGBQ+6IhUo
soJ9MF9boOpa+XTEnbKeFBskpY+ImNsLpwpG5xcA45330cB4gEOSRX/BGioXg41KJ4pGjBuXtR18
k75SRDuEZHi3Fhtn72t2tULa7NrzaLS8CVGMgfIZEoyuXkQ+e3DdFIEDPfTrOtlwlF1LNpSn9oax
aZxTCN5J4tP675m+eLFhZWetVqwfnnbfSBQFeBAQZZ7H3sosSzkpwhmDfIfk6SHfsx6WroqxMaMj
O0OP+9Wn7WrddGM34AFMMnqqm4KjccKU92+itMm6NA0JH4wWq5mRntIzSfulYSIlp/nfbPaUovZc
wMSq1tkWXAK9wqx4RVfVuF9DSbJaTSiEvc6b6ImLnuWzkB0cGSRMTpIzl+LCn0S4IMggk9kI+qD+
o4RUluBCb4YTPFHNsZdbywb58vzU+3Rbi20Orbzd7DMmG8gpKFNINXy9qkmw78C1MLxLdA+MzgN2
khPJOgybsCe01sRHlwbSOfH57KAvVKyyFHR1S2x3MQREp000roxE68Pn17A/JUe33Q0cPRg/hCpB
sd8ktoAVmFDpYHuLHdIgyQBdl6+bGYilkXKKpJQK7KxJeMK38FtS39fQZP9GovEpkp0gF+skrGGh
nsd1R6mQyYMn4OnU/7eTX0tv+2V5RD04cxNdx1iOnKRvfCU7/G6mbfWD9SvVsMYCC8/b9fDu+1Tz
dgqfQKxFbZ7VAMILkUwTVrVc7dDRga7AtbA8f58hmpD1Du4mEmbmmvp3i7nfQGrTVVFW11eTi2EM
YTOKlGyrvIFdTTpTR8b2fGrjr+96LQRYwpdp1aa4OfKFDTGRqx2RP0XvgXtGDjC5QfEVoBrL7+x6
IKcQ+ZCAhXk2Q3xGzeLI3aJE5zWbAe6Y6pLEwdmy6N6Lx8NzzwUuvEq4NXWrJ4oh81Z2gbG2HNDg
6mywEkLy2t3PbchGu9FcvgeaXgiQXAofH7ylx8bJHiJsFsVhFtcD/VJEX79ppauzy+4mevbVXrLO
2s/vBJcl6tfvK+ixy8oH9fxLFea2brzoX71iJJtLZ1pLoF7eeVt/F1HtycnrxTQQPaU3h9DS6z+F
HV7R3PlWJCMAdlF2Zod78C8TGTmV5B4xLla2IGvJJ6hmNLquM9LZkYvwobAJuOXkDXCq8JhDprz5
VC1Nks8PQ2PMKbhICtEwd/oOd/ljcgdqDfRGg8Q69X7ndhavgDOK4YBjy/SymJDes5qPfNSYHqOp
qCql5nhlk5P0UjKcuVw0mENkEsaTZFfUQk9yhIoSBjK2WPk9aKbGqZyjqatUibyTccOhQ4ZDJkWX
caz0yyX7Oa0m2JibY5CjCqAYMzDxwT4rAaIG0pMV7plTSvbGC1e0hQh+6bzNO2N3uCjFXjArELN7
EDjtemEOg3BP/mb047qek3T0jB+zk2N38cbAQnjsaFsTw4CPmXvW3ZbSLzSOZ9fFTfky8Q1g1vZ0
Ea2EAKpwCdKJzAQ7IcG/TyggXXUTaLiuSDZ8r2ADPIeIgbdANya+ogxK8HRmsh33tHLlCzaDthMc
rnRPdqcuwhuEdPXPcBqzCp5G6Lxz0fJwX/Y5tuDQjKw1vjgAWvPEKb69xyH7Q0Y1zWHYedivPaCN
tgop1iASCJAGEmMhg5EIHW4YzIGY/88hJKZAvXYtMSlOz9NMtWL62ozku2rL4uYH3zBydUqEuXTa
Dsgof/CFdoxYuVLUvd5AoZMH0SF7eia1R++lbh4PNd1ATodyNiUbGMH0VFM8D4eIYNbq7YV4Jw3k
t3sM9iQpQXsJphls59gBPIku1izTVMum/k1/OKtmmgdbBELG35MSsWgDKv5ny2m2fGykDydWIeta
CAJaveadri6S7ztMq2wN/wjTTLgzqnnYehGTNkigRNMoaajF9mIZCV2xAcFP3ZTd5JlQmZDypLXu
k86fnk1Ql+y/ElG1b0nWYb/vlPIqwZ6bnkOd8txiIytgcxwwjyBVzKNWoz15e5JRFcevy6mp1HNt
xLpWioGYT8qXhk7V16FIC99IhNz0c9xMvpQuDIW1qKiLvvqwl1K9FkwU/EAZXqPLWyKl2e5ewU07
iI/yrRL5Wg/ng9WjmB8JTtTyjbZcN3V2K47DDX1GHQ3ELMgsB5kJZWMahO2l//qsZCcBWLuEWuuj
Ov9ykVBNCFzJT6ejLvBqt5s4cR7AHZADiks9m5AslPd9AqN77aUgkF73G1xKriTl7FiZlsajpk2S
CXYdpLTrwxXpmbrRVcoo77j1GPLwinokzY3SGj5YJz7TvDymdMpYxAE/7YIcOSWkl6n+0kc3fKbn
5K1mfYpz6OTBhfHeSV78j+CS9ugKEogHdsTPq0csqWsSMSsicTxHORRdroqceLaPzbf8KoLHwYfq
j4x5bxm5EVPKjv0dLz6Mll7eDEvacZAcVsWgHERd4ZPoTTYnOGaT2OwCZbH+B0WE3dz+Ofb94PTW
gyoX+KFrmzSJWTPnhnNfDG/H7KcKMhztaAIO+CeFqNNVheNKaRPetxrScVIj3qcO5oULITIKk9ek
TsI84liAmcbMW0T1y4UNxMRcamAtPOzd2WWVAY0e4aHPUQnp/DFbAM+c4jc39/tfcLa1PNBIbmwz
wx2ZAJ79o5mZi7QMok9nxPQ3jlFCdAWNxwSCrtjBNn4/Rbwz0VZzvDWkf6JfSv4kaUMoQ2xqGYwY
LnpkoyTXLIK4tj/FsX32vEbdJFzyzTUjWvillUzMsZK8+L+Xq7KXq7/EJ9wIgNp/RATs98/y6A63
S8Vo6fYzkbEhPFDKrT+f6kpZl2ynzPfeu00k4/tfGWfImIwtG8iWvQH8PDLisHLD6UCCNQU4rn0I
Q59DZ34oKtuC3X7mB1qUBAsIB3mGpQNuxYEvEgG6UFuVBr1xl7bZZsvPbz8j6zIBu1pdr+BfxnF6
41DpoOz7j8vwB+nnJ7GvznvEDXzplwXk3uDkuJiaa0LYyf9jQymqkrC2+v1ExemC6PVwl1gAgHv4
93b0lnNMv4IeyBEB5grkVtM9VL/yVgIDYnqMAug3k9RQD+Wqqp9sNioD3KuBuKnVNKC8W2PzRirp
elCV2mDsK+5Ubuy5q18Io/kxKclZ42K7hRvrcJgl/enp7QHUka8EhdQaEAOvZ6w8sHyW48osutCm
1rGEQIwELkkh14kkre3mXOzXdS7iLO2VGXIawXa0I8t4/MnfiWrF9sZGmYCU7qIBBIf8eoMJqI3I
ygKo6nXFARHFGp6aLFb2Sj2K02XuXxBnlfv7tV/pYBXWvkwksYFqaHgSvhDVtL+WuvPdva/5MpW9
RQX9SeESGaglnPN7IxMCJYLYSxUbhzLvGtV0Wju9zniICOTGmzlGwp+YJY125mq84vgQRvxGD3F5
3F7AsqdGcymdyr6r7+Vsg/6pjS3BAQGl4/GRL7cGDvi8RqIdJXCIzg3EJdflBn2kGLHTAXLOjTlG
ITztENau0eqonNchj2Ry6rXqW20hoMeiUztIBhzQm3VbMk96A1tHfSoccww0S0+JCGGKRT0EV3zC
ODs0LwFDFznTD1eUrO0HqyXMNLl++kcAFNxfGHXFvHuXkBEXjRhiUllmohGbwCJYqfh1tok1g+tC
1wv1lM6nScSjayq6/FjtTTBj0LM+d2ZLY+cg64dpc13LYRUNEhQBPkR1aQDNeTaTjHa7xgZ0wI4C
fu/o+QZEmXIr9qtuQOJIdknIvzT2/v/emxxVpMyU6WsymymdV167v1MUJxc5yL/Iv7BPOUrc6cTM
e9hgmlYPGsoBOkEN68UOKQ/llmYEHp0LNB73FkTys1W+oUbieYIqHxIRtkvGS3IPzY3Bty8zuD8h
impvIk7wkGJFLOkWIUrTYfzzN2BJcF3GegEa5EQdxQyis1pCA4k8Eu/86zyXIE8T1RNkBwCzwY27
IUJuLa7nrCz33d+lG/hJ7060X9IZaMztU/CtghNydqFY1iYQpwX57e2enNTUthA0Gtvad/ng+y1X
AY0vyK80yrZlLHaLv9ukO/oWU+KCVuKvM42+XTFvsHpgWesn006fj3RcPhhsWIwvNLKqdcDuzw0o
XURXbwbh61IEKViuGGLMC1Qm1ejzCdNUiFqPnqrCICe23OMHbVar5aQJUZrhxgjYboEvK6JVYnBt
OBkqi43kkBbbdCKfTJq9AYBoyyQxVnvQ5T5GKPnjRFga2O59y6pqcv5u1mjSHQT23IiNBbCpFu1n
azcq3NJ24DoyIQjmUOm3E72I+qx4R7UHQED59EpW/53cf/KxpMK181YVruxQodZNIsPs68yckJWy
Xinq98ea0vNTVPs1+LamfjXHkvDw/o5jmtQsePoiZUb+UrpN5jKUrnFIAwvqxQR2wcPqUsVR0XJf
1mqwlJgOg/BgrplfuFDsj/x0Aq7PLergW2uCaMKb1bANOHNNFTVxlgBuilaebZSKXhNdOg/FxeCZ
u1E+M7JlRFCKWpQ65Z+YKvwA1KieTIhzEKkCQ3roEbgibjYnRVizNZEyNvTyU4bOffHn9THueUap
Oyib8V0cJcl7blmF4vggTZnXVk+Bn1e0bZ7O2XuWU5UTWCEz9qHt8IMdRZ6qCUth2AjA6IaZ6p8z
9Xyp/RlhiBgYRA9GAlB5ctxr+NkSsABqNQEntdfSJp22r/8Ne4KocnsuIAwq7P7+5Lm7crMjdIjn
rXx+hDOvafvGhW7brJcOo58Ycv4gN9q3L9bBDmBwlyTHM13qp31da8rigRJlSXyV+YGjzYB7GCTR
pZktNd4ZZJRlUHWbC0wf9jBRbfyaMTCHtmZ/yBcLWH9YUXt1WOI40jfUmy/wQNhpF0zyLj237i2b
kVZn7knulm3X972so/A1KkFkYk1ZEhJOek6hE/DkLDeAEW7ORImEFhfE8Vhc/s1VEkPTXaEw6+SJ
VDKDHHIBTfTGm12bywJdFP3F0wzLiGrrNWaMMn4EuCh1tFO0eO19marwCczh8JQFU/OdW07/k7Tk
bk+V8La8UCYE4pQOR/zrGlh8YTjKkq1X+zo0JvzAShSXchE6v0zxJYb3rk8F2Pr/wO930VxC+afh
pO7xuMotSicKi07t/sKzLgpCAa5lI/tp64RUeN/xQrYNgV8JAbc8B9P2XM/4eq8wF791hoa0wzHq
vQEstOmiIIjmP08SuClCprKhHkG6yGhlxXgSD29Ur0mO0cblWC7A6iHQ2JiwWLl5CoFT+zMsLeYj
RJQiehAXeSYGd+Ag9TIt+DBuUlu/jWxNY0G6bzqvNiG8dL4aKri6Xl0q1sK/s5If+g==
`pragma protect end_protected
