`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 139136)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9KNavgxBjecblo7CHyC127sc3Cw24XMHaH0+FxRAq4ZSokiUCc1dHfvh
A9bAWDNRgVdzGLOnHTehYnMppMM2LME8turcIHnBnrlEo3bbYpRKkjGR0JqMCbcZF4jMFxLTVekQ
1MwfmALs5isoDbG4TCtl4UfNJDK6psD2lgZO6J0gnnw11PLTdwW7bNwhbgA4XOrwZkeUVA1HeN+q
E2ByVh0jp4gfkWq0boF/DJA9q7Ow/wRQEsudOhJDHl7brRxBVUDKb2kCfiHgW8fbDFRouLyugbEa
1Czyof+sNLOUFTlL+TZtcND1KgKwqIYhaRTzClg2a8x02DMBYOtHyyHmDFMPF+53z5wREU43xYCM
BvUQA0JjAC/8nqyi+ETsa5/3BBrzdgYinjINFF/lwPd63j56n3f77K/kalQX8nJrk6ZD7pHRWcWP
uN1O69dya2/fdZGXHkoLIVXWlERlz38VI4FFZFK/iiFNYGTCMbWTZ7I3YjvkUj1cJ+eKUxGZAgxx
ZGqMfEKaCYnTia1lB9B/VFu2suiohKBXGUG24ioapqrOl/fibz2kuaUJ9DyBq58OtnAgNRP4Mf48
g87ICwzLjZ6qTmPpc4q1CDi3Jwc7ALkLxd7CgHE1k/PMR0OFSQvoUcaPcGC8gHmeCw+QC0f+sxyN
bSmDtd58LqhjjWGiklsAOMf34cI66nHp+e+akosbIV5lBIL+4gVmvVc2xB9TedIJhEczcxFeO1eV
V9iDMdU9s421QvnoQ0Muvmm+9IU5prtV1zsmYLG3uGx5qBRwBpgLo9E1RUAfH68PWsdL3vqhGoxo
JOGijeM74A8Q1WgUo8wArqSvRBnhKmTUJR0gVDA9VxV/HKXCxlomswgzewXvDh8ecXb/Iflvnf+2
GCTCZcc0hlWSuOXIzJQtnQmgEg9nJ9XHa3EAbfstL/NK5qBuWEJcIMwRCdrDqcWcWj84RvlrG1n2
wQR33EmVgxBhG/JLIqy8EeKilSZdVftl99OmIzAVI6ySqw2tvhoHe1HWYNoI+CCl2WqWdEPe+rVB
h6aiFyaGKW3sIoMKwXyy4DOXk7XJMBefxdtmG1vYAsst4+LadxzlIVo3WmwbJ+fBP4CJ/Ea+cgjx
8odMnGD8yXW4VLNGpotl8MqoSB+QA257BISQLO+N5glWrYLc/oMXN8/XqC1/S727L7bRXCyHBgOU
+Mr+p7joyiTq/LJnmaPGxSSHsTBaU3z8udyPY9FndAP7423Mlc2y26PTKwEq3ajFoeffdTGmY7qq
AAfsvCtxUxHtYtBb8sixT+4adjEv0VM5sZnfakEeYViaxd18uG7NccsVGZP3GjbiPLuvTTbO98VA
SHdwGx+bss6KLTaMAQoqtH8Z7u3sKUintgQIznrbO4yxsxjznKGWqIE+NeTq4aBK1R/R/Avz76HU
YTfkxSsU0Hj//h7XIsRD64928rFGPUJ8l4kP3tdgIDIecDk8CooABGD4u8vFoY8j52O0KyKgfNlE
xKt7lVJpQZLp9TdFq+fFFHSaVeGsFD05pUE7KM2JwcNNwnej7WSB/WyRqi4JsTgZBpD/4n89eaQS
yqJNNpQiRnKzQTXHuqE4bZ9eDmJlbWvpSaSMp6eFbGGJsblnzC0pNnYWWfY6zukhNy9k1iwuY1gx
l7fQQUihMirljP+swql7paxYx1Zi0cevDfcfcrjgdWQagOTczSNmNpBEN7durbnijViLsZUaJdvt
NCZG6ccUszVmgb1JFkRfW0eZ+T6wlIdkg02xA6XicasrfaWEsDyPJCiQj5Re66PIz7O3O2OkV2i4
ksKy75cC9tU0kb8SiNhFj6U474jlz57yVO238XHS8kGynMrMXTyse4Y2Y5xBWpOWyCv0M//weZLD
NDh6Lm0xgE0Ivw87+g/NI5oWQ+28c9/dk+LRXp5pjpCPspwyyILmaY7SUHTckMBwvdc5WYtluyeW
tXg0UyW251/Fj1uu67EI9xoKdIQOOKSUCEIplO13vvcSoGaxqHuItSCdXLEEVtj9o+C9HAW3GsWm
04fYb/JGtiBPA8ekpiKg4ZvqlFxHUS4QxkWxHnRuHIkmQlRJH44exYw5khdyOEo7ZR0tNjCMmhuw
4SPRmqwqGZgIO6FugMGTyeS4ZxfrQp5mgePlCrrm/t3FNBu8HOvKDU88CXB8cimZwl9XoFojpTrw
0z622OcLWziO4Yxt/i5QKv5piOYy+8Y0FyGUdOpvHQBqhe2Yd97E8psiulPU0UMXnY7r42hh75MP
u6eTyOAh+emROW3eZq4Qq21YY35Ey+zK6ZvyVFj8eXOHQ+rfu+LT8X3v07LzP7CXqAd3qwkV+bKO
cWCIZboO/1b+vo5beepD0g0cq0ENnQQJ4w+A36S791s9b0ouyNXyiUBvKzgL4LddJwZb3S+2l6vC
h9GDX/l8dHto4nGKxRBNU8H4hIsMS4A/7ZMHjjhe2mRhV+gr1OrO+g5GEgRjwtC/s7MS/k+TGyec
4b21FlGMcq/z0XmpFE/wJtmslkM5YfAQghz5DWnwxHOmEWWLUUwV7XqcRUEa26D2g+3WlHgG0rEL
ZSdhbvkxsN/Z0A9VhCFHNgt+TGCGREjhNbweU9F4qR63DNX4QPraVstiWs+LNIjEOsDb1iAWOZyL
kyE/Wjy3V9DD22fuJgbjrhzfS/garBKrhVFu/tvClZCtH1F2AAS/OvuK4aUtMDU+lv5WedMOZLec
nSpYKqTKydGb4GFD8XTt0RRJVgb2OC5c3DYakJIXkoE4W3UNy1GDifTjtos85pf5pao0XGvHY/6w
CaE0xG8/zOhwpW5WeYFt8s2zRJAX7Bxp2U+gy/v/+4cM3rFdoyx2XbUVRmBpz6qZnr5UFTYpoOIQ
5nduaoObaW45OcwhU00tYfPq0nRIrLuFf6mdwyQg2EbaJ/6KjkqPwDnCIWkuDVh6hqd95cqHZyhv
6t8+ccK9u40HONvL1Yd6qruLTilIKhj4UeG62bTrXfNb3v+DcwuYho8QiKHLrW1NVGdaQy0bG/XR
9VHNSu5g9eLGTc/cMxwmP2a+s8+dYc9H+PVygOcMa3yiA/Z+V/mIWVxPurAWlQnw0+Aw/sDsBokM
BIjoUjFDW4QVFqT/z6YkEp7Fw1blmT5/M4M7Yr/KZ4pxLKDYVYH+M3wO/b0h0tapIDHUTp/lzqAo
ME5tPAwey9drfVzww9/U0kZrArdgBK3oaA0xOXrz9WxjymFZR9cb+ww0PuzkVP1pT/thUU9PZ46f
IMQ6uSTFylTBEDuseS2ROGjEq6Ur6iOrnEweO1WgRlc1aMTxHQmuINa+zRizYxlvHyB9ZNa7CF7w
adhrGRJqWO/TCY1/133WfRGnP37xji5DJeF4Rtd08Dpk3i5RVMwU0bpnMvfQYrtOPvTiLxnBvGWx
JJbUyG6Rm2Qkf2G3zwwGh+5UjsjNHbh3KBtiqrx48iiFtAk9ggusver6KEg1/6oYfa3k3jqHwW/p
gOp4lICPJvYVeKdRFn0fevUUGUR026YoRPlfGnJIZWHLNnMvJ6SBqeLCzK0zffk9zfzYeyBc2rGW
7OqTjbrIAjNa/PBBCVDonvxcH/rbMvV78VhAGQYskU1HiKh2fRSmpSjGjwfrOMvtml3jakZJM95M
eUyBsbuRUz3aeQDWFmYyMqs+EPg7wQ04oUTycqJnX40WhtzAZUlKb0Luktl2gFai/U+GtDPB/dkx
ladd0Wh3++zeNqc4s+n5TNHhZC/AXqO8CkV7QAtNf4aNRnjrunbkDzZdT0/d4bSDyJUFpcYb8pNu
ytN8NltClaoF9SB4XN/pC184TBnUToW7STE+vCYUu9V8/7vQW1a1njyL295AQ8F/NYbv9hEkVQCY
Yr5kPhOd8Xiztc8hY1GKMVV+H/9pwZC+Wsjw27HXlUQGx9UbZ1daQNd/2Uxw2mm50512fEEQ4TcW
wIievku33r5A8BEskuhwMRuVNs+BNykDjlhgNcD3RtPDTAb51GeE2staevJsdt5oxVV9Ai6ETyOJ
G2IzAbXAtkIAdS+EZF2BHSXB6sr/siHq3RkuX+Akrf6JpQbLpad9QG7n/hi0lFR4NWFoKk16geNI
1jv+wYAgcb3SuA8oC2K5rZ1655VIpr6kj33dqv1eqpcYiBRuUZ8r33lBmXjZg0RiBlZ5UHfWRk7D
NmR7GA7vBJtKUz/LKfMvalB9udG2f3Nt/sAyr5/vfSevQWQ0zPszzjj4zVR5exm5qKGGQpQT7xyP
Odq8mq2F5GTM+S4rhIjgt/BQ59FgRAy6ccCvSIiJ8/lHlqqNi5dnsAVIl2GSS393HsWtTsaOhPT7
1dbq8UpVcVXJaMo3TkSi7yh3mOTi3JQmL8M2AG7mdsfxnfYvWC4KbyW8BZOKHGu7NPQU0aELpm8Y
wpwbNj7O8NGFOZuvo51aED71d7reXNLVvwg2ABd7HZGCpE8nYCRcM3y+e51/A9MsT3XQuLcUkSk7
agfEWWyo0PZU6Yyv9jtNSIPgPIOS483C36jLmzxW4/Me9skgk0bV8K+TASjDr6MdzLcDM0dPK+EO
RDbI8SwidDR9tyIc9gRZJgviqTuoFlwkzcrM1GLJ4gNlPl++/IpA9ZZa7mvVk9Pnv7qeoyt/uUlC
bOos3cVgmKzPC8Pe7t41uST82z069A0rOMHhxbnkqNDc01UaIpU0vPd/zDUwxdMLQFmeVUTHgwip
rM4E+rZV8+dYk+eGmaTbcja/OJcYdm259wck2+xrYqc81ZJ1yg0a/Isn2y9AgjEjlJWpCQ8xf9A7
+oaH7VKqYx0DSnbpmz8rsKGK58OLKoLKqb6sJsuteP5QxI/mh3P0ml7j7ngUpyMM4UOv288M6F8e
HrAeygvlOGe3iSyWWSD1p8SfAzaFSmVSxspx8oKvIxXfTCYLOtpqVrR6BPJ5HABLA2l2fMq3mUoY
SJ9IS4YvL8xZMXmysmfxmUHEV8J1cQeKdPXAkljkBkzTXWrS4dqb+GwBFuLw1NVsZTb7+C/VM9mp
bNWdCQ7ILdzAatkoD6kvQz37TC2EpR+EkWulEhElqTIQpRv8Imk4L5+th94xwYWBP69bGqd04uv7
z2e0GYJf7qTKfawauWa25kFATaUJy0KNc+EGZQzBDr5rVwGxh+nWfb9I+r0XHr8vQs6mGqpa3HF8
JXVav6E5qp0arsr0zncC15J+zC7ll3tbcjKa1MgezSd6X6vuU9Ox2IJSGl2CFd9nIAwi+oiitCyL
bbh3FwwlawEWMUIrqW3H2QW/n7mEnicbT3+n/ESsZLuNTXr1GXAlc0ZZD0Vj3PL4OCWgGTQBkqkR
FbSxoHumOOi9KA0V9tX09b7Apbagpl9IwZx58HAzv4pKtAZBL6gqYwjLqnNbr6G+Xebizt0dV1ZL
4tqgZo4XT+wbbhk+PcxX3l4m4SCe8pNqHmCtpJwMrGtQwp+qJ5Pxmw+RuyDNU1zF3ei5st2v/yzY
84WA5uGYVTPau8oywn04WTCOUNo6Ioi3Jn3tBBQh41GZQotevZCfCdzNrQzvGTYXmTmkhoZ3jlla
es+rPmWNMC6SH4chrZXZxHgaX9RMG1K+gQ1qAoMoyuoa03mP5Omq/MjxIx7TtshNtrbeB7k0o81r
rt2ttjiq4fc5qY3i67q/CAh6vNS/vszzSrGlUErMzS2TfkAKleCjq8W3dFmAyS0R5ZHE/kbPasY5
H9KCpHZgkjXOjhh9KwCn4sEvSbOUK6/0kJXuP2ewlZ3c11j2xd+JL8chkWlCADSR3O75chOGfbRT
skoIqSWIAvHjd4ZrI1moHdYd0xq2/heCFot2/F+9mNcHrCuzd4+9fFqI7ZZ8v3RTfKYFRjJnIwSE
sXFw/uPhUkzkplhWcArFED7fBjps7xvV7qopDbOzz5USLHIlZHY8WDUfHNkcXYd2vvvmzv7QuSNj
eM8J/7oLZZz2sZis5wcnZkq+ZGA7eoTdl5bvcWTFPmRhQ+B3i8Mt+5WmAjn3j802I5c43EuNz8wZ
ftwtnB04y4uXOc8Y76mx6fprLqLaf+mDgM4x/6AWeHBUZ+ko9S/Upq2VQezuw7SWYz55+4f58WtG
ANa2pXwFdRH850TI6f1pyhevVnWa5v0s6Cwu5ZIJzQlbG6hVsZ9hCij28dbZk/mdRPbtNsOnsHPi
kjiiMNlUKVOO4fn2hJrB3QiPjZtUP1sj8e4LZ8WbDV4ReSHse6NeZEc8fm2C4SY9LiAFZV8EYh6K
rkyVjPuy3SQOuAY305Ov9lzvsppke2F83ZAiIoIR3aSvFhAal0HDsKCM4jKqb1iX3LTyi7Te4xSB
kva0DuuISFn8olbR5Yli2emyvSKFFEtJ7FzKBIURtwD/aQj56HRuyKcVd1XMkjAbxw4NeRmvRuLD
LdRKHUQUhrPo58ofcjSZ1nTuXsNNIk3wlQ/i3p38N/MpGNoqZpvgYl+1hOlEAfq0Pk2K7UIdPIB+
eo/O4RdfG9czUUd5fJajRTpPje0qD7LSJdKSdzWTgBy6s4PXrkfB5N/s6849+f/RrsWnRKgczWWn
U95STeMWmVVehcoqaR0a8MdLxcUegmRxeMcdiM7KOAoDXMYLWFY0D9ecNCx9HgGmcv4yqyLNeBwn
uY5R6KIUcZuVs7nALSqlnzCP64u6NqFPtBF6UWlKVJsGbwT6vULLPeHzhb6CGkKxJsHt5XTRpDJx
4YFB4gh6F8aRk+LXZriXAaP2g3jY+1DdYAkq1tupvoZ6VMzTKjGrXOw4ht6OsO6nRD5IMoIEcRMi
8uYv/wlACtdY7kNJWPIjwkCfFd5Xq8hvMDBVedagGHxKqijaaonsw7Lcpv1Gu2ZSuA+yx6/0OiVl
N2Vil3LztqNZGfHRr3dvVZUEfup2eUdanRRsKRPNrMd4NYbNmCBVJJAo8cZga4Y9IeSJFF8ypfZX
EckMiWHjo/FliqQHRoKcbQ38omSZDjc+IyxPqe6EdhtZqgHlz6ywZt0vD7aFfxdjImgiAjqvxywo
eDD4IkXY+/hE4NWeGOFfFSNcIUSfD0zWUdlsg4rsaPz4IvvOWbzNVmCdtUVp04THPSvAnro1Cz/m
Y3vDgySRV72btC7AD/1KmpeoAyZUxfLt1scilZfJ31x1abMj9/44XYybDwBJxbBYigOxIH8m4gjl
ZSSRQemo4vv9nhqqmgOeK509+9QPx3ALDmRFqWxvXUIrQsV2HFJD3pKHJQfGYC6ipgYAngC4t2UH
N8onsLoIR9cqCBeFqMLMqQRP+ZLYJWJ+iAJCVNxS3WGoLJhhVJgNMU/FMjajy265xaj6XdWWKzf+
4/MciHMjXigcJMJ7irfGbhaOFY2Fd4nvfkFdzXiN/K3X+oKxEUIj7vbetzMJXnFeBZsJUw3ifx+E
kJQqgU+25YqReca/RbsRgon4ZSwxcWx5zI3g5RWcBsR6xkSVwvo+Wk/yRzwYr9/Y//UXDOqbB/nx
IdzAINVGG5+xHmBlaF2NyEW+VfvPnODeCqGn4s+rVFo7APoO04SWQFMtUW7yHOzXfHyrYjVMSujN
SnZoRFwgV9x9n4FIg9poe1qKEAgs9Xb9c7db6kentC49Ak44ezSnCbjoVrHyTyHydqOf09zF6bjY
Q/NJz+4VoqlZzXiPEWRWWiwPvYPTugfX4ktJ9f21WmGpolKoXpKxB9HvOCwMxhHSUUIrXPEOtz5F
R4dGwQdFb5o44ak8CfhEfqTuvkSlGKm/tBfqztB4Jtql/BC4ARqEjg6TkAsF25hxidChI0cOk9IF
aTQ6FU+Hjb1sFY8T8Ewpy833voI/x8qFBlDNXENJ5VjlM1qYv1rkgB8yrykEH500uk1b4J3w6A5t
ts+n37DoO+kieJu9VrymaCzOQlV99o+pF5nWvjlcNFCizq1bSS+v80fcXSeD7tgB/+3b0OCCNwGD
Np+z9Q4TkXto+pIhJ5SaaSAkkHUTU8xYzlPufDqQ3O6L18jLM8Az6fVmJ4HQKBgaAACehmDTooTG
Ubxt5+RhTnYsiMAs5Tq8V9F8Mc4ILwBLjUBJzAf57QCQmY0On7jVSvzssq5aDLyr6UkfZR/1fCvP
nN/2ekMdvDhp/tZIm6P2bR3hkN2GMjGFundU+7qo7b/GY6dqnk3Awhga/Oj7SbEYZg2nl0WQpxf3
YqfCiviCC/qa/VFWcSmV9LhOdatk8jaKUtou9uHTLZQfff/v5ogQvzLl90ipQsTLiuigu3PB7SpS
XV/o1gkTJ8J6pUnoglOrLK83ePqd30J3eD+sr3vmjszgVhLTIMzvUsha0jf26mI5DPG/51p2bYXs
fbQ5Fc414fFGLXtEalxGHSUUU7ZSwr/nCySDInFjLf8+1JJJTj9LT1JZOQDh//sxIB3Q1+Uof1Ny
43I91ckx0SGrZ2BX/EludEwWHOePKgii1xUWNxLI2TcWl3KvGVDSCB5egExZmVCYbTRvEYj/lI30
0rJHRIfkQVDiaOLQnk1Yb3KNfi3IZKqCZHQEo1YmxfP7UmFuxcBHLSo2Qy3XWik7+U2KrF76lByD
ENzxe8J22koo/YJbDm3be/1xhX55wh3K0FabUZ+Tcr8s75H+HaonuRzyi9uJEa02f7nem1IK8lbz
6Y9DS4dhG0hRsDsz5cMkUZq5XV1F8mKVndAkxjTfbIIqsGzzacrnMvKNCV9RQa/eyKPuqzfdx0Pi
a+KNlflQlzmv99TFeS9rBsGOjVuXCUuyhJ+Vp3EfhGy6sXfrrQ9pMhQGrfAPesLM3Tay+FvoS0ml
4XbORoxK8diZV05oFkEqAuZqRcIcc2Z5uXPMy3eGx6S1iWSYQu8HvBG9nrTJRWa4RPRHhb+zHBKm
vR3UJ/lr1Pw1oLYtL/PIT26CSBx4do0OYm40Cc4LkpqbvXK4SdsmbBpdxPlUY+L+Rg/5AKIeJCq7
VtoTswL58gzw0ZgqFTTaxZ5ZZNrnhukQ1ZT7HIPiUDKCnAq3l8wBDffnSkz1dvlwQjIInBbemgWM
55QqD5a0L3l0d9YMWDcGj3cJbRMWnTy4UphxfU0G86QxPCsH/yRgJnTtV1K00JKD4IxJESpQWAGE
Ujad3jhDJLZYKmH+F95vbtM3ACY0V9moKG1QoXrXrxt1cnX6XtzHGNIoEYbPoBNFPZ0JUtKE2CAH
UntgBnbbTwNN6yUB0RQS9utwljeF1ej0j3MS2x0C0Dlpx+4MgczwBG4ptRVdpAZdT0S3VlKC/6GR
TkeYzvdoV6din4dSpeNzyBWQhgVIRpHZGm6tJaI1U4eMaehdAe7LT6vGBNmliUg2WwyGSN3e0MxQ
InzyekKnKit3P4kQex6qkN2tHU/sjkgct+GeTmIrnD5gZBu480go1r1627C+qVpBMUsEtYVIe3bH
abFghrtpQJOqX0kcgMND/S7DuUX7p9RH8PIGjZKIB/vsiAnvSY0YQQXh5D5of2tQdjxobTCUL83h
vannnF8AGoOia/TM0iaZgCezliAtXOY3Llpe7/QPJsJw1W5uSc+/2UI7OVi6C0jlZjmYOalHy4Cq
RZmVk6f2Ou3zV7S+AV1XgI1WgEZ3Jl85fM+w8K2OGvnbQCcFhSENHiqtEKyXCRaPfbzNtcLKjJRT
UlVx8MfExmHKCXRwHXR4h34N8ySNVFi6GJfBxm0cI6KD1+HKg2HZqgNZyVh5EGOMtbi1c3fMRDrP
mT2UYUDGPXU0zgHSdvK89/u30sXJrnB3hLzlNJG+DAw2LrF7myuHbmJRkioseonYqEdPEqXABTR5
8UkGjsanmKZgdEFneXoGP0s1Q+A0fPk44xe9wUONpI7T36k1Gj/DgP/oDnzFRRZpG1j2Is7UnGAO
A+Dof6rZcBtC2MXpih9ji0gjvOIEI6GyUitIDwW5R4Hova7smetTKKgD+Gaw2Rp/pLKksYXF7CEq
L9xi0b401pz8YWsHXHe8Gz9lT5AwMJJf59WioLcF5h4IYhf8yFHYaboUZx5nINxFkgEcbyDZEqbD
Xiif1t5nGH1UvXej4Tq/REPaZIGfR+KCNF2hnXGZp8hsxbV+hI87ir03ZuaLI+Og7rjhfQXqOS0K
30E6qj4oVUQmgXQDtYTdVM9awqIZCG8sFuZGeCMQjno448xbwXWLZFbv0fKkeOKuIBEoJ5B0Gh6m
BaY+icYP/iQ0nsAaA8AUhCu+HEbuatf/fZhLsZ1xENJmNwMG8KKQ7nzoECgU2leNSrRJNkG3lxtS
Q0b/UXMKaLy+P2b3jbibu6f5WwOkMYEfpurrau8EYVNAWkwHiB24xPchisXWGZaKzhkxIxAz1sgt
YqZx3BVPtFLT0vwTIOm/tgx6YLZSlr1mh+HVQQnI8IF0Apy24Ihckp+8txBsnVnIDH2TYIJ2gtc4
9wu+h15uWyUuuD1wcWanW5bvN3ZovH4MLwmkr0bIdB1KkklpZ5q/p8w1Cv7u9NKnuPWqn5kPrJVE
KKFScby4r37m9PEoVHPbEfkv2fEgie2GebfBNU+RQjyyVRjgk0vNgqgS+HDCpyTv9A+8efFnwNau
Ux7zDldi7e9XGVAkYhn1gxJxtWOwG1tKTFcDgZFexRgC3gfKgNjWAYf9DatpvZHFpS7o/JEEnVaO
eY13WYfIofTUBfSYYxYdia3uxqQArefERuwPd2IAdefy+PGpwho4ezPLYN8zRUnXC72h2kuHNilS
h+GXiXZ4t1MepaKbpmRMO0un27RR6/Bb9ttPgJIVeOglcnDkC1mceybtFW1dQNf/NAjQMV96ySs8
fcRcovF0hGsrNSWPyaQtTVS6SaUrdFYU5BJdCXa8GLKv5KmpWNeYvX2g86SGbekfCAK9WR8CVI2/
9Ed2BjrXvrSrFXUPO3u3KrBxk0uEDWWbn78h7mWCnC+8L/qUpCDQMmaMudHtTYJxvnH6VOPg68Yw
LtjiEpGm0mvKBFSlMsVxy4yb+haug0emQvv4fhsUeKvBtH6gulRiIlcFkPGDEgHy7PP6c4czdi+Y
pcW8Hxxa2l4KDDH9kdikYhH2Ah+0Co/5FwQ9ey+1cfk07KL/L3pKZxm5a9dh3xZ7D/6ulZ/XMiHJ
HZdLry9mFbQL2xLOpJyAUoUN9DVpD9dGIEAUXpXHZyruDlKBe5Y80rN9pQrcqAkU1AmQZTCnMvma
Smsu/R/lOFYP8ceQM54r9kc6C0+82HE5AWSLz3e8mATYIpiR3BJ3XgftBYWSmjiX4+qeLEJxbKNX
tMzYLT4OTWrlCkIEc+gWVDNEClceINxREzgO6I84Epi9OWWEhziQ7Kls/pTEWFCkjTQIX2TrKxiD
evTMnx/KbhWIqGb+PO52+vz9VXbZPzHPLBD5p5Ozo7DCOPdF4GTClZV0QxotcQw7s7Wc6UzgUuBK
KDFlvyRZubUb/+sK6vzt6UWnZq+qCOun7APlyiAqKrvTcgxnycBj7g6hYw8zldVpVDB5EYSU3NhV
0Dl721a7e+RYfjp3muJfJ6j7S243mOBCoIwsbr5Oohi7TP5NVp5JYUdCYMp2V228ybMpUSdII0pZ
qTYdUXY/lGp6EgpfY9Nnp/RETdPDSVmbe2Wo/teIOaS7CP3IcMZQP94y4nU+d/+eGFVJEiIepUrp
RJScUc0eeQTniB9CtI//KYukR/w3sQ1gh8tppxRCQNjYvORJG1SpoonR61BJYcMhG+oY4caR59Up
RgPm+pr2GQlHKFbQURQ3qGa8y2AeOuc+nP4e2VzAxrYAjRa3R9DdQLsvbeeTPAW4uxY3yPHnBSvc
lBjIYBm0uXUnbJqfHuk7JrBF6m+U8WQIIg8R5P3mQsnRGJidWoiaNRU5e7LEj6VdoYBKK93Tlgcp
9CUoCwV+WfF0/4R80G2fHKENqxIgf+E+2y2w/PAdQOjgP92FKUcTarsuPhR37pp66iMM5Gkvm5Ja
crNYsKpyXQyfkyfNd0lY7szkBxyfFsXe6EmU/+u5nwIndBVY6AlRBnTq1/eQJ3ZS2EV14u2U3Bwg
H0czXbf5SbQ5dYYtsHMy+yn9CiUfCvr6cBUATQnnlOjOFjQ2CAxo1AmZPfntJMZsM3aJTjJKWGBV
TorNOHcKbGA0ExXIfH6B9/Yh6yJOf4BgjWcCNw+MC2B2yKezqxhdt4R/UM3ADM0SALlEysFBtrVF
HputHE0E0NnZwn6k+GwzOMat38cGgrPvHfAJx8WvDJoDQXqCS2sRfaK8AAiIz5xMNjolB0fcNJhc
zLsyfFkwvcCGbpY/wVPuWGnhHT1fHjWNciLfZiI2pEU/02olg0HBGkByNwCvQqHoHNa3OYTkjswF
HvYrxuoH/4NMM6Qyh3zuF37MyY+GwSqyg0KmQTGmcQiyYgg7aXVnor9sSJiaLgX/KglYDMlgJTKu
r+ZD61AA2Gc1RzRPZyssiaPGhCkcLgldSkjUCa0mltn2PQQIiLNzhI/rYxK/4IHckLevRCW8SbQv
9itPFpx6qcdG+YstgLJ8p8YZrYgH7bUtZCOaP9dgIpWk2mpU3QDAL+T+zIHmZ/iTQlNFHaBV00aI
3g5GbjM0baQ36BE6XJg955Hvw/j+YCFnc3s85VWqdFe0FbEHueITNLvvAhsQO7f2HtxNOU+BbYbc
WTEsjNGPBx0AdFYwJOha9QyicrtH+K/686H1klo+AhhBsFWIqRWpghFgwGUtoflJf5YsV2nbD7RE
WDGbjr/2ZS6Bp5tNWlvyun7cgr5QnDnYxnkXOBxc7Cfo5i6B4MKALM6q+jHPaAahgu7rXUDGUYyP
PJ2Vwl4ZoPqPgqj/uGRqN5RqfitQQHQsApO+CPoQH/Uo4aMLpDLhEY4XTjAiPEGwDLd3B4/pMYRZ
c6y7dDyGUCRkdDIsq1RBa+lnb/8c8GFX60pfHz9ljXIKlaZHWLVjt7fK7j0yQ3BlBA6hRAd2A4C/
w/xgfBppUL324LI6CIkGeCB03pd5R+8DHsEkDBGh0dbaLVf7OoaiQmonSeIMmkJj4CwDaRuFFvH4
KjIZlli681ApOSYuMAqaLxRkw5s6NLXtRqvFwSUJ58JMP+W/4OM9eMDZsYt9PyMy7tf9mik43HDL
bAtXmEcaJdoprSWKUZ1GUOG82424iqJYse72LsknUxmlv8uvpxyd1I4SilxPh/t+RBpAnarXZ4ox
AYe71IN1wNKJFMsCO2ANVr6SssOB5b9I3F/XwdQK29/5Xdg2kDTgSuiCnWc1OOwHabYat/geSkex
uyBaZw/g1dKCEsL5ejg9190xyKWUUUB9ltwk+r7q5rKewPNTClmMhOIU9Jx288uBe9cCVAmPx/WF
+ZPxT4XndmM46C3apvok7SYZoTbUqLRIgBrUcOjrgcwcdc5EfgJ70W+toB6RFan1DpooSDkUiDEo
pADPrD3Os+TjuiydBJTejACW7epANtxmC1xVvDxU0aJEVmLQKger27y1E8fIY+hud5nD4sm6tn/d
oc0Zr0teF6mYFG6cGbM1bmnFTmp0yDAzTDcfyjCifPrBhctLHBo1CcKpzYyXCgFUjUhIylqVSmuV
mJrD/E6ec/+P3R5wiF63kzvR449TzDfcub+8Y/xQ1x69G3W81L97u0cOs+z+1jQcpo40hK2Gm4Yv
e+ns6Mx2oKoI7uTXEsPFNxsPVorfxnZUwGkKyllZiessDeRmjxQQAoWdKE7zZ8Qn4fFYlDtc1Lkj
1wQM5ZtfXHnkuWpqe7iN+dLRqMVFBt93AadXQbN+wS7RuoKg4w1nt9EGuYlQW6vLzqhVF2jrP8uL
p90avn/BTEOkdZ/G4QQZ4obU6mt9LjAM1B46r8FtHUjqRbvPyDsyN1vaBijoxYcY2jkQceaO33Mt
U/Ay2g1Xj37Brbxplq5vkpsyxcH/F/vOX+pXg7e3CDoJ3+1Dr6rWlMpEgDWaJHgGu/gchQeIWd5B
fuhlncpqWLObN/eqHDCv2A7IRIBKJHazBhfDJvqXnxbqcpOqEtiFUFRdNEiGaMm79XGklAc7t/Pg
FPKTBpXZBlsKOePZWCvOD+33HddhsT931GoIo0rOg1PX5J4lWHLTOj226s7MgJMDD1vcM8nxb1u7
xfFEATHB1NbalBB/+bwlE8b7WQU9+zfUx7NTkoUkRkEazsm/o61XSOe+yrE9TSAA1nl7oK04D+tE
mkGqjjZ+p1dA+vSB12dURKD6Pz+0XiaUDZ0tsP1F6HnV+ucH7bz9XJ5mE/PoQoNiklKDyyMWkUhZ
tq2/RqKSPr70OfBG3jvS69RCRA8OKwi+OLWakpCByAkFbUnl8rqAWWtU9YzjSg/2HH6JKj2R3EUH
4G514gUDDYzz5wHnN7V7ke7kAdwPieecejgq9rx/NStSYDb91Pbxj+EbfSdqeNUXmOl+e1kbH/pY
hxlDy7c3jFPWqC/D2MPd9J/SRNusRxjkNTOChnorp+clh9lstu3Nyi7Uwo7MUw0mzX0aXFY07DGY
f08+0/JeVi3z7HdLtFbYWTqTUepuv2llay1QyEV7sxuaIRc45zw9Wan6gQTzdg+aN2pCpLu8LuHu
IoJWjlpSiSsINvs3x4bloG/4O/jJYrCf7sRlIwHsUxFBcEAxfoUTTK8kY39lc3svqB54e6DBmICg
myDKPVfpos4YH5oOyNfKcwXFUbP7W+1OwF51y1gckyh96UOAQsxfygfvvmLKNiTG7+sy3vdkPMDh
lmVlIcUk56Kn5J3MQgAE6v0bJA72VeqpUbSQLsiqhYZSRWhl9NqrJmnQtvtnqTe6TP2UKOcIrdRB
t59RchRF9zG8leYBgxugVk3hUsxVxDwElUywvcYmZ5aL3qJfGVC9ALHA34EOgl6oDNwTi9eQg/c2
WK6muMLmxa7CXvOj42H02pTEvxtDNCL2EpJybEtI3fdnPcoP9fQ0pQIPzrqMnE77YeLV3tHZ0BDV
bqYsqbC2220bugIxlA2MEnEGPLVWNo2j1gaBAcoGdtY+M1/PCWNzUIOR6e/QmMRZLVo5UUms71PD
Yf+9fRI8yUel3HvWO5f2oesMS/bxDeNavgwXojvsJS4GrmJZ2joLExjDiMztZDOBgsaapbU7I/U1
wL0WqzRERT+Vo2j7INZygoZtMoKjY/x+IIIbC71nb378af/PN0DHEu427ufbyB3iDRKQDCszIF3u
zNSZFfXVCD+yVxRCoGj6istbvU04MI7oIRSdRmi82QHoAiB3AVm4ZbSCAQmeB/meC8WQbcOmJ0jT
voUkXGlxngTqs53zwRW3a+Pj0cbtYSfO9TndvtU+1VMgsNjk+SkisS1Tgy5IcS7TlpnfamZYk7Vd
qbAzCc/peyzlHY4YUi7X6hbAefBO8Pj4DcfKtmsKah6Z2KMPLDfJ3uf1rl32T5KgLxbpg6mYV/hl
Zo2LNFszpvEJ2eKtwGPp/VvYXDE36fC+hh/iYEsVyjgZ/N9Meal+4GRaoaOJtlFJPML6Dvh3Yft8
QM1RZiTMlvXMrNl+rnzDTOM4xPB4P6nYOCoM/SsWwJwnE2NLXlBzJDllutn0P3gE5ItlS0LoIbuD
8loagjJnsYaqxJjun9u3bWoesFHRu1B0/UV1TZqLbHrYxLdPR8iqwL61x5gUWLCrSkkjQeKEDpTY
1cG5MzJGiedhlTaAF72Q/c6HhWd5zRrDU5PNqJD6BHwYISWE8W3CeMDzGk1Kne0Qm9OB852kuxGt
0m0kvUFiFMCfFBuWFrlmykF/Z9EtIe1y3MpsrPSFhbiofYm8GNAUbzCZbXDJdOdSmLBJAKsoafm0
ITSub6ijGssyeC2RyO4Ohfgd/RKsY7JQkYSNFbJL9xpzDpYo2Z8jecSCjeh1yQpZMEsbzAE3uH7X
kCKmQybVwimvp7mZctPWO/anW27c2iosdN6a+E2t/3qpuar9XCpOU/KzBPnncgUDGngEWickEDvW
2ySvERliNFCy4PnlYLpFBzJs0HWydXo4NS1Qs0scCtNFxt96OiR/heW6Qn7OvHR9/qfg8giMDwls
3VGB/q742PkZ0lNsSQmQZ4kYiCtZssxIM/ubuiFBkafiNfImjCUDGVCFpomybyICjx2KCtgX4gyt
GsAn0Qas0JWV+WX5F9s7K0yfjZ/xJVunnJwDpWlVqdwBoyMkiRdkQheYqOGeOn5a26M5vQDteQ2n
XpAgoxzzTBvEST03T4TIKZrf9CL+zKaKHlgnuzpIKaVOjweiZYHdUGK2jW0fe656iiBcKDVckZyz
d6FWORhO/ucVweOREbJhOHm8GGBTr2HlrjjehcUEaVsIZu1j2a5EWCi0dD1KyXcPSMTT1e9yY6PE
SMn/LJznnWq8U98TKhVr3jeRZyf6RHma8J1fMxXY7CVbz07FA70LxRevy3PmXuWLG+WF0kRM4XW1
0O9uzsCH+CYECSZ3pWR/wQWeePuSq2+48uygk/+7zhHo0s1T0J5oMAzi1q71gfIPKpqL7/mcmVmo
Z6Hu2RMzrhhAXlm02RA/mSN0U5lXrgmjgcnyhUJ5r88wN/sbweE9XJCo0dUCkUQvi0Q3Yn4IECnt
awyFSHbQ5G+PhfRXg6EDKhjYWtAOjULEeviEWuvOy+sk5u7EJHb0dZibdfVFnqj8tDjhwtK+3xLs
fuWTkj/+q4iEOcY340NhlpRfQhX5J0vZlXPrz8NY/kMFhYz/NwygM576ItAQHbUWiYko8HcYevL6
MSMTrIkmhR0Uvf3zvp5yLUpsVKLglAv8pEkbPPAiVCC/wu+cNxQVzap9x/NHQWsDiYFiKn/LD4Wf
oDkWslYKiIem3Be0NVkcrvj2zM3qP9D8FiSyvQrRE6r2VFuK90FFz/kD2noqLkZTE9O8ZefVKvS/
jei3FmlYbXnInN2FqYK/AwVkkYWTNebtOtUi8eH64OAagIL8HTjAvht6b21HX6Z9DrDlEAatl9Vx
n+R9h44AhhOR5epZbwEcV/zHRnu2epEzahaIzl8QNY0PW5p/mXoG8d6SiA6LwiwXRBjIDnsuQPz8
HtmfKIZS7jNuKw/18iEGtX9vHu5jBKfXP/fPEAoO2PZZo2gNUC3QTj1zTCx9s7BiFhhaB0fJo9o/
ksfMQ87mFcthvfPqBlBMEgAk9cI1OhvtdUwJiu7o55ht5SZkgCm/3ea4sUG2UrnOsEkYnXf7pVnh
iOMz9/9I2TWxYvbTh7J4AKM1lg1UTGntDA3mUbIfyUVmy39nJ2vw9gXKpzZRP/nzPA/TTagZbmpz
nohKLjNRlyIQYOpjBxiZ+qH/u3/MmLKlL+COf/3W1lZ1hpR4DpW4uH5O/erCW1pUoZvkQVJPJ/Lq
bKjwQXlAyR5zssYeZzW0jE+WjjEkkN79ws3xyKzjOfKX4njcFpW/HwOupQtLGj5d54WBNz8GJlEf
SoEQGyQEB+jCCnQ1Ny2w7geEuvbjOW00HgdmrledO613dB7Mv8BEaqwUIKVxP7cG9HKvBx2EFgdI
IQe8sCJDk2l34RCzjNe10ol9/4SqoEH2frTuMetnj59KlUm+cYuSHHuuUZCEpCzUaabBsX05EkUF
fp4rNjlGEZUun9/cDv/jS8mAHEXOIVOETcBbQCGAR0ASRs96V/mHy367WbNoxRswrE2Wwhx2yKFK
kLX/JkdWxRzBBWfQafcZ57jZyRrjbQRqo8PLglR2yz/B94kd9RK1J9ki8ecnIIdQQOfYWMJ88zLT
P0xDc4cmHB9xqtX7m1NRJ+BMTExrbsQ++qEWrmt4icYrvjNzNS1OF00hv/Pd2YYisr6a2H9DDrJy
oG/ckOXvLFdc5s6TRsUhpDtkgz6PCm9n9oBjrfcU/Xy2Y3OzCovdULQuWyv5dUybU8NUIhYrlCfS
dd8WcKqyVPK/7Enf9Dq5v4WsUeUp3GR2WWGaBFVYFewsLm6TCYohdRNYrwtJpFDxR68w3WsxHLke
Jwk238Uax7BC8EJBHFyNt73KCv8I8ajP9+RW/KR14nSj6znts8wD77IQ8r0Zfz4O4z1TQm/k1KCi
rS8GfeLrL12CdNLfc2gGcmoxbxKCo6z4WAbOhaYP4wH1legcka7psSJ0y2NmbneN96J1gKEIuw9R
SYVRwvD0k94W3ji504M4b2W7vrqHyE8m3BwAY/mICqANlxXzIUPm70ljauzXCaoYiPVbNvB1kAdT
Oa/an7kXxCUWDVNsN6q+OvBs2xb611Vj6Ny+nmJLH9pnjCSCMj5GqQBKTo286HBbnILMToyhnY2+
GS4AvLa7FPSuzMkhqkY4lthA8NM7Jh2ypkv6ka3ojBmNLdFCUPy/8WGLtR/QP5Ea89xmAFRi2WSO
udRTJwG9ZQ9pOqJ/Uj+ogUSVGTsz3br/IiFShwvtO4/iYaUO9VslxLnHiyZcagka6o86rZvWknft
KW9ctmcmwfv72FWsjX0Q8RhqG89gp4JzHlG6NPtQJY2Yv+fVpXlrk1yZ+L3/5IQO7MLFzyyy/75m
l54RNgoriKBHi1xMN+jW78RlFAzPFDqQ6wAR+JKUPQCj9egCHFT2I6KMu4RoYvKLnQqLI4QN4gZr
obqzHag1dpiIPkqT7UP7rqp9n6np0DpXtwHArShrkvJ7fATh3QxmJ/blt7fN4vB4gnSTrJwV+c79
DqQpgSqR37AfoXdzQeF2BbVGtoQHm7fhpa4Oc6zsqSmWCQ7CTAYlc+ubdV3EHk3uVaKD59ZabgL1
dk22RhWetjxfWqu/yqxIQL4tfOUZm+cugrAMdFIUpU1SopDdqW1eaTZOgnCRuWONy6AeOctZn5jf
Ri3WZv88UQH0yHrb3s3jUXN7tVcX55fT0TrNpuFjh71Q2ATe59XMLVV42LiCCyJISPG4Amz9OG8S
a6SXR63stRlg26mV3H+u1fuJD+AY7ih+84a2BIjJ2Uo7cTrosuyFJ4fFksLkXJqf7PGdc2u7yr5w
6LDzfEpbSVWnfWn9J7fjNG3OZioyhy8yvRBNmF6oCatx/DOYrmSokL2IEYVyKZXg+urLzKkIsapn
VY7yvAcUKDR/0jWBmOyn6HT5Oion7HMiZGETEL93kKfWv+zVwVmXFUYtNuBHJ8DLSv4EaEJ0RO2/
KqHHotVc8byAC6n6ztk5LluiKfII8Ckg2jML75b8zKUsXjnxaR+Lys7J1+ZtudYxvm1G9zk7oTVe
VIWnbW3uQRV7j6ab2rZOIuqsVV7HTbS1xvwlbGfR+9H4dI5laBJzXlPtAQ3jVsClFgBHd4ZMD8bl
wHSStd884EGGwFXpWg647vtndTv9pBZ6U13A63T7di3WGB7tGyjbaMrHanQgnh8McDTPvMF2TfBH
ZLB+z36jLTtPpMyolZ1poH1027rDULI5izPUPWmOLt+mktssVKSFbYzGVhkjWniEwj6JUYK/pMD8
QUwu6OutVPsdil162B7anglg6M/4Nk18bcj1LKLKPrAsR4YixdpZbZZbIDVKOzHWWcH5oP0VIXOB
hihQL1V1BInVQdsDUaS09stvhBq6U0hxpyVrTW0nl8EibDa6gW+4OpYvRh24BPYPQnc2KWbFJF7v
ZB36tfFQxunVlqXKfAQwrvLC/J3eaG84nNhONROizsmDPhugfcfikpQQlchb+j6AI4dpyHVKUqkj
N+95+b7DE2AawfizRGDYP44s/HbQjc3mne2qisrWZ7L4HAK5o/h7BHnL+aejbYS7hAdt8agHRP5S
Apz8xp2OmvhmNGyB9GvpWQiEZSNC+kYVMIdK6pzt0DYkJXZgFu0gpW1tul/ICdNzX2uNL8FHjUe+
dWiLMv4wZe1HDQR9eFMAth5/PvTlqCwB+tHmAzRvR29lZsIV3pxvbcEp+kByzuqClGA4ple5JQ3U
Gasc6RXG/lnXUInr6rchFP4AXF6nw/Z8WFPqBcVPW0tgIxh8SrGHuvU125ysUxWDbPXzmNa94LJf
L+hhRbSGTSvWcUPmDMBBanAtHnfx5OojUhgEdrhK5Z3gnTbGvXrRZwC4kipRN2GDQFbs4dzZg+vI
xWVocfjyOqP4MB64vQApzN+PaahMifImFmBvrAODMTZfQ5qoJv2slOyAmv1WvzsAWmi3IPxBPdfh
AYSGf4kBurbA0vSJKY9pSbZ8tgWZcI7YEI8VMnyb5ovA+cTYCQbeedf+E1wsd1/GE74dliLVDQYc
rdqCXHshFsYlC0WhIz39MgAxvHWSz+9TNkVnjFRwzbXDHPSTs5hWmNHcLVI+vwaf9eDSfkKDbaar
iORABD3zcp2yYnmwcdCwfOzDvdorndAv/CHVdjKjJaFLRYQtimOACTwTdIaqP0BWsl3/2YbW4RJ7
tQ6dakJ6AoD8sGJCkngSRXu3feiQrOGBiTjsCcNy+UwWIiGSAEBuY9/1UWML+bdGom5mgzBuakeO
KuIr7ZjbR+yWhB/ZEhxUekeccTV08I/Nk2LRdW2QXzRhRkKHU/lyEx9Dio+B/7YF7epsJfElyQ1P
yCYlb6X1FHpjvD09S00928BtHtUrSUr1ot0MB9Ia13rP+M2+w30iZAy09OfiHvfV35toRcnKpK59
MV/CI17Km5UaTSPzsZrRCPCqop2cAK4GuMm0qb4fObjpbVGbI9UXsr4l70p6bVGbxteE383C+TNw
arYScslByGDufdA6CjSMfB1CkJsg1CDitxxnhud230m4OnuMryqlveqvHBIZ8uOp9eHWotJFGciA
0LwYb44lz+4sZ1H+7Ox/IVAW+BWWCrx+moEUvOHtkCH7BaDQg7Vd85cRRzFxY49qRslKhSn8LcCl
4CX1qvUYYmIIM61ABqRAXW4Xwg1aUqPxxfD7D4qzQlsx77+3ppW4air/uIkEy/tsbyAbRBs4ShFm
QeG1qdQ65Mnh4oQNTpt/QH0ClwGi3sbCb8J+x6dIsmCU+f0Zn68Bz3Rz9Ec/D1nnqfRtuumEzPkw
htMtbtNWRIU23e0HZJAluSmILRFuywKUJRkIQA2fr7cLCbAh4d48EoeQEyhIHpPPQNgJl8/lrRfq
ymtiKuilcPjLM0FH1czCJz19CquJX1+d3qOG1EVZ83UvxDIi3b/bO/ujXM14+Ib1vPIJAQ8b3tKn
MWF/SBokKtoJnEGcY0lh8Ca0HC/NTPCtYt6tKVkM/shaOkTaioJHBks7he4PXIe8QzWFT4/jrlRX
g6zy4lET/Q58kJjpzk2oXXZg50jf/emQfIMil+yhyEq5K9ph28rkRpwZn+rbjt9tuOLuAAXpcx6O
JeJtNLMGF2FifRV46vzsL7Tl5inznHD7GZYtXB27AXu91f/BwEQ2NxKYVjuNCOVtJFb/dDdCUJKn
AEwQeR2T9kE1DNXbTFkaXZajrs2BMcEj/JjdzN3Eoj2A9KTN9fWfbcoWwHwNzJcjkTn9TldkIqBC
3mV2YFM5MNa736McBmJzzA0yNK/WVu5JXqyrvujFIGMDY+y2ip3+sXi/5vj6dcBzAik+RXuS+mRn
EM/tNzsh14CFcseJXlnq1fQ+MUpfWnmzYkd4faFC0qsqWkh2Ot5kBYXIZNq+on2xRLxV/zDHYsBi
a372wCVZPJw7GM0yL9P5w0C89RNUUtpCz7wzrZT8fbZ/1VOl75K0zmJdWFt3Fk3BVhi2zaaBivUf
x3GIC3WV11+lVmIojtny1lOsnHvcN0vU5yGHoefvHsd0Tg5V1MoLuoE4tspTXvC9D/+YcoJTpU6o
WRqghQla8AMq7nfTP54SSAn+sSfAr/wXIY9JRLTNI6PLLm/t1lozJ9vhf2DsmBK3AwN/E8hbppKV
1u/BHl74P9bTnN9aVOaY0Sa6XhT55GmljtwGoz0sZCK9diPZMR2jmZEMRNBMvc6x/YRcJbGv+tYv
qRdveraOtXuaHd9evngTe2+KLGKsO79+O+98Xcda446z49fj+8nlQVMMLNReGUtbxUNRvRq+73Cn
uN+N819WgaIboealIJ1bBrn4ed3s99omdqSVou+hTAYaxAN3Mp/63l3F5WVlAxh9Y9uX1n4Rdfrm
5sD02/IuvWE6Bbwf5XKgMKP1HvVdOzYcM3upTym1ZpeAsi2gYYy80slA0dx740jMCwVC90FWiwtq
KP3ospy94UC4/9+px4cDdFzu8ZcO+1w/Db5vTyI2rArD0Df5JRN3aQWKP2jEDdeedvU108Aq7ukO
kYKmsA7K30Y4H3arH04aJCmSDl1FfThGQnaka9/LbCdCzvr0fEjKp5KUo/P+aneRdyLPsLqFnXe+
T72KOH9hzdVm1qEdQFbhM2zw5IOrOkvrouFlUW3oaXutjt+xIkIVRcDaIqiv7zQHrTWp4/PIlNiB
mvPEO79bBVuiQMkXxe8UmFJOmmmvWIMtyVVJuaMMMKIHiIErPlcXti15aP2P1AVqtKI664kq2gPr
1CJAxZo40JPQSh81F+y51ltlJudvqGvvoQmd5pR7dtlHospeCcB6FepxhABRj97RWGfTbyCgWyT5
IA189EHXjmq8yhDagzHgJJV+M9iEMFWo9ygCIu1C3DmRFSNwHSnhKDWI2/DvRB8zTKt8Ko70+xou
OPVw5Fm9PeSPev/Xjk+kJ6g41aB42iotMbBk3GU8whpKEE228NjvQd1INH1Mc9H1tBSu8ix7MfnU
ikZm+j7HClwBtZxwDyrpL8Fa7YJ5nAEVWV4K4MHck9OukqEl3iOhqL6h4aDvHmOfJfkyHBKuixtb
kM/o3NQA2Bcwr4Q0tpH8m4WNKXOe/mVbm4buNHaAVzoSoqkc7N5EHrWDV2Qj+cST9TU17229YtXY
dWFxUoxBAwH6kWJIht3xbikwiDgAWDUydnMFod7FxCY51QhcYcRU8m4MH6kmfHgCzKvBRIeQOarn
K8qQ3pMKLpYceCoxTYewnHDE5iBhkKQcIaepRe94PTZQmXmfvgy2ZTtGpP3uWrobL/tmQboSpGOQ
CsqRVenVli/YoYSAefvOpDqMX2beQM2lMms//lu/SGybxElBUDHhFHTletcY3QoZh9vP1s7QGju+
k2M6/czdkifxum/gGsIxzi9d94Lj8gG2Pv05oRZS9L8R8r20DfG4Ytx55EY3aYPW2MoqvzqK7z+L
KulOQtN2B58h7jD2iI5Xw3fIJmy0jcQ+zzhiJG/8pgFNbxIrJLRMOT6xEwJeur/6HTWSLordmvEZ
hD6nHMML68p4IItDalEMMGwuhe+ZWwvPc7c6aGgKr2VdqmmrnGN5LTtaRayfoTEI7uEG55h8oC0m
q9M4cBeDaSBLyL0qesLaaG/PP7CGlnpTpn3Gp0e6NqyurdxMgYNDeQuKS5eu4vF4bVWlefPh2YKT
EeeZTRZwxZYK1iUwWBAdZv3wMR3Z/iAURfLz1OxlH/oxuDTuagcs3kZU3cbOsryE/bmFhSoFJdv8
ZYriRLHxTqgPSBgh7WCcLZBnuJWdgB3aAOPBNs1h9rIamuj3I9myhTtNC4oXglKEHPlywHLz51Tx
J+LP+kkXkiADmzxI0ImDb/fEfPxnprOjLUxoUxzxbn3SYsjAncJ11E/hQSyRuyxgw6WQ6Kz3sEYu
tlO3HW4vEP8SH09B0CTaVWVhkP7ZkGDvmIz41KPh8MDaWpDQwSLyh9KlcwlVkhMtFKJD7Q3y02j7
gBhxeHs1/4w0XWR9Jb3HS6SDWB3ntZZRzT4IU7T/78h7MvsOsTcHJJ1jDKEyOcIkml7FFnXnjpzk
vlvhhEAy6LmowZ4xrlxSgk0BDuV0W/ANn1JzT5leAxEQ1XSzyBsE0OL7jRPqS2IR90SvfBLzBhZJ
gRFVDMuUFXPNIuQrPGNNKAxkNOYFFCUHUF7zcxcIBm9NZY5+NY4gjQ/OFYQahVnqu/ZX7Rb1sw0a
Tfn1NyW6HY5FeCxS+ymKXN2YIL6IDfkUY6vgh2Yg0GU3NQEoAFDInxRzRkzpFu19kfnZ8uVsbDlA
LOpSb6SHOoSxK+VHHTyDSc06/+IkBDw5bNHMzR+LwQpTIAj2QlE40IbYmyYaNxsGoiA3UMyzGM6E
qmTUQgw9s9Q3GN1ou3bGSG+iuw9fE0UIhRsbSpv/f5QXf+X2WXwDVrM5EWxSdLowIgHT+g/RUUS/
kBgrLw3Gt45vQloRwWi7g17qrqjRVKcGDrO6V1yD6gNZg6+9g/LgHfWu8yoN3vLKroRd+uWqqsme
CPusKKHIqIr5Unoh5ehMT82PQEynTQbRmV1t63P1WssfZhg/lDykUMu/MT4bywL9n2RV/DFomC42
UO8V7cHjsQku4BFLoXgJrsaz/WhgCrUIg2AMQJNDVEyOxzEYXoNVQjS5wxXdldU5gvcnJ4TChuLo
xKk6fsKUF17Fg2AF6YM0XlUSKrHMc3HR6b2ibo7CaiFTuEMAOoYZXWo4FsrVGCx1bYANt9bM6ocD
6gZSInwF31VxCnccvJol4bpg9e74ltBrWofpm1ad0zhA79YiaakbUE8Q5EnKhUU6SqfdSVc+IEmn
DbVV3XHhNRdwKt1YJGLWmX8JXKLHiBlD0vAc2YYf4lBMd+Lt57sj+ZJpfpoJZmMNJjSsKF2OcpXs
thrKmvauBAcGQnpgFtojUV8bevuEenCNGYUsnw1yUOko4U35eqzaFgqGkKo9VKCOqMZhvrxkj9ao
drUMxZaECCbqCLtZuW1XuWqJl39YaehMyttOqcJ8G0wx91e+bmFp66UzkW2uAIXfB2yTMyl2Fit/
XB7m6T76vC2ngMJ3eTEsclAQ2ARuC16moF+GCbHbaWII2UuJAm+UR8TvaVoh1bhjX2J+gkqV/7pY
dCACQi6oPWGGWuvvzgIkoq5vD2Erny/wcuNq7/hB4ZToabcSlcPYlUejlqO64X29mz9AsZanLiA8
YSDoQCAngrEBMK+IEoIABIUt9pYJ3A2NLzAUGAKqR6YKULiM1HJVrz7L4Nj/VMp3dRNqf44hNa9+
DABmoQ37g9je2cigcG6Oa2EkU4G2ouRX8ZX7WYWcLSYfZcAsm776sFdi2Iwsz+Zd4YiREdI0XI9t
Sl9A/J8mmMXFIKQfzNeK+N3/eTaYlgjzSfggMjme9eflJO1BfMZf2A3Pe8wVKxIR7ZyVbHyOaT6B
uoAIgY0jJVgtKgfmG32ItAr5TyVvo0x2p1Aa7bBwYKa3kVjBSAEptgTWjbInzJJtfT6/qyYgymzz
SNS0Z5S4iGcDHGl5NxPoHfpPF2ykC9Q2OHCqdM4yZqTV3dC6vb2rqypGXsR1gLkKSISEJoDEs+Oi
Yht3MoUz5jLk8W6Re/MdugoK5G21Joknd4WmPyOQyWbamOZatewEEfzvEb6pT+r8wC1zSaNSklok
L71rG7zk5ZEVEmo4Qbp8ZJ+Ptw5JZhGagztyf3YOVB2NMLu33RZli9ihm8XsqeZbQugZjueL5AtK
dhBdRUTGv+OeL30dXfWFFH6fI1MK4Yk4kVcApB6smBO6areYdLNrGprjpj8nFc83W9pNHveWoqjb
DUTMEwMWvHPXeGeJK1egVICRnWlX4oNobgjjVgZuTjC6sTmN+0Z90nJjErMmiUsQ4+TDwlM3vkYS
HxeGBt2WKcwQBX682mWmw+dSoc+Q/SBmwo1mpE3fOe4p0bQo3suRTiMHVb9E03u/Rd9B9NqMwLLX
oxkMV+ObViyoZyvwob018V95EL7IAVssmHbQrR0zC895rYjd8/QX5v/5tVbGe0linKj8kkvXpMqj
6R6LfJAQ2j3LtXy7pUtchkwUQBfWvGZSFyZp0f9B0xzNoYmI5/4YyVeAUKaaYHc3Ql/+1jgWf77h
SNxWbwQQCizPxQh189ldB9Th3+PB8s/J58zwVk/I89UYpP6mkKT6kgbzMCzUSFyhvhhcVYPNMgYw
SSGzARfJz7TMu/arA6errxwlBh3bQw32b+EaYvav2nOXe7VA/QL5ZBimNcKwppKdVaih99XJR/Fy
pcRj6AUGlA9VxIByug+aJFtWsTZNykJ1u0B6SugvzOJBFe+DzDIDXHV2kt1RO84ldt9e6EG0WTpq
e9U3d5XGUxohvL8FXEPi4t5+aK8RnGQrGbNIAi/RZTUDndomE/n0yR7jXAc8CcuT6rSzcB6e5mTn
jkNmxBONQCs/KNK7BksC2cuvTitGh18VvWZrHM/8x1q3nagKhGxrcDYXDzNbRqF8jo2aWYjo4828
l2J/zYvjjiWc8DvfnrvRyYpqqqhwd71UpzlrAAeBp/Xnc+3iFAgMTnGHLTiY6CPrVChe9rqivUE4
ILNzA9aOQom6JNK9IWfglimajF7zLURRJer5dFoDjmjOzesxY8Ho9TyUozAiIRQ+m/XXQEnEu44H
WLAtlESjAGAiOjtbcqOdePO4j+tug1aa4z/1r1DZ/Sii2kCLd+cqOT3xVZdynta11WUYQWm1erK/
WHUljYtXMr3djOq/I3UFgD9HeTV/4X2+JWEFhhpNTExfBwu64P1rqhSRTSBwHpA2c+FiLrfOGbQd
02TaNMDIxbQvb9osaQn9pQ9BuvLgURKioZ1TlzmGdo5r9ZV7zN/+egemmb17IjVt1OSol7R2JGc6
6lpCkDokc4yOZHN1VORucqwsocaubkJcFoZBgAqXNC/zYdywUlWtbltxhiLWpv1lr40jPAI/RycV
Ouxxzp7sjf59WvyD7EQSo5do8iVCCsfrxsU/jm9X+NufQx+z/kq1OD+o4ISpJqyb3USnR3TloFnm
wUulyXin4YFADddI69Q1qG+BREXmbKijAellM5iNB7Lfmx8txCbGeSjCyk0M8CgG3to93PbxdO/W
bWKHP6YMqGushZkXsRqv4x1Xqj+J9qcohHnaEK32QtCthxMjqA0oY3iOkrotV4HZSw2XffWebYsF
O68JTosXFQhG4gPxW9NRWnFwfuDuKn6wMte+olrd+EBuDEVt5wHdhGOZnSC0W8JPzRuVDaZU7La5
RH4zVmDTGQZIbqC+2ajR9BwuihUs/nvf3nX2Y8czCn+dGG8EVtINffoqvkfJb1jYr04L3+wCPfYO
9c5J/Mp5qfj4FxLBqQcEg4Muwc8YtgxxuKrvBvmSM26Gip+vwIo8x/UHYByxZ14Y/7ma5ayCQu6I
hryYKmww3EXFm7iVoquonZ7VLwqNAgeZ1+9ZhUlo+/dRK+nUnJmqYJWVk9tCdKyJUYGk9uy5PyeS
z7VQmyifKZFRuWwEKIrXRc/SV9DKpep7LH019QMFMqUivvIWf/UpBP+xJCjhtP04NMwb5V4GC5Nv
2jmf01xAnwYT6sENAL6+2GC5JA/xGKKaYBaii8SoQqvyKMoW3BHOvs9rbpHAKB+0YTut2W3u6+iw
Kpsnpl7XjBPQWy1yHq/GKS07puG7yzbT1D08YnYl1MRyYL3Tfr1+M9pV58b4PdCGdpZHVqAwDFeq
WP9BN7YADpKz0/YRkWtuPpLCUIsE60FZdh3p/hggA0se0YhhCHRBWTONobpSSJ8WqmDBjUHVdVYs
c4pxWoNVN1ZagwRSbybpBOKPuB+yXqhd2zWEdxkGkW5g6O46QVBEx+Nkt2sRo5Ak3+2Y4OasDtkJ
ObaanT+gsY2dF+KLVSSqgJ+eJ7pJ4vHPJD/bDYOTGKuH51ZEtPPLCYkAS8epSjz9WkO2hw8cV1vZ
4JO/JM8lHp4LdvhqiaFYTU8u9J7zumw5XXq64WDwJIzs05UgMFoBjWRSkgoEL6bLfGvTlOJm9Ycj
j4AEtNqe5oyx5nM8cU2tmMdaX7aOVHbAuzgnJtrLfM/MqNmQWcGNxtqnCqd00ZlPzbP4asSYBIjU
O4eOPuL+zDf0diDNs8ZXOqvs0Arf1Il5ot2fCC8jqtrfX7CntE5xKLyRbFjkKPBzUuIZfZsW8vbU
Mwm4mEy0U5jrPCzNyWtWK1QNjnlBCTOklF1Q+QHM3Q6YGmqi1gtQH+Vlw5UieTJon7ejmPE2+AhB
juQd3RLZB31pZHd4e1YCaN28MnvmLBG9qnCFqK3KJ8VAsMf1Ihc8EiWPR0NA6pVo+cSM99MrT/22
jkp1RoNjmpTG99QofEXpf7CtSCuT6mI7HGatCxJiEDXW1tSPeryKZHwgOLZMObeG6Fmz3JP0y6XE
OjkttBrHZZ/bOH9eyVves1sumKxmbAoBUhJ/BnR5rpaHXKUQ7A+1AwbR4W1Tv1mVP60ruf/SeZ1I
KF9yjuts1HGq6UqvwNJyQdHcKflZvYBxvW//wKXg5wbuJZ2s2OaSPjmIWM/F0Iep0EJZ6Vm4sYtp
CO9jiiXl/tI1mKaaAZtCwIp3ZHWNzD/KlCDmt3Jfl2kvS/vXjIssv+xqFVjgWZbKmbd5MuIpHGbL
tROFoE0OrnB1+93V9Jt/ympGWGJ9HAEZd+EDrEzZAGkp8M7NbLPT7pubjvzinfQAAGjY5ZML9ama
mgNA1XoIDFjUD8pRoRUSTkb+U/dHZZu8A3NAiem5dGWAOz4FgRz6rAzzOZSjnTwM8cYRdTkVTMvy
uWu/wIgDaXMo/BSPp9aNwWORI3QyedXGUCHivJjQq7X8L6Igf1A/syVL4Q71ve/dEEcwl2v0bHGV
ukpa2AH/uFoiIpLtWecVcrw7mJFlYoGX6GfM8jTXiLdf/IYGTpjPBiflvLitwDbMAoIEpjcgn+Z4
ARRjF0FG/XW5KwuJTn5PPsaE51j3HsEcEi9b0dBPS/4ENXiYS/Adr7W1Ami/88JsbiCcaBSYW4eA
nzvNM+lBC7Wa6t7fNdxQgvlWsW7j3w89mku89Fbm4yY9lxeQEOjrmomtOIcoWo/GEpIooUBhUlvM
fPBxjrSBq+sUegRqdYtPYszO4Z25lwmGS973LNAxPLalixZu4oC7Uc0jdOPtdh/tGCkgk/iLiYCz
0hoDWC/E/oVbqO9pRFauJ0ap0+NmhJzUznKKvRmwqqgar3++b1FGPeShKiDnK4XW8/7mYrCDbRac
D+FxZTeieVlzk5vtU2v25Osu5b7y0ygjViko9edIGtcs6zzlbkQwrMZS8mFLwS3m97d+WgD1g+mn
dApWy5ic/d0S5oHWU3eP//mRNNxWO+QFcQOaW1AIGwuSbwWLmmUEFmXv6HMipg+aTdt8FA/zU14C
FTrEoNzn+uqXF1iXClpXFu/E5HDV1LRyf8IcDz5Gr3WHLvS0wW+zW4BfLtlxajaMyt/Xrv6vR6pW
iD0GnHBuZ5WpDQjKO2auPRCQlCSeQYnUrN5sJDiY3CjbvdkebOjObET3RwJYJ6mDyrFcz06229UK
baVyEMlM/X5X6HAk6swIeCTwtlq040tv/EFhAxGgUDntjVOfDuQpJgXQXpA4b0Yxgrq8bTCwJ9E8
k+2XWlPQOLR/s0GM7w+NHuwhvIspNU+Izm2VUqYsFBBxIGPrEaCTBa70SsfZJjljyf13h+TwshyR
On9HktbHf8roqBXg33fKZne2v2sa7GEI2dd8PGELDRs7phKmMDJkxxBttlWl8ynYyZyAqMNSGvDv
j2gZ/LPBpSGyLuQQTSxw6QKRo628s5ggmiH6phQZjEpHN05e0RnHGsLP5CFzW7TJEuELqVmQRez/
b4T1O46ntZqaLvIDdrIxHQJSOveey//B3zHgAnv9z4cbVuCYpKriUQYkooEsb74Mhwtesfptb4hX
bp//RA6vh1fMD5NUBwT2Sc+jBCG2+yhqCA4nDAslzPdFLFYcXp96NZJhmpLUCY6L7DlR4J+Qf8/4
o1zl8MekA5PNdQ9VmqUf5IM0n8br1HsnKaUyq9pXhA9+7vcfEEh3FYcAMWtomAFrB298XuVfLbbs
tOydPPHEH4Qkf3OzUoH2F5NY9bbd2yiYBh8LQSu2m6dPNimHwfSgaPCjFYy26mVBIPWqHinUXYxs
dN2rLpH53haRtVN6XHU3VSnQ82K2YKIwOs4zuns4ypVqhuScphullinvIXPpX1roKgE4Zqo4eTvm
vPMZnoboFqvNnZvxxZhIVFfaAlRIosK2Yq+U2r9cBVvm6CQCIeykK1VkE3MAHYdMO1ktQHvuv4xB
WVpXLSv1Gg/WmuNjdzTxr8P1ZgVsLBZpbWeGpwZUlNz0PFeLHUek1Nr1ABEB1hHa/f5c3vHTHyPv
gXrJEBjmpYT2o9Yxy81YBUNAke8L5J1U0G5u9DLuMHZNxN5kyI9n52dPvmbbQxvkmLjPpLWbnrbC
JqGjsxf/ERbbK96c/I7YRYBSQmKcNR5/850V3kbaHPm4CrY1NPBHlnUVJTxijUQPrSvzdaVehKKz
6KiCVIjmPloV1Sfu+jdxPIRsP89vtfwxk/TzU3Yz6dJjPQyi4X3A8e0j9EAkvE5hoGDATCocC0pf
xZ83wlNNhsjFYxqBZPvwIQji6gJEDceEeEg/pqPwpk3gCPQ8p2P2pB49SH0B/3xV4y73bEc86aCu
w1UAp00dhcYxLfzgOJk7Qc9+Xr0hEEtoBPGk+Akmn4eQ8dR/H0bbcKBtpROoET/RNLm5GKb2rNhl
L8rdxYq6tf4GKoQoLmBxJZNokIpvuKrEvOeqgah48S5F+njfeh1IbyvZ/UmebSzwlkVDJhQBAT0/
3UozAMQiRRYmeaoCVlxpr6z4c9N3QHoD/4qN+axj/XtxR9kNJjs41WHwLJfjwY9TcnvqTO7iipa+
2eFzMU02aoElOXCZ0DKnkDM7FRwTkuoucSE+wdC1aQGaEq2LbLzIGsB3lVKkexo/jk+RCxJ83ogE
wQn+wQV7IPv6BFYZaOx/pjZl4w25v1TF23yt1fN/AK2t2qWQW8WunirLxnF3I2Zofbqr9FK63d2i
tLmQUzjhvaOjUUdMaC5HmdPggv7DdssErxNHurB7dMMsU9sz9O8hJE87jlZuhflV61z9gCHlc0mS
ZvZYA/mU5oQi2v52e3e6wGRQTQAkazXoEKCT7s83UMTvY2iB46aeFo5eAjjf3jxifGmjZmoHkOf5
gXLCzfieRkYDnvSoZmmcYx28B+VZ8DP7bOZeDrDVFqI0k+D4vcYRK2/k35/oFv46rLmeD55vX+5x
NvwH34SBk/HWsM+kgc4RQilTH3vKU5SbY2Cju6eSA2H92xe4eCR4rmA1qbJqnLplutXvfzIBCdCX
6AFwEBV388Ulja1rLm34IEFPTOX1Ji0m+RU/exlbBa7CUMBYhQ/6VWECcvJVmQEjwY8K9zS4zYcw
KC8zefX6DJCuQ0mMJecD1pokA5Y9mbacDwi6PANjWXTCHa4O9Th+EJ2XWfD7VfmP3ucDur3EvMPp
EgWy1mFq5u+dgXEEdaOrsVKdI1C/ituMnFvu7/5M8xjOi0XTMC2c62+eJRbgQnE9n16pn251MC4N
NCQMe/79FHjnMdYWODgdy4Uan3Kw+JOoRJCJsV/5AZZyO5heBDAoKZRBr2zYwGjyjPHJf9QXHr0i
oUjYxC/qRhsWqaAoCwTw2GDOSRMJuvGdlnLAUFAfQ03NFAoqcm5jOAQyD6cOm4vN3IaqdND6fXTV
5DPHyDcuYm9n28PYULsZ8tRMHvmnNiVBasDJm/xnOO/fa3nr0KZukg1UM6XxuaIUS5zcy9f3lq60
1w0vVcqa8t/6MmWd64MB56wyXH4aQmBM6LsQULUCX+QkYoHRUNCu1wdQ7lOrVN2xMhLyLqdI/n1T
g+dBeDJ0oozbj+72skX15WuGIqX8R7x+1/zdJogzR1hpyBqFcHAvb8nxR5vmQLwLA4DaBTZHUS3+
WEFfVoBNbzjGYbnzyRgQuC/Eo9hK1+d4SvGD8QWeC7SPWPoo4o2BQUpGsSGvMnRPHrXZmNa2GjRV
YZLOeXOv/shauwxc0ry8UDDIIeMvgi0ZNc+hD5u29MrGYDyieyd5qSUH36SlBTEkM02X677HNkgt
lic9nvoKrT9Y0nsF1UDHN0Z74T64UAdATtnf6plDp0DmMuCj0t8S+J9ia8+0kloXNDL5Bp4mPptr
XZo8VSq1X2xN8JKAGfX5m24tKl9HxBOfO8K+iITC/Dwh20rqyNRC55n+vc4QcT9HsnfU8Z0U3c8x
uCrQQ7fjMGpHO6G986Jt+ZopBH+ktACtR1dKFEMA8NFoFXoB2aSZ98Sp7C8DNn5FsgbpbS2qkXtl
35SxCGo4dnY4JbVpcnXrhVga6N2zbBbrWsgWATWxJjvs9Kh7SOFNpRn0ML8RQIEphXemOEH1GlSL
riA5fuOm5QZ3jR6Qjdu+PK6dAstYjFSkjNJVz1Ypphz8Wwizwkp55hrgJ3aMYjVbVp2NhqoEHQFO
75yhbUG/DpRQQ8rM9SGQNiMp1lLahxlomfF/6ZyltHZayKx7q/5fQnaanypKD4gzkHcmqqJFqj9E
EZmKw8HEFwa5SRykXPdJkr4Iq872r+Ddxkf/K7FRMZwaNeeF/XeSoUzRhr/pzzpeJxxilfsmIjDo
OsFT2pAsoeD7A8ucQCxL+naM7Y25YqwDmINnCq4lDwiLz3GCN96KC0taO0BbWG/5zqh0g/Prku9r
zB/b+ZFRxz3Zt2H2y4JvnKM4hVwAX4SqmmIYa1EP87Hw5qy9cu9v2Il10FeehT2EavYU1cgdELdx
FgaxNE+ejx96JM/uyeY7g5IMqHvwtT9Ssko1RV/wUaW6BzZUP9Tr0op6Tpr+8pQaVfnjGoEu077p
RhD5mK9jkyNqT15Zw7hs6jJK1kEvUPNFwgnsDLUUXo+y8zl0Es/p3wDKKGIkPEKhWAbIYMNsU5eZ
MCca0lOW/a0xklN+q9Qv4db0KR6dUnl84ONgfQc1t3UQ/9iUmEFsdMYHdHWJFCrjWAd98hDFhLcA
yuAL8yzS+m1aUFp9Lc+pOlppWVjUYBLzn6flhtYjJwuRy4dVBdW61aKPvvnhPuZndHJFnNkMTPCe
VHh4EPT4fVS7nqcX0PUI0XTYh9iEAzoIRhBfpqTUIp6Lo4hosek9NwofgquK9kulctMxj83PFw6L
dTER/JPUuPjJLi/Diz6DliqRpJaxR2xPjN30FDvAiV9eGBpZR0lnxn3PReOofzOB7AQUDRkYR49p
grWjJbzoDXGkTet+mI+K0RpIcSvs6bViyf579eiDed37ZoLYwKiOnivxGbaFCRwodgTO8TypPspJ
3C9mAVmn6rbniPgwRFyZ7/5+eM/TMmbRg9PAS/6Wf9iFmXvJFwmwD6fCxqkIKjX5L1NjqABKCJUp
Sb90Qd+uDpRPCto1d2AGGpI2RtddWimMVSCZxy+aJKxXB6nXKEDu9Of3Q5c7VubJUpkRvG4JJ4u5
4Jv+KdU/Ca8Tg6mP/l7jdlAzO/oTLGBfkM3h+/xTbEGClC2k20BC5JyxNXLAH783tkaMV70LRvyr
wVBVd+Zex3Lqvn3gXMZgErXgl0EXoOaT7xIr0sUv8Ui98UpGNab2m0J4pO2bF8CiMUhy5JpFtlpL
eL6KLS1QDAtYa7lPtQv2iUjUyUxs1oGmy95jl9AqbAa+brfm/aWnhNK72EDEJHSTMWvvy2I2LFSs
/muyLYcVSD0Gspu99s9fxRqlwpNOFPbEujP4C6P571GRWcuhNLpfuT8wE7u0X9yhua5pf3iuyCs9
gHJVtngez01OCYBYCOT44l/6icx3/gbic8OlHhn3ADcC5nKKio6fDrKDxvWMfejY2RimBre77j8V
13sQGhTgSeiZ1v93C2/50cgrEtf/Zbi5wCIS3iG4uoTHOtNfz0YKkTP1vRdf7Co9WMYFFvvf5Qf1
3kretoFGRr3wSlq4godtAqqxNpQnT7vUHWb9EtgX5ZfHXCbhS2iwj0TOPZH8EG56yz++8XJC1KUD
F9yq/47i3WDJu2hssJpgZha2fm3ZbXgEaY5+GvhWw0VbG800DCTGMffH7h2B7XKX704k3xPJL8Xa
MmbbV2/wsoDzDyI2DOEOHa0k1hFM8yD2ylCHCJrt+ngBqIdRiY5HyPtrbO74/6pUbYSrNZdGHBKP
Tf2RIa7rPmHHnhO2jC5sDECeZfCNg/c/PdI87rRmG9dzlhMsQ80nBOKNB1NkrPWAkVtXaey+nFU2
MOwVniWHF2ECKrAl0VI0ttveCu8mKaCJBbHJDONsrtiZigb+QrAyx6HCIS/LfpiB0oPKzjkj4YJ3
IDuAx6dzknq1q5bZnKo1XwCCpFtirlkIBuVYTvaBmvqBnTpzQNhu0IvBjrtgvESRm2jta+A7x6iD
Htu63JeTDN94/ou3YN4VOSLxyKnnp4X2ODB6v300QXZ9eJlv7SGSR45sVHr+nbbZ4yRszhGaf4+5
1yojiVwPjP4qICajfIX5H2nW21En0ybVbanag7QT0lnZ0TaS+pSIqOlosbwdAoHLA+oMqeHNhaH+
XDXtkXDowX8Yt45bZG60FWTQ5isjBBK8C5UI9RZYWcVizOgnpQ1nI2GHSmL9kjUK+SeAElUd5eNa
vxOwUy9aI9yll/NXVtT9YB1u0zIdDiWa8wzQLrYy/zjZYh/pfdykBxUoYoHJoQBXVfl1zotiTzoZ
59MMExGpYWcVNv6b5/R/B0JOGKih+ro6EXYXuIX7Kv1Af0AyhZiVQpOUDtW3uaoFN1NqcV7ThbXE
8DV6qELOtV3BxzQOS3e0pi8nzi64P8JBEpHxCtbnd61p8SGaTaQMfDKizHKISsgGJcr4TeyFl4tr
Pk9Nno4dXsrxhGnsnOt3Kv9DePbV6TMlgmNp3OS0WYLFc4O43wruWQGVzz4IPf/iXq3JvasZKUKv
r7Vfk4VyI5gj/wdt+WHVI1rz+p9iTKwDaucjblrJ43L4adfkbolBcntRCapySYnmep0lG+oIc6Mi
PVx1eBHuR0CUF1I0FYu1CPFzJGkAJHMMU8vJBy2/d50GH6hWMynVgvpAVz+3QVlox8Lyba9hhbMJ
KfXtDI+kuk0Ju3Er4WD9DrrQYQU8GuhgPMAdxkRPTBzi9gJ5Yi0g/SVptolroeg8lGxsVB8P9JHX
I4pOgglhfhfH1YPnRHteI3n84XQkwrrBPhNGStbZLvgu4rhdSF7qy8PKs2hYmKusApQM62+WA9sN
LOmwco5vTpPjCLDhGk1IbUtTZf/dKyV2ridkbmcRWl+zI6NuSDPqqFNBCa4S0pnt5ijoix2Z1D84
RilpFCuP/xbPyfbzyVCzPEibNdMwAt1AHoH7YV61kYShwDit/xFhrc1PGPCnCaAWV+TatW2vXSCl
992VvViqNSw29IG7LhaCoQttlNMMRJmVleXaMZ8h5DId52+4zJBWoSj1W75IGE2ihqWfg9W4rHJ5
yra1zz0U+n80IXQ0En67aRe8ljy5HzCtLYR0hJ7KokX+rdgbt7Vn+4KdcTn/vP4ZP6ABaC3XSESl
q6Ke3/pw4KaJYdaXgWOOo5Bh3LFjLgMVyeLi1Gyz+XTaPYB5vq6jf1F+pP1X/um+lRH0ZKmlhvAw
Z/X7/NloJAK3xQ+c99Nh0qhgHJFxAes199yC8qlXmwVf8lumTOx8RJhOAYSONB2VjLMylz6hKN0w
zqzMPTah+/n529T+GZB2tIrz+lAmw5II+J/wizZwEam3pGP6M4nj5HWwH9VkSWwCA4CRGhDgbS4I
Y5VZ6518D9DYxm9sn9H4BJLYidNDa8JjT6uDk0BeJFaeQv4PRwuozaB2iRDNZ7puR5FuVHsryUDp
pZ2wO4sNwnfhfxRrM8sXNvGzIh+jA1DeFFVBS8Dx7TbGbFJqgpccnHqEVDlbersz0cWPf81gHxyG
OnebgNnS2pZrE8riyND/SOkgv3StQVgpqi2RiaCHgLPAlrBSUlhoOl6JaLuZGJMBoibc+F5PqOc5
DLVOWjHKkv+ETcKB0+uYwFjHD+EI6N703J4taxCI3m2Jh31Zso5NONnTQMWTx498Kq6Qz5Tsnpl7
kMOAJv/YXha9TPTvlKiQ9GxaByyKt8CRAHy/zH4HqoEzvnmNvLvxdMLDkX1EHTK7NUg16m9ETijp
5NFHxD9mFHvZGh2iDHMfJ9E3tZGTap3JHcwurWgonwYiG8MlcX5ZMEfF4RII8olrgrxLGsvAB47d
AWzVVFq0q3lEXc5u6XIknwQtaK4DsuELZt1jAleVure6e1Cx4iTKda/babnxMspyUvcS/SQHUJTV
p1iDIzjeq22zzbaRVmY7p/xqjaARpdAhnF0FmkldNcx1ouh8t1qwTBJL9COvUlxwMfWnkWWfzyUk
VOXMtSum40cFWIzS1kYGqKoRmGyORtUjzDZImd7rAE/S2pBm/JZIMKmCi8s2MmRWuxMqtZAEcoy3
P63oMkMZsEdwAZ4QkjwnF7/6m6eqt/DO9oCkRtio5qGikwl0j8LJeKfREQBk54VSdka62iUXRLbv
ei+xdhPW0zcLL/Z/PRmHJ02J2aE2WvSZrHMPaib8pW8QTFKEaf5zEgew4rva0Yu7sB0bJRYXh1k3
BSParH5rCkCHQDSHatgnGOFr/tDZm1bEE3AkkYl6W1l9Npe3fIi6cDB2d1c+mcpBDRkb3uq/HXsn
wp9qJ9FFCewnRd8wp8s6W323t0RHWv6rQdc5Jq4mg0H1EYlNvHzhrQnLvprPVCLcQAE9ugj0iZyN
WrBQVA+MIgCfy6t046zE6331O0Qk7rqPycT6MPuoKCH3SX6HBNdZENATSRqys1J0AYFHZB4vJrku
Kjaoi91TZZkALhyxw+pd8h5pNnzneGhffYFms0fkF0BYCMnyQTBkCIendCr+kxJhHAXfWPkFcF5V
gU+QaPZn2C265nCjWGU+iC6BVYKc/r5VtyvcpWquBpAVpRGCswf1UFce6pknfZ2wznQUGKPpMiT0
3PnDaYuQGbHdVw4eL0AGq5UAxvvI2jl1XkK3MB31TFLnKEfBKRzzQym1q3g/j6yF6f+MFFSK1mwM
cFQzfWvZSN3ficz/i+MHG5v+PdWqoNFRYDs30w9PMft/meSp5h+W6r7lOeMvtRVlxUqgLfS6vpGM
PsybSjoVPF6Wev2Wb7Acq4HQDztCoA+TkKNWiK1vdd3BVKxAuk5xQWA0IWeKUNbJefYXdKV4L9Nt
Nimlkr9TCiVSkMg31vjs/huQdxBXL36QW+FHhODqyrq4C+WWUE3I5Z9MZftzR/bXcsXpx3GE/xNT
Pw9VEZUOIvH5w5k/RQobScAKGyz8vLlrlgH4+pBWybTuJ86XdMEvic4CBRVdu8H9giG8pwk6CIZn
DAzG/7o+s0tDCYCA41/OlHnBPeN4+j4VH7mYS57cGihgEVTiIh89H1BkSLjmxbUIUTZzKBCGYfvZ
h6eagIgxSjBQVAH0TzgokP/v4wl8nBdPDvutqiD7HT6bkfmD4O5yXm/1JF1Ta2sVRisYdULum11W
YctdkGrFleJ0hvLoX4NiEYkdLCegYvQN1ad9GS3O2uzOZXUt1WGhiQeEzkWKSL2+OQxl2BarUL3s
oESxssqqs+xXr9oQY9+Ca6qFA9JKBEJXAUXOVC1jZk14/WFZ4bwDJ9Q755qlJXeD+gdrK5eXQSQX
7L+tXRuia/y75qllxedV0A68q6Tb0BScCLwg6lEoL6I6hM2y5As++rT6kylMafCEDSS04XBLuf8y
2vzM2J9bV3fuVn8nxFQeyQJpSvUUKlcSqfIwLgjLGIqSkdwTBsMVwUdeOqtZYjJebU0pxhNfJdvY
i2Sq2M8Z6Hwa8X618wfLwcmAwHvQrrlM1lXryYXEb0rF8YdZs+pXnxtN0c7OVgRldAvP7bwsSUav
+QmuTM+UMqr8GzFSEzTnwfZJLgzVxVcWCUiWCvWt8sNEJGqwhzsCuprJ1/tWGLwPUa+r2WnoBBow
tez7xuF+eRFA7QxxUvyK/+4sQ8C0jquPSNtOmfHh2rhLa0awUEXa7uGFN+fim8DEq7Eie3VJhNT8
HI45vDM/a6bBwS7i8wHPClgKX2Se22G3yPjdmblgndJHrv3mpkhZfb/G6FMwLjIEezSjMjtCX2Dt
BxqzxUHxK5Gs7/xXe7+6KhzsA3sK4PZPuXD7UOjgZyz4umYVhGA7BnSrfzmLYKQOQ0or+5MVu8g7
MTl+bMAquBOhCSGY/9ORfNNo2sxSEFyvRqFN+Z9dTLu/mN5gNxapXiTb0znaWtzoO8Sh+BgRkhws
ySPgr0vcgltZVMT2A62BpUiUOLLKE7696SlIsIRIa1+E/tktX96U0bi452DC+aIqy0lKEoUQDQas
JMldW7aBWEzO9/FhZxz4PCN//cvpzSzCJeczyVT86xv8z3jaxAFtwUrhoa4pXEMS0/mkjCo5GrAn
Rb6d2bCQ6YDOAsILbb9guRZX/dMAzGyTAv1xp5D56I6G1at6HCcW06XWB4BqMoZU4NSjHgE0kuWE
K39vMOG4YPXxQOspANyTkOKVRDfgnyg6Plo4QJLTHY0KA4QRsHYZWn9cSA6ukH1QOtWSc3prbGfz
n6MlC1dr/77ulSZFs4SissSN9lASxH6oAJ6zkmcOwetXWmZyDhUgqYRzJ/6SfEfbheYg9sg2GaAi
GvDtrbamT32f/iUQJMqOLQlo4e3IIftfbCTuHrE673CSu7engdScL/p0zdhgYlTE9ghKSEhrmL6n
u8MWMYa+iA7gnnLZDVOxOH6RaMc4pbVan/qqVWVXXu8TCWhengIev7Y4LFvp1QGmUThW7Au8UG01
g4E3uH2UPcbPO56tcrXo3STJjvmtywS5YrAI9wZ9mkfz3Qz9b2CQtZKzhv2e/Dj/27tFf713tjcz
YgAVxWT1GJRLIAG4ttU0I+cVTN1eKh3DAiPzDM+R4yR9vnL4l32MKexgj6CQGhzbIS5h36ETQ5zr
fbMrGEk/8jkDMokhDyZekqhjdLwyAne1p5KlNlFJZMg6NOZb7BJ0yVov/stzYy+VdOrKhiG7z60L
nJnBnkQHOHJBAqFBDcR8p3I+k28B3u3uvDaIX2gkbP5/NKLaXlwm8wFGcP99IjcsosZBkzT+7Og/
N5QM1XT+bY4oJZPHNIXBhuB+wxdhmZqDgqlSF/vqvmH4O3iJwVziqCos4SZQUZc16VQpI3SAgJ+P
Rgx846fDpURjeEU1A00Eskw/VBWOfYwfZvjbCLtKBZZqfNyjuiyZYtmgoMFNSzeKhZ1PMfXnpTtJ
c/FK1SfmVU2HtRXSC+VOhx4v0f4m5Ec9i0+lBRex4LT6VSE+AVlzXXPoQI291sE3eC2vGcC7e6iv
lU/dKHbYhLQnTH3AbQwGUK73tkyg1h5OgVSVG8qIFUszsN/lMXMpIOsvDnidGx7Sd6EpJik4mh/N
h6F5TTo1DFohN3bSVlfYgdR2j9BhIqz1XxMF4tqIreNvSjxAQWdc3J7DZHqfLh/UEjtwWB042TB8
Fu7C6nHwYaY2y1d1jIPpkZgG2H9TvVAM+cplPMYuuQStgU119lr3GGEjWE7iodFDYKdbTZd3lgkz
IhxvHS7kh+/1fEWCEOwOYvgAvn5KoruXQBwd+PbT1j+2ytP7ROFeW2dQkvgyuLAJ6nLJKhG+XmVI
IbEIYKRuQ7sB1NyvsXBlyUBqxHPV84cWJifHKyK376PiPSaF8LjJHt4n+iC5+7iMlz7dWJkLUVGq
ejcajFMkpR7UTnPAWVmv71o3aCX1a0ILJKkQLRAtzwdNmzGENTH9sAdVV0hRyF6xw4DeIYKBER7w
l9BOVc/rQLGwyY7ph98TGSy9HVWbGvsORj5arC7j0pZb62prxzXC9/lUJ9FvvceU6wWYiXhtVUDB
dhjE4vJx8/PSNusQJrVg2D+VveOHeCjaCpLWYWETFd3W/KiUwmqJaFPB0Z/9+/Ol2KU9t9kWBNvY
zsWbt3V5S5ZPRic3UkY5sYQnUczQx9DIXqK4VC0hRgKa1EeDUJEq3xiSpYVyPMNL8THhhF73/RVA
GKMblzb8nJeKQfZIPph9+gNVE0KEUjbYE85TcLPrl71cOXfj1fgbF+TrC/hxVlLZkD0ummsG4Ldo
N0dBSnpdbAy2Igt0n/sJaJfS3wUQRVjNcZxA8wdAwNE/SEGJUOwRF03c6saUPzr5iTXWbBbqby06
7nJlcmxS9pFIkswb3l1VWMT0wP9+1JwCD3UDUXI3MjNzW/ib4U3SmJ4vTxeQivgFlXW9witnKBLp
CztV6RSlpzI//EzIk94Gv3x6P11p6lyi6GJvU8u9nJ3G9AGiC4lgqvaUf1GQ2YZH8cvPUtUWu6V8
B3QeAll4/GFA+hz51tntMmIYh+bdSNgLwZXc/eLT25awDma7T//QmJa6InFRF7QT8KEGA/GJ5XPK
0OoLiUALEEM6EA021IaJG3OqfAoahv+jsv8zyALb1+KNfLM1pKe+C17wUN//dIZHpQREw6P0HYIG
QbetsTNsTloqgGYh9n75ADP4b21YNTnRujWrCSwLrTgu/+Y4y61AYrBY6sIiYqsr+onW1WCSD4YZ
lWIVa5jEKWgpxY9FD8a2WPDJDM44AGyvMwY9Ca36u1VS/IMlSgXS55B2XdNyG/j6ODIM6aW9LkTl
Sk73GT8YVwseLX91hsCnLMEfcfbPTWa1NsBLmt6O8ZuMDLjVOa+0lWJSsgGKCI0ydC+6Bv5/cXGY
7iWrkHerYC0pc/1FbkkK7iRIGCeIugpmY24m3EP9rCcAQLTkJydCxL0mhDv0jV6ZCJCQF6AnyipS
q88zW6P38k/qPOw+IjxEjtu+Fa/rb8fjFIvi8Jklz2xAqFKw8jMSeTYHuOeDSZ7dLvLKyVlRTrUB
ezweUBGgvr6xEMTm1u/CbNUaSbHOUU3g0nfO3umU0tXAL7rS4nmpkE6qk8odf/6Jn4Dl1FhJ9+bm
y3auV7+TdaSTttvclnUi5ysbCTGDDF21ouX/Nab7iS1za4WkTg99h/nrpTwwBGIbQozvi1huXgeQ
odKYjmMDRCMexWG27+VHaqnW9zirlGupNdOICJNa8+dg4mdRhFhJwI/A91AKNqNydNeLZE8FXq65
Rd3QYripX06ZDxNf4A3m6UTA6LPTnnigm9iHfyI8GldwKvIFiKZESG5Nx2sTjZsg39WSXVp7glE2
pwlANm58r90u1EHnyclDCcZreKD7SUttZ69kcFf3Q+57V7uwxwV//RGNgx1L6oJk+aiMbm3TTNl3
vGsUgRVUkgUd+ELJxDPvsj67ESIAgZ/jpUtDo4iz1K1m3F29aSh6HMqyBtGzw7NtmKXylA7l1uSf
jBR67ZqPPRdPOp9EBgDj0ZTpNYJaWYSuykGBmGDP/OlBdghlvxzIDcIwvaPmVyyHwL8WCYPFlqP1
UiQkk+vDQYtZWZNvHziODFmSSQxbCc3Fhkm93fINGtbniEA5+/vLqJ+Mxv/Qrj8sSDP+VeX1wLGD
UNXOc3dRVj6mvhs/cogZbBd4p/hL9rjmUJ8OSGtW9SPh6qpNzzsv18py8bT3Idnvc4SCl+/lz4Xs
wl7DXgfRixvNTIMJeWaw1EHAKMcFP48tStIN0+aXsK5o1JuwYyQLhy2HzV7po5qUzhs8v4jN8Pfv
oz+ZW4+zhifr3RGxOpTfkF9cOrJym7cevUFtjhMY9R6LXXhRdU4opmwEIIa1Is+RDQOj4Kep63V8
q1IchZx2p58LCvlAx7t/iM3/Y05F4845O7jEGz/uOTxzHHiZdKr+MAynUQD+cjRF+zN1/GRkiG2Z
YGzNOkxixY2hNpOwem4Wec89ki1Lzk/3VsQxb0vy9FrsUNqWf7fH1xviyHaPyuX/hJVHmkDkjSZv
mnlPjAjuR0JN1AQNpcFdmBraJ1EBkr/NtZa6J15sRZz54rAXqkfz7S74w04ZFXvMfia0OIvarAzR
NXLk3dqkXwdBU3TdcosYRwlPeuHXe8ar4x+PAJe2pfuqozE72wISfNkDqLebk8TClUhZdBoYk2Uy
wVgVEmBAFxlP8ISIK8OFJeXjq0sVK5SUDj5w30Htqsq8xouIp+KjjPnia64cquXDhF5TeGLLG9XA
gVHKuI5q5+AY/RiIKX+w/tafhmzQMHa6wpMDyt27J6XlRbF9NH9T/xlSaNWuTbpy1j63ltWoMd/G
plorJQOT9/TpzM6Pqmj/nWyhJ7Ap5ac7B7RUzrrNJQqlBBwwSnhT6PQn7reqd+eyw414398cD8U8
ZKMPY9ZZ4DlOPhRohXQGjIAyoLkBFt0NROz69DFrWc1bLxZBNjDuq7JhDPGQyf+NE+s4AcetiOX2
Lu2BGIj/MSEq+j5EMEejgwjUNkpTur9UEM89Ib58FCJ/qgMn6GtYvempahBsx0PVBu1lUJml9P1l
GVdXHkBkeBU6uOGiPaVv7v7wnH71rS0TJrxk24lse8JFPEAED3vRFRyGlcoY0HvvwHtuQPRIIG9S
j06mzu1AAAjRrJLUDDMGGpe7cMg9C9FovOeyKpc77bF/psPjYsrRXnm2OC/UKOdYf0rgL9qAd4x9
kaTomkQJwIcpR74qiBI2TZD1eH51dEreF8iDF8/YrKL+bEcW4oPE6ZRQELa+Bi6Sq6dFR04ALVDV
ax43HcLgr8RzJdZyxyVNKs306AkbPa2W5J8BvLr+oNWFhjI9L0++0nBtkZ2SRqf9tcMGtozMF8q6
afmpmR+JvbYVQvYJmlm/XqVpQY2v4qgqhkWv+6H+Mh1GdpV7B81DkeAgDMiBLI/+CrS1bf9Hxvya
klqrNsuxbGqdP6dHaflOVUDDZE7YgNeSbqoaBFmzODmQkG13DLZiiHUcpS/YPGnoDhWNljH0FS8l
M/dYp018rQJj0gwqDKB2F9aIap/gr2ZAXE2LOgjIV4uRDo8XNgPrm14NC4LH+GpX9CpCgTZ2wR/s
/Aua194wwUcEjQuc51sLq7iATaBYRsd0gMrjF73oS3dPGvqwsXTj6S8OmX9TQcV8x0jJQV0mKldC
juojXD2ix++0lB6u93bm67B5KOtzMxOn/7IzWflwmGwlQcMUMg7i3DLk3WD5pNm9ai6uzs4y9Pmf
pkFcuW1MXMXpQTogUGTZo1SK92AYA6E+tgYkJwbTSaNIIgH1hsSOQ/QmoVR2HrHvKI8wszsozxR/
atF3w72eFnS/M7i4JDwD3S/G0gFckwaMrWaJ1iP+pm5pdtq8lDyf0wMlHWOZbx1IiAysR45vuBNY
0Ooubo2Vh95J3LiIpGznz8KGpIosCW+nTfGYqYCh3M2MocR5zq6UoXvUysumzB4QQUMnWQjMbuq2
LkTIIi3xCWMgdkgoY66CiRz9z3ko9dY+VB+yeDWDb8QAJfH9KGxrWKikAtn0fjC/QRSC6L3KAA1E
m5yubUVN7YEXq0l5PjKJTL9Q+LUCa/Kh3BCo/JV9PhF0iNUYILCGWVwpYHc89cbWyqYUxh6/7XIZ
e7iCgSJdSrR42/GPMqziYbW4C5T0I/PjHOxX0ZqxSaojZd6J2QH/zhMCGPAm+iKpivDLdkLRrV/d
n1SGt48yI1w1ypzOKqcZar6Ke2fpDuGiN56QoXak5LNmbvlaJLcQI0miY2yOyx5lMTXzFllZKgtl
0fS40vBlWfqI744P9ho1V1l6tqdAg+/OQESFX4Dt+BiZ1bClM3Z3vVIYggJvAuJe3GapqlHuK9w/
aDKOdBDavDu7d476sNjnfir+HLi98JEJOjtHkXCi/7kX1MAre2X4eC/CfQx/H6weeVP8aYLh2SGp
lnhGLmTfaNVB9GHS9vfaceR0JE5JcIiCVR0Vr5uO1soeuuySEzbr2HC96PuERqSBuM2Wx5ra2EBG
UV8AVMpCdbFV5aSoV6Gd+eOaITM6Q+eXtgeu7cuuYI6i5ZEOK+EXtMOty69gM6VwoJaS7/ZVzzIo
lb1wuy4+TbWIQy0qSxiyvPDBYqM32TdFO20CJgqTsd1O9rWzP8gS+49iSUgFuryzxzT8EIRwxT5R
X/uZkIheRUs8xxZDlMxRerNEE0u+tJoLOaQdzJZ/a+dW8q9WL/vmDd/JHPgfGI5+stEzF/HKn8O5
pz8ctW7HqeFTHp4HhklaQUUzOUqDG5jYCGH7ggZKo4egj8+idhEstJCwnaHQRdQNNR9LiVqDp3yd
vNr/8SWKRVqtNUpzOrG+YLYxZ1LPQ+8lKd+TxvU+8cvWQ5E5PVuCPv0PYrrefiuj+tMvR2PPJ/3a
RJPzyXxszRUb0VWhgcV+7qwdziI8Su0FXjy0pVio9FArD+Ee+rSP3UPEc2c9Tc/2PXjedlUCUY+X
2kpCS7szj1afR+TSNcDT0Xu4wxxbRPtriEfrEmnjyiJ+wb/o52tIk7JXRJXdv9pDw3munFVYVjSF
wOPOulqSkj/lk786+RDX4DJcSDG9qVo6rrYxgZCVvMSD+vvQCAOFynXk4D7PEbbiFTFHGo6MLnTu
ddx/L32I2ocs1Dg82qd2RAYDiuzwyBKdGZdhccFa65m2PVf2icKc+uuq+IAzwpY95m3SFrKKaEW4
rE+nfqXEg+RXXgo9M5n2xp+tpqFjy825h4V8LtEXP4IUy3guZCCiu70jm4biNx4xz+G2rnhidU6Q
JnyP0lqNDxAaEyQNIzlxMTJUoKVT1PK5/4l8JzD0JHxmZJpnbuWTEHa0BK9ECDvsIw5OcTRB3B3C
7LYotBW6yvYoZAS/bazHSilFeTrze0v1d/rzStx9lLGMeAloVQZVNcvyXfT2ulxJeiPnEJZEv3/j
9GeHsJSUqr3SfH2+e184BXnNxaUf4xgQGJCsgddH2vD5Q9I54ATQuiBS0tQSxP8d6j83tDrHJunN
G1M/bKUf9bCT9e2zruKadGEdFLwgEclspUCxyWF4OB7kUxOXrjBNdLRIsXYAR+KRf3Ji+mbPFiGC
y6pHeCW+CjF+pssg1IxItbTFrFPe3FRjOoctSs9fW1vemT+IMuGXvkax59uIIQzIdppyHPLxGQge
13PdZjYIWks+9yD/MICvuBrN3QNluUuXx7twBCp6xDsZMm0wrFtW+EoGktvdE2ndldqIqD8Sat89
bbXaxBgBrWLshfoHeIaKb2ocDKTPiq3qeAFqPSqEXZnpdtAop3nag2buVoVvlxsWs6jm8+W8Fr//
PG2dCLSR8yfRRi3dMix4bm5AjK1Y3qcJgVf4olLit6X2p/vskkAxAj1VSn3D+AiSL2MsqamidTiR
HLVLKaLPHtqoCoYB3ca63t2Ty5Z1iHUF8zwLFS1XCmkfs0IzeTqFBvKg4mIqtMXgg6jcXvn0mTvD
wRtOIK94hJANdrpzc3Pf9E+Xo8vrlAo7AtFRsHRItdhG5TJcrWCylO2lolhhkJezcnVVh/Uo+soj
B0Zz98kmFAu6qye4VYG/cXBOXzxtUiBUN8PDaoRXDBNoeR4QOPTTvT5DhHRZmvWdgiWT57178FZD
XMhQDwy1/mHJiYuLe7HXE8YqWNOHDOln8xmHogxW9eqjqfAwrd7DZy0sNwgcGY8TtGpL+jJvh9u8
dLJ1Tn03jLHiJebmkLvSf3JVSCC5brEKj/PPBNK27Jbll2sKuvIRviI6Qx4Ird8zvQPjxO+XLioT
xJAXm7KrCWWPlrVC4LZ/RUu0vYQrgzjYQrwYMfr8HwPgMYX8XUvGBwPqGn8dqm2VkqYlXTDPnzF9
WEm5ZBxJ/7W4ec/aPdgoUhFlrUL4b73PPawma/xgTEsjN5Je0LNTJTk9HNQIuq71BCHIZKzrgzWl
tuGiahvE4zte7wBk1Ekplw2fcVaA8vjaNmpDzzGabVxpk2ddPGPf+8dBrU/MTfVSnuWB4IXvYC/j
J6wtdKt3xIwCFTbZtc2sbhIIHQh/tzFCkuSGw8t3HVLTskTCMU0PiHqHZdw5SA1UkF9Cng6saw8D
6VyqsFWaBh0DsMcw+BeRS6/4yDaBkWicnRwLKpZmDS3cIanN9fJ3mMifwFl8Hz3tHMbpnGuJ3INb
jjrEWiBJaUy3GuYZxEhpyN1tW149kmlNqsRAqPe0hTqBVS7fymv1RJ0T6mesrguYFyRwBLnDtH3s
I5A0FTv6aP4qsnWuOBatwuYjX72o2JA6DBdEqbcEf4YuSzVYmCBkQQsTfEKFh5peGdEH7t8qbxTc
SuwxxAf+jg62zmyXXnPlbNiAWAtNFnQFZ5nTeNs/V8HZmrJKzBQiMKlVn3J2hWsr9/sv9hkIYCvM
a2AgfOunzZWgusHC1/85bn7hT5YT7uS/lrUNgAF85nnszZsxeG7QINtoC2Z9DJSPCOJsOItyuCE2
d9Eb+W7sxYHSXOSLReWf8FFwtywk2F4chb2zUt426xP/cbnSqaL11TfuQZZ7m/ycyP9v5JlPQMgR
uFo4kt6mcZG+/dV68Xu91UrO4x4EoK9hZjR+uwUBh/GfNr66U9Z+ZlwZQFyiPQmuqE6cCIDcIEIE
/267tXN2bFpaFlrese/uqx+xaJP98KpNqcbcXOT0BSKL/RA+x5qBkgQhgXhfyvqDAkNhJ0jujOSA
X9qWxpHqWnSTBsnxmCFEhz7RyFvdZ8YFovZfjRScEGxDY9vl0Q4ZhWQAFuUITlXScVpLhokv0cv1
go9hiTzfveacgnTKqNp4fvRH4IwWQlUhBvDQMOSaxNQnTp11VWG6ipOc+DMoxpTd34MsuYIBZatf
2I5GLYgiFw2HTOouyXjOulgn+6M0H2pcxYPLKtdD+4WsD+KdDIOfKcAt2enzY4SMnzLLorJJR1jr
em8YGND80+lmSFI+/3ruN70wD70CCQWleumjTsIGtpCxqGM16vZtaWVwXjrQzTpfZmuB5rwRFbRA
mB04xv/x1n0W7+oUTBBz+9aCRkwsb8rh8iKA7Mp/MMKjZA5JzGcslElFlxD3GcacaI+Jq9NzYFhz
p2rn9Y80oIcgWxBr/m0vBdhul2VRHVwUC8RuUohx8RsbdTzXqsmkDHI/ZRmap4U12Um7mkp1Zq10
0pOBLbaSNDMitKx28z8czzGGxaLy83ta2uVanZ8U1DCSbSenPOu1RMECp2hV4XskGSxcQ/rUbCjv
RNFxV1UUXbp+/foZhB/6Vy6y7hs4Ns1m35ulRjduGEVL43Y0FdwBCYLbXoklsmLFLq1ugcoBuYXi
4PZk/up4l11DSWFiERM2h0yiJuCoa1tViIXHZsGABjuqT5ZfaAL1pMEhsj/jP+Tb1R1+ojTEjqZ3
BBLBs/zL5n8Um688lB8sEexdfsJQy+jKQTDFsMHd2Bjw2kPe+aa9wE1E3uRHf1X2lfAXD+xnh/30
i1pboE4D5GjO5HYleRpbcGW+9WXVlA+NnUnw228P+4KvAqnn2iGmXdYsxx0vEX5N+DFo4NGDnV1N
0Q9562x4HfEIpzJfGFxm80Mql3KeKGY8L/hkZ4XnWm17L+eWZe2462MTYTAqqhO5eEqrzjfq4zw6
1Wx01qUpPOaCH4w4Cw/GXVYdZVUwot6fBQjXU+LphuhH5w3bfYzsqj0bQdTTnrufpyT84CgWVQAt
Z+Av3paqUWo4N1Dv7geTziqYI/aq6WaggdI1vsJ77XrcLc27doxMuiGtb0E2TtBh7pbNd2rbGv6R
BjqPRDcseIgDmMW/tXLy/RtkASrLvwUrtqvri4F9o3HmPmm0UPSDn3/v0jDVAsaBPZCFQ/ZUf4Ir
7rziSCIWWs5xG9pmnUIAcAKmoJsD4xwoG8zjkYdWoKZ88VpJcJzOCBcb5OAgsf+3F/3ZRBFg06BN
Nv78D4LH2PsIkMi/rbMlGeqeWBNJSiuDeIoVe69KVDeBd36nTDDlyjo8N+zew7yJJ1KQL1bfTB+d
TMBComEYwb5FIs0dRYj/RDT4+YjkfmqcUC7NLbRVZdF6UJ7Z+eTWGTwxJw9xs78FcpB+OOLmLil8
Z5WMaDT7P11wiSRy3KVrZJ+ocA3oWH7LFGsJjBh2eRI0yOXTn1gYAOB7LnGXLw1b286BxaC0eRzu
sS8wcRtPpbEDBZjfXw1a8T1Y+ELzZR8WJYH+wvb3/C9q9GHe7QEXkSIQL8KcxXMy9AJnIf6ivQTT
sd6qIoE1/nE38QYyTeqjbOgPM0zsO2XEnmfY9S0IIfftddBa1MUXfF+vcBaajZEG/1W6sBQnTRc5
ysZZ7j1lJTmyS5M3fvtzs9mCKKDHt7Vfs/+kdadjHBboNCFGYayRwJUl/BkAhJdjUqAYpf0P/rDL
/WhpQjXBQEmLSGcr+1/BgxRxoftN2cFNbxBD6a4Zj/TWeazz4aByiA47uGHKEH0gOIHK15B25Rfr
7vt3144uTVHwRS0gYEACe317hUaz8hP5hby14jLxp5y3bFOp5/9VobGuHHWzatQ3YlnKCYfhZmFr
cVTFuG6CiKMPLvry35XWnhxO8ec+cY+5f0asfXnKzsr8wm+v+BDcLM7VYuwoECyKYlkmPDUaOXw3
cRWpVJEqGlkg70qdrzVKtRVNys+1pnhctyNJfx8+yhHhprBlF0XArEtEsVMaB94X6c4aTYLzWZkE
lkQJhddbDXIIitW8h+9eclZXL/OklVD5zLAtJlPu6f2p6pce8XnT8hSgxC4A68R96MzIH+MFb2/x
s2syG7utdr/8FK7Gx100VvmaXpF/7pOY6w+Hk1zTdyqdVcNOXyRFkMKwU4ekCKo/mDE6uU3CawiV
Dy4ZTg2dF7VPFTBwvsP/gD7yp0cKb/aK4TKz7v9+XCYhWJdkkVsv6OyXPDh23a3rghC3dQ/nS6Gv
WhJoDOxBbjr2KPE0Qor0OlZDw9LA9L+2un3p8GEUXVvmSksoqfFOAkmAEu8eL/3CAhR/tiH9T7QA
d22IAFOkhXV+7X6aTnGMcJ0RyTzcgWvvrHCd9lhgSl69bfpi1CbRT8tOA5waIMeTnFQ5MaPnFJla
OJT/4XX0aLIZEvtperj4zCJhP+KOJgAK2Ps0W47xzff+UO01s6KJbbQcRKtM4lTz2hsGKxdQDGVo
GUIoKuKNKJqM8ZnKF6w5bCg9sWlGoNlwdcaq9RlkHYi+S7sOeI+4SIusuSn/vOTLzcMCkQs3H/YM
BixQo7WUWIm9071QJAcn8EMnYCFg5I1xt76qqJ2DgiH04O7gTNlQ6R7wrLpMt0ZCXxlS42vZvyW4
RtT95rnO/FrQVfzyx890lVSqHQKg5i62uUpUwxOD3j/TkTlL4wQijTH/8rEiMM1riTvm0VGNTZmb
NuiaQRYlOdk2yHUaeh7nnjUvEFQsvYfZ6fU+Gyq0xXD2Fa4cFkhc5/QX8mJnkurQ+wVYavh7rncV
ErOX0qGxJa62z9f/BP/Srp/0zfy4CXt/RwP0BCPl5BYA6OBzqKvfRc8EnKTyy1gKGgpKAk74bc9v
aMS4UON5Ha+N+Ke9FTbJ+7LPPXC+XoCloD3q12mK1CFDa4/TO1Fu6K0O0JGfpremDrYwF/P6/09Z
U5QWnJUKvvWa68wORQASt3zMgncHts/weS0Ut0nujEknJxycHMZ69Mop2jZPX9VAXbxIfKitKoiY
NLbvY/R9iNwFX/NW0ABTHUimYtOEmauK7VAJ6I7ajPpcrCPMIYHxHqrlmxqqr+JvVArpzEETVERQ
6sEhkM6VEUxQ4lrxvpqLkC6LyyGc7yNuGf7T037b9ffD4CduAE7gI/kG47eHrp3XXSK9j3pYT7/P
HpPt21fVM/13UbSz3EYcxiE00lU2JlMnoOQ8wC5qOxgukK+9MB1SckgQC5xb7DzbpUaAkTPqXw0o
FN8oBg+BEiTsoCg9lTGQ6kohmGXx1ZH+GUEyY9dfOAnipbf6OWzp242xtJwRhIredCqD7/96t4QL
8VyEcGUuCTt6nQ/Blr0au+VNzNeKxha/sJCdm3m6CBTPr+VcIQuL4y+IFYlCyY2f8dS7fcanLptt
/iVo0H5Ed+DRdTKwrafLh2RL4Jd9I8++kCkX48bCoaQL1bhmyiFKZr8ez7ZLEEArJHyMzdeTK0zp
jsRJeJJADfF1jFR0YmpC6EkZD4dGqxcnee1SKT1N2IvjBFf+Jb1KNyndRvEA1OjuG3QG6YnI8dxG
DHzqvF3SpiZwjF4Co/Y0ERQbT+fU6cMTEOIdjoKiluTdqxFmdU7DcDXoWV0Aqk4r32s5zTlj8nH4
uDs9Zh0vC/e46Crv+ugcx7HLAhS5HEsYUeNaAgtZqVe3HvPxt3pyLyByGa4i7km+1e+YPKmRt5Ks
v7KZyFvt14ZeX5zYEWu6CD8904TlBMXE8bG+rta9u4adDydtPP+Al4R0jTI6eqtxNWUag0q6p7BA
AYDV5mYIPjJ/Xb4tysI0kgExec61mfHPONOMu2xE3E66/x5JEygdB1Yi0dHK00Y4F6qHNxnKpSGH
ffpvs9xBZauWwqAk1t+gO476v/QStUO5LEBvyDvdf1/N4tirQ03oAqmnbHyp+5PhogWIfhTEpX5R
wET7RqmC4u9vFOhtoo+WMl7dFmTxsTBz+/vlVO+2cw9Zo++XODtIEHPcasJC9sEYHGpqBUMtSJGh
tYCRsVeazsvBk3/9AEpMKRAFA4bLhFLDJWXPWbxY/POAXQi3tNNwy/2L+nIodIjiOG3aBS/Q1wdv
VcVhejO90wJDz5MOzDfy2wrUNxYYcBkkv97UmMFTKgWCDUacUlSXG0F83TjitJkibwdIDar09DO4
GqXqJyLXMqbQJSiAm6b1wyovw/6QuDbb3N8MJGFeWv6yLPHu7+CZQ7taeChfsVtQ3NGXTdKwpNy4
n6Jdh4tmhATLwVKdppI6H9RCv+bSwaGe1JXLKF+BhQvLdq5edLQbt6gkzSeLMvBRSv358iNU7OOh
oMhxAB7bPggz5yT8qDZFGMwVZkcFGtegWq5hfUV5iGzig5E+n1aKAOxm6coEdJqtHihimvoX/uww
QW6vLAKFbDHCVmHOHeloT+dYclh9ry50ZU50+eEYA+kQnmrbqEuCdk3L9XMK27JiZZtwLEw3jYgx
l1xCAZR2n5EynhEP04tFe9TVJVtHXnAKJbmcY2ENaCJ5GV7XqSmgCv4qjeIuxdf5bjkUO5tCRQBb
h2Gzu9mMEY8h167GaSlDVgUNdMXj459xYpFyZ/oXt2HEgBQ9qPmpS43ItXs9gLLxLm7w8+or6GY6
XCVIpS3/QjY+/ve4i+j8Op9G0ABSmVq/hkAdA5cLZJ4cFLTeW11jIVvNdyHiWRsP0amtl2IhjVOX
jQ602FkiEVEuyqe+Fq3FARKxd+Ojn5PqmJZU0t1o7TC6ajE0N+YGTpw2Bn9MTJJYcw4qlctv6fPF
k/jpHOqaMV3O5DkMrxYls67EdiihSAr8xgxOjAUyMWYotrI+P4XXhUQCeHOo+oPwlQTQI8sCK4jH
Vmsu+qtYKLVu2hqoby6B9U3Op1aqUn1V02F9n5vLuLV1BE1Q9kVQh4z2mhNC4mRPXSmpinkBLtSc
1hi1qXN0UVeyNG4rg3R4OjjXT5g7Rn7p+ovYVjRKAA4W4xhYEwJ1XS8WuZEw4V/i+lJWO+Ew2bTk
umaQ+nMBDK3l0HtGOw+Xl8jEhsDszFkl8tlQWhIKMu7z0duwJLHjFR5/OkTxUPlLkfL3K5J4rTuN
9vEW/PPFVRI7jqsbyI5FjQVS2EH2grDrZmgWRCewcsMtt35Wn4um0RfueUUU/qyCX8qDhzFipHN1
o9qZ7rRUgHKwXrG8FCDhlordAsGOD+3VYWhgeLatwLZY7WnJ+qhqEWhX2MCxDNxbBIrnw808CY+k
9t1OkECyFN6ryvABbTRjq/pkOEgCvYf8saPpy2vsN5IqXPNu4BfVxcRqmbpxK6ZySic/QY/94UC4
wG4FjIVpTaHqx/+0wpV7khflyoZ3S/gEDiAsbia1MLqRfka4o1ubjpxoOSHnCpWzVwzzv9GnrT9p
+3l0TOfLQ6CnR3b4QjVAtgT1cpUcLQ76AO5pIdTRhnZQu6xfnsGRQy5A5C9Pu9+RP86vAn7cHzQM
2JT6BDf1Op0b0u9/layuoHRSBnAZAHI/xvr1ZqTQcOr/RQYi8vGUDw9fti/hUN0t0g0tSTPFmf9q
y0x7IQLcRKH2vBjG7U2T44b19SJ8DiNuq0GJqzlKwvVxsigS+PB2tDeTSlYfzkA7dBTgR62IJWun
wGLKAUf++tzT0RSyH8mgSKbnUTt3RbzMaZLvOQT/6hbi7C80+1KeEzmYQGvTfLJ73F3LhLzRp0Md
SILhXpK9DavB2fM98KxJc+/RYUdTCP6TdbeAgUkv5aaGr9gHBM8N8NZDbNPWYmol40iK1WQ+kp5o
PXaOWTPb/xPGg2QsAQVSfaBCDYRZxMe2yh5uTWSfml5tfh3sybAy4tjgkBphmhGgtbC3b6JsrTY/
NGJph7LOMZI9nBPg44ZJAHG2WjDEor/4DL3KoXw4IBhbbuE7pHAFDfJmkpnXRk4ZbQG7e65cwEWf
KgcU1KKkDqwFz8TwvAkfFx8VuW/RYw41o1LCnHD4QCSB253OQmVok41TeRvj0Knk3VXYqbxbQ0hm
djOMDiqaNxWFrYbDCt1XoJqE2Mex257L+3uvRjWFjpqlQ0016FM5XGY1hwpGxZtq21/4trf7ekFh
4GvahrsXqiKHGNoTsJEMxCTKr77fA/jsNpE4F9RBaI9j3cio7vK5aghHjQISYuipNRCmxPhMA0/y
nAmvgCq/YHGktnViVPmvVHwchjw2cI2Pc/j0fHmX0ynlHrBNg+iti1acjSdrXcDy5sCZo7gOSSuQ
SoddYP39D7eQSXeSBBl+2CJg6S0UqEXtrcNxLHiMbB9+SHdWVuTzaQO1HDVsQ78DKhYHxEZAkmOA
+9jiSjN9M+6rnJJ2MPu4Y8+jzzAQGLvNGU7Kv+ykBXVcrQxE+H9QqApHFEb2S7ew1jdJM/ny+yjc
MAMkiMrW4iDPCXrQqFLdTTf5KsbuSqy91ympamnT1VXJZzOjE8NM7IvNSQzZrdNL4FKSsv/UUTNJ
wSGcuDIbe4xRCrdvR7Bbv0YgTf1Nieqo1Hzzb1YCC6mOfoNnSpEl/3nTQ7RoPnc66cq58bUbN1Bj
/uUcdiPW55Nb5PJBuK4VOcLwvMqYrerM+0z9bAOX5KIt7owwl0pOSaZh32wPN/WQlJj5FsjPvR8h
qzqEiK88SemAaGx1YbBo8IH5sOnbB47f7JqrCcE29o4APO4anUu24EPfetRAnDHT90FZxwrrk9dZ
wpJy0mYyZlpJimJvvfpHeAoUvnxk5Su6sJvNYS+h5P98lmlG9RlYZMWXm9lvPf7+iIlkzeFevm9i
fr/ZgbUOiSmdRCSF/nqdYiNT+xT5yaqYDqfBYPPs7rJvckQ1w2SUGbHx7ToyVQ8VDTXT/ZFdIX4P
1lSvEg9kCxf9fndbbxvz7oWsm1jzCL+s5LmOPbBeX6lRHre3tHpifA6/Q2VE+Vc4mqYKRITJI4rX
ua9SzPZ/NqpR+mWOpumwI2JCnIKX1x0FKZIA+vNg0hzIsElv7dD4nYo96mHsOM5hYg//TSWgkbhK
WOvpNWpEbgWfq8aY9z2kgrbeBAUy22uWANb3Clie8DWk6MNRNYFif5nKHCqpt1Q24sH2WfI6Itxn
+2qevMTPaAruBUZP5ZsKLBcJurrTJIJiScA51O7lCR8AjptuQm9SeYWQwGVsWqfea2gBKC3sNm3R
XqabIV7DUKvLfNQyAlqgdG+JXRr97KVCzJTyepvpszniCbvHHpmyTdEPW/MCrXU1IJj/3siFpTPf
XfbUUeUNaPFhcD5reR9CQ5QtUVP8lDPINRyaU2QcT7BDT7x4ussjlcrkAabm/hcH9ihbBPPSbvTb
xk0+CsYlCT/ihRP5QDuG99210jsgF/8VdxOPaHChBgPkRTFXquj5qsvcx0xk0P8DVG7LUgKFIwYs
WRbzOEFllidCy/qZNrYtuFIPrJUZ4UeoqMzENkF637lJ+KArYrbm0dNLX8Q0BpdR7lN/guVQefS5
2UmiiMjX9ECZyCZknH+6j54Q4sBkd2tzBZDrEco5CPvt7IL9dEQRPTxSiKr64JPc+cmjHjDELXQ+
zlKz/QL2cMGPKesAbUyPW9X2uRpGYUaID4NFIZDl+AJorVwnOpvxSeO4NmoVaiVX+9Y1WiqW9yLf
nk9/SuM0+LJj9D9cPdgzrHbMYDsJYqjSR60mADI5Ij5e/FgFtHGqAivzP0p4pw7+Ngbw6bJ9yEoW
QQl6VB7HhZrRoUoXaqQhq8m+xR27wVEL/TWS3ab/socJBXYLTdznPLKnQ5lkR0awaItXFeZfb7hg
m2aW0azJY2lNc202IHd4zNsXMW06hRqcEUdeP9uv4G3nVwPbrxIC9wRbucZmiH3O/Jm0N+bBuE0l
+jVZ6ABGmyUaLQjNKq7ebdwUEmOvoR4aHs439Y3sMRF1tR8yHhjaWYYYc8n6wRMoydTRMbkabSsh
FCHHbgZhS7aSYGTypybB6QsJLh7uChS4mPhql+0o6/3ealpqO7XQklHTlfUE1q+7ruLSBKMOVqeu
bsgOU+MZ7iWNjV5d5EhGejh/MXMYKNF6VjB/lkoOLC5z4J1+KtByZYbOGZUHoeRpTLxjlYyG3bR4
SdZl5BKI79Q7x6Mo7sQadAHpL7RoDzcxE4yyuknb6tVZaKBiIg6Lvhs93ulhnKYF5Ini1rth0sLY
zo1MYZFrPWTYi+03QuGCX2OXAXAPv8lp3ji1B3Hks5TfxEQdGz1jHESjuOZYKr8MHlutst2QIAId
lzYJ4ZICCr7lCYuiVZ8tWGMsVQNzMO5WkmtkWWMSehsfftyf0bYIFqonn8sfsICZF/X2q2J5iFFg
ZebhkqAFnna3vUI9L5DV5jZNERw7rqzerxcUW7iJFMDWrtA4eJnBeYuAubvLnfPVErN0vehUyghs
7xxPWECDtIOdWzCTCTJeAIUlvAIj5VD9QLQp3WBrDZybV8zlslrh528xxHeCfm2zfGdAn2acRVVx
WXsDTny/+NtBET3NbgiAgudOgb9RiLcFchJqKlyf/ESFfht6nT01io20L+QeEJCGeJ2TIn03H3qk
ICNWW+QiZFNdx+2kHd/laAxQ/oemKvFfiHJ6LOgOwbq+vYnq8cvV15qwBkaUTGoXkob6lr1bA5F9
HocYUAwW2g+HXUW43H+UGScHg3ssVezDboNMxkVf9cbIClb/h8DWR2uj4T9NJFoDX17Z5niduJaG
0LLdMP4RgeJM3c3tetE0LH5HdG1r2lrXXOPawZ2CSY8FsYt/j58n6ojLrnF1ooGhubtA35fvwS+c
7Dp8/rInKaMX5d5Zw4fzJmGJxSef2XnsqjQ54XxKhAuf40/QInP1ZHz45Eb5tTgHvZAYXAXaJOH0
265RVoFVZGRINOJ7a2z7OfxIZGQ0j9jCUNFqGpM+G+wl/ZXWj3f1Z6iuK5HW86WbxScQb/bQkFdI
MpICR/A3It/JrKHeWhMNxiw0UsnDmtnQumNSj0bTI/71iydccntQucIb71PIRTa7VV4dEwSLTo2x
wSX7J2ViLyaNSYdy1v5qVYDZs/WhtR8WWrDcmgnxBsSOmpZP/XD5P6JvmaJhf2LDFBdLVHcviJza
afHQ/CZIIBcfqtVFWRNGlxpwo3Uz8ptyVO26/FXyugTkDA6p9ynkWAtzh/xOW9StZzf/d1u4XRi0
hdjyMZHbOluW4qeX2KwCbZ3/fyp8i/vQy0ZDYOANnUS9YUIbUUsUA8Dr3ziu7xv8suZANwFllqEs
rKSIoT/SfPZcVkJ8aiUAVpkqtWz+ErDfLS6EveO3zMn/2wWJERExg9gpIrHH4T/eDwjvxJkd/jaV
qmHRhq9wUUpPIXwS9dImGGXu9PWU2VhItyKkx6tqvmLxsQH29/L1Kcioxr9kBdnXjGAmdNIU/SsX
uR3TM7206eeA9BIgGHXJGoVjdo+9ilgtp2p3+Pq1GFjlB5Ym4FlsGhbjYXw1xw7sMuh27QAPZvM/
V2SZt3/JKOTMAAgA+tG2iIOroj3Eot/WFSwxxOc9hTodbJncvTVv+y0qNMBB8NnlRxKnfKgTtPTO
dBrgkDPb+fj48OYPqW5m9p9U/PQmtpeNQjZAr8TIbWDcAfIJ3SkGzFi/PmngNoMrDLLbW/O8q32C
LcGAfCIKuHMfc1m56mBcSqJ27bbbFv+yERcleN9vfaAgWx6nwmgY2bLhPC7fPV6gTylIyu+iNrM0
z9LUXtboqaKY/K1qC04w9YtyLIyrZ7oR51qIq5a7J49WD9uUy0Cpqb9ny+vSh6wsXZRkJifjBhYB
LWV3Png+LHSqMMvH3HFpPxgOktbFTpwWnQTk7bNShFOwf7i8W5kmqJuS4s7ZAz3ZU/D6Rqr5b0s6
t71bX+rKIUYibhiCNcpcZS4O2fmrqWMtEHRXbO847IdKESF9Mg8MyHx92mNv/GUaIGCKhbhCCBRe
LEwb0UIFQF99ej1LhSuui8PWyimfiwsp1Q7DiDyNo7WKRe+koFPCVR0rAaQ7Vzm/if7Uv/rs8PiN
tzI2DSiX/ECFLFEuFzEjZx93hDGlDBIL/hOhTnr4dywp6TV3rBuNAxHZjs26TdU1W0h0th94BTE6
3bv2uIF1BISrzFcvRTVTrAr5I9a4RrHgyVW7Gryl+5P5POfFrHHySFHNxCfjW4C+DxuHcBEa7AK/
NtX96ssKHIkuD5nHa3y5UArc+AQm/JC8Bj0ATSr24AMrBxFe5ghCjqSJofbBmMO645rBVbPX05Os
AhnKhaEPVLODueTpr3Z2PDESpJ9x/XhtmIB5ZMbcXQQ/arDt2vkRrWwP4M1sfOsDhrY1pWDHPsbq
6xu4pFhHKqrdpbrxgkYJ6YWtcmmSjGCybeOVHgvO04S9JEd1d7UsJP3HPPXGqzBqhdEt/n+njqxe
2Sm838PblrP/429l/mxoWygBFr+w+A2nvdz98wNsr63tXnxGErXF+D1m8dwlpjOuZ547w5tgOBB5
ZxEy560uTQoVFFquFbPGYk3CPMadN51f4Ea4IlMuSMve52u+DI28+br1NHPNYrKOxk+bbFX6frHu
KYEnzPnOCZjPupNI4OdYn3v0u4Yk/O+xgFJ58BaIhEC7C46+xUzuHxNh0yNvJ48GLvYXi86+hCpQ
sRYfo847XQgz/3ORZaB8rtcQcPcH8fUeoSlbW6gbP3tqxThYmNLwh3+knCjvY1ZDs6nC1ABu9C/M
2JRJ2KDDPRoHaVfAuIwttQY+f+Uaokh1tsRhIxb7dOPbPCKxxxfML8aqQ+NpU1lY1bW5cHgthI7W
qRD5U9PneIeXQFb3RPJHiK0qgQQZ+C4j54n+hsyXFEWcVoUzRYMFBxhtTJ/4XIM8/Zz/CNjUWiBF
vctL3JB5G3VzuSKrjazr6EVmAZ2EfRjMqxqIaJBevmEmQP7f/BgPrk2m03rVrthx07oxEX8Nmgyu
SXKPY9sr7Esm2sKyGbS8sF5Hb8kNIdtGy9Xqd79cj62h/fsQPgU9hKGgJMzihN1jMjcnbRPBliKV
njmoDByU0Af0iRhvs/tXU+d5mndY/cJFK7Tb5PonRHI7VDl+50gM6w09cVuIyO2bKm2vp9Rz+sGk
M8zdjd2Nh44qTLlTKVJvKXBHgqiXSEC09cL2mzx/C/2E1kmorN/yVwp90T/h9kPGZrFu8BNq+qAC
yWBoRTWL00quIxPrzWXR8pDs+wgyj580S6KvcyyNaLOn8sIm4ARtY+9VMsdqne+3Y6f8a9G8TMiS
La/GDf3BaMA7wUOObYibBz+IQNdyeJAwqRa+F2I59tMU7CCl/KzkJTCNcDoR8AfixBaVAs1kX9PO
bfhG2e+reDxxeemhN5u0yJUcGrt+XLi3iBCDvxZPwkjfrgO93JhVbIVUtVNX3FpA31sum5jefjXj
JaiYGWknFxQ6rB8qGUvwTocnJRFfNxd+1psfOc4TpuVeG79qmNh5QURSwEpeWrHHOJwUVoTJp/Wp
hMmL0XGM+3ECrBd6W99pbYp9mY4BWLZ+xxO9Vxe/3Afdweo4L/LRZgg7xqrOmdZD691jMsRtyLUs
3c3TS2hBH0xqsxV4rCAjZ/71xX8p56I9tQ0isX6pEpEJ0ajEJExRvneXkIkWLkrDbZAyChFrZ9aD
6cPPOQ6ZDf5vjFNtzbIxF0qLlBIZiWEo1v9PZfG2p45bYB1JRgX7NgIt799wzqXpDCGVwXM/pmUC
gnbdxuLf4ErT9jJllu2Ghg3sUOgPNJ43YXWyv9Q65u84rFGksTRM8ea3wCctpG+xltmqvtqeJXSC
W0AcRzpYJYIh7wWLD+ldbtV7q5OZ67jnag3Ik7ghKfYIDOYPAOojI72ORVVU8mo6Zng1qk6tQbUf
L+8Ou5MVGjaEm+KOFs8/xsEFaX9f1FYg/hvGL/EM5nGKgdbku7vLx4oJBT/hVIs56xFj1JP3Lle2
sw8NFggQ9pf7hmIIcDKW92lGWB7h1VQFP9uYxAX2PhGiy5uQwP1SYGRgVvlm4yA5fJUo59ma6jpb
/aTEsvHd76WbElyGFSRAavfv57bDFWv7K8BDKklRfx6fI1Db25H/rXcRQo7zjiBVCk3XneOikf2p
n8KnlQAfPh6F6Deey+uHojSO/ttROVb7BcyT0bfCmRXATzON9nz2YTgarXhys1qeII5q0dTTU02D
h7bhte/VVt1Ax1uHlX7JxTuXJGPuEXUMgkFwebPrdAZNk6eaPTBIWFtuGfBZTzGFNMIjtPoubq8c
mJwUMXWuf3/cdMRuw0VSnwx33+TCMe+t2iwQXQPAwR6Pxd263xTH8779UsGqXYEmOiElFv3MGf7s
fwa4pOT4OTRFWcbM2EXZNOw+lZ3um7kJkhWXOf/cqRgT2kleT5L2vzfog5AN652AtG1YWmzhwbe7
vssWPs4in//jgHz8IDkeLm4QwqWCv9AEV4y7z8/KKn+W4ctVuuHk8MIvpQSwcXml1zugEvjYCmxS
OTtTljGl9vlt6ZBxZKxz3ohfS8ZiBBnYd5tZZc6oMKjko18nffXibtOIrbwezQrOinxY06BLKL/z
uUMMlnBRTohxpiD3gp78BEmm2OeveoBfd/gHkIGIhkwzKEw/GhE1bf1pbg3DNP+/p8br7gGXvSgU
NWLtZkNr6rQU/GZUAMKhv9UvUVgMcDLyk896+sFzvWWnHAAKxTkCf8Boa4BdQKOkAGiXp54uuHdT
NWCPY5oGGlgxwPn+sOol6Yfzg4alvPnvWnpWGba4DTtMAes2RJwkSGW6iXeXQ3YlA93EAkOLsGoF
9DJwAPR406wFx6qywldHf99qyB/XbDpnhJy5n/jxmpVQJTFC68NSfOrvJZc2WtHp1Bk9dDzHiKNm
pmdtSm4ywiIKjitdHxMzqCG7nkFd2WiDQooWEx6thyarZMi7kGftkSgdvw8ajMgnBZYKws2/g3tp
TL5fTMiL0yUcfNbaWjQOiZQmFoDjSE1xC9tLh5GtTK3d7XG566qM0d9VuC5hGvcrs9Ztat2m1Scw
Z9PCE8uCzn3K2LPuefNaWXNzChH+Q0hcreAHlw0utvfyDT7sWxwbe1TL8gcJcI6asPrKAF1bWuIT
XiBbeRiAk/G9YkLFitbGRzK9hz1HeoPw7bw+xIPjonza2T3Bgk7C4amjE0s1RL+cZbpF8/NhHWtQ
50//dXpUfsMDNo0gq3tprvYklPj+gg6QfUrwMss8vAKGgWy162+aWHjWd4c/Z8FSxS8jUOTGoUiO
9ogg+A5BHXmJbK318KwhpyJYUmgHCWb+WTjGwhKuRIiJLssJ6yFwuCdYCXRTHG9T9XaIVryLibTl
EpTZx99ZdUt6tGs0Y2IgaLGE+ZwivKsaKxDq3UKmUUkGn0qx2u5z3/yBOQdqapK7pUoupQLhY1B1
EU9079ay1zN7O1RTgZpdHUBWlnmQZDAXi7SHp48KRs2mDy8mcm5Wv0fuwajYKxev3TS4Lv7fXVQi
K+xwKCXVdtUnP9IemgqEIZPY3SLlGjQNP5LEZHIK/GQ+TD5VhCvJ2OOE5TAyNTEn3q6MBuo8B6kr
n+vGGoyFTGe/lnL0cXqvQIwG7rid/j3Mf2Z8zLU8vnSV1Clfglt1cBBYmd2HwmyqQHuOgczPwQ0E
O2O33/dXWfWvyyzcRIFzCWrXMk+6iXNDEosarTqXd/Q0mtaJyJliw436iVjomtWGBr5Zt2rmu17x
vKt0rM0BoXICV4gfbP6gVTvtwuc3TW1ghCMnqYaGIOSmN4W4i9lJ5rQUvpXIVfIBCyXdey3qEysS
GxJlHs1bX4Syvpb6kJ+QcI8WKNTaIxDkhPQBfYP/mQKCJZ7QDFTtnhV4Cc/ccdVUqg9Q2jbGQBuD
x2d0mD5Zp7uyVntDyB4KJGilxckXmqdnaYhNjZGEllhLoEzqxkWGXOKYPXW86Y4AmLma7An4SPC8
g2LQURFwSqNSaN97xZipw6wOVfrO4HrRn7R45VMF8RnWdbOS8Ba0uAosF077ZEU0W2jRvVkJ9ebr
Gf5roRYjLkmBePJf/dmEMFvRg1TEOHOBIrIsZjkm0U92gXl1gITBICLxazLACuRJSpVPceo7Rh+s
NIA5nzvSI2rgw286qeUSQYDfivtKirippToroqjAVzEpB9azp90JmDFXBUf2BYJfFFF/m1rqalJ/
bztQttme/YFBxcX1TOQ/uFB2gQ/JAzh5OJFthmsMZl0n7S66/MgX8cvZCyeKQduIuV19c/SKzj87
w4oQkMWTi5hWfTZslT0CX4zp7bZtH9avVwlvr5737WtlTSwMJfx3otGkZGwcPZAW1MsIrvOsHaar
6iCD+9JD2C6YCHClnBXERsi/GtMrXTyeOHMpHfvKIiS4PHpRAfV+MKD0gFleLVPxodOpe5HAkPRZ
x8t0IGJ6Fu7hjjT87Qw5v7YhZ8VqNrU9V01AqdBCh53fVjIeWtZasM96SnmLDj8HFwarfnYnlDqY
ZVlZymxHFjSb39lvIcf1BkzFz8WzxpddoA9peta348WU5KPVzO8TAe5rBy3QqnOjDatmP1DVC1LJ
5o2Gejkm2umPxDYyJjd/SLUIuOAmZOaFNA47steXJVo+f7Qct17eiL1DmgBhjDzwN7i8bA5SkV5u
2L1F2D5eJ38G8VMT7cQxLVSgTV2xCLnd1vGz1ENma3L6dHfKq6whY+tTaOZ3lvgD/mWaDvXo9166
9j4aXnXaeLk8s42AM0WerfgAZfDQ+N0UfEcHpMNONYOWi8rBHxF0kScBmGF7y6qd3O0T5QJrfQLu
6d1TbVUedrn025WrrlwfRR9plPYA0jfH+b876HRfF+xWELzbPAWwZcFFfhCJs/p6xYy7WpLxyiqN
gYYb0W5RHEKDURBKt+/FADBFFccqxhTG1tG031VHTc10U+csMq8wlyMXt17WXwzoxna+qu7EaMIQ
llgP8GaZtg1LDfng3cAQw2QlEiha0tPrlYCSFKnYrpGFEKPDmKJCSqzlhWWVLqM7SmL/ADDKNcvQ
/N2+QEU6z9jioSZY/TY3zNL+hiOxiQsnZMqx3H70/099Dyp3Odcq7xl5alkghkV981mEKXqlgoGU
kdIUPJTZJGCZRmQt1Rp0qrC4ZrMC4U+O+EeDENnPuUZ9y2097v495Cli1x19OF4PHPJgZiizNtKg
+75RJJzj2X5PwyI/kIlh2mPKOs/DD9JfC1EJyqRFazeRdCZ4vTA4MOIkWn2duK+1jzrUFBn2/WXk
HjxhAKtmLHYZtNipdqAez4U5y4c+Cmx+rztkHqmw6gh8mQ1R87kXQCjiiL1Vf4GNd2uZBydfwtc+
sg9G5QiQIsUG3dvnMjkrwxKk8/S/6AyZTDQIqKgJKZg6B689jkTqsckZsf0Bk5eQNL/ucGG1E/TS
DUTYWOls6TuW/90OabHhNIWl2KDgzOSfVxfMozRFz+LpKPJ8IPzWvnR2Xeq6/7oX0kySrWwseicm
CTUxOvry1bOg3l8vAlDWnhmwwlAaS4fpLKyDs5/5bluOcj4tZbWKbt41Zxzg+K7oDNhTMiGC+HKy
K9kTCrj8jEqbnzmHHhuwYmMYVtoohKcatlx3fCQzihnJUAwxYRL/X8tnUM40u4Eivi1xw7bjjmVW
HADCU2fwKAvZk93f17EB6Ype+3kIn+MJdT0w2r8jkd+qH1JsZIra/rIGwuOINA62lUFJqN/tmApW
ZAoJubn+/vE9fIpCL0na2xhQyVid6E0adJz8x8d9HOayW+L+nHZaFIwhTe5nTj3WnufwY/PazBeE
0PXflr/Cu0+pdhzD18RXGyrqAlsqZRCfeYf4NZebSxlvdBuITFpmhbaXzENT8p+HevKRQtiWJ/cW
c8uLnY0qaer0B/QIN/Bhns4qN1jeX12JPAsYZDfSdEbq/8wIxifGpZjPiHVLJj8m73I4ra5V3TZY
zUQLGee+EA/vqTHLMZMR1MEVtLS/kXl6Ce6BWfIuxnigQVQ7yAGo/1dQwtciDxQaZaqaPQcVX9yZ
C306JRFLRcy0vR+UV9+6rwdcmmQ+ysYL590VvTxcd09a2mkAtT3X2rmWBA23CMpjl1e1gTCZ8lKM
h5WouVLa5a4p7Dzb68Xf9IrstaXBVDbJ4+IMR9ZPO903GsS48h5f9SVsNkihCVV2tHO5Vq3MdrNL
Wn8iHuNho2qp/ZqeOIbppv0QJ4s9vo9yDAgvTv0oXXrPaqlivCi5yOrKvrb8ZVzAiUXoMVp8g4VK
/1ndQAIdU6nFY+EO6lW64vARD3tK0+TyJq1REvaHk7VrIjQCKZOoFYufLpoY70/G+BtwTLQC3V66
1oAK4Jcx1fQdahgbNSPHRHzfXVSPYPqHvROy0a6UxUI2Rul6qor2Q4E/uuNriX1gPF+p+upbDxBN
HyYsKG/734AlBUsSc8GCiXJc22hKRlmS8dkponSmExtsQ3SmdqQ5JutVxWdvNrFGIN/w9/eZylFH
3gQwHHDBj3I8ehu7rcVMykRwkRiWsF+64IbiHEZ7zTmNUWhxqq7KtoA/1bi+4c7R98jLe6XUIX65
HNffOGIzg8Sw1TDTbu0E1oqOWvCvWo8a/HPOUG4S5a4G3v924O37XESbhS41vFkXyrlbyItmtn74
axUfwbmmkn+2LxRVT0m1thZ1eLKVIzDCOOKcHj5qPYKcW01VDAwGC0/O8V8WIkR+F7pqIfpj1IpG
iak5wMzrOp+1Rqzf5GR9OsrT3pc1SUvSUl7yzmX2qB+1E9vpIgPZk2I0uSsoUlCZyY4/ZraPuqUP
u4bxg9IKpZYRBJjFpn+ro+hNYO579UAGCe+wBITpLJ3tr/k12a86z8z7zfbuiqE2NbGws/YJjUOH
9AEx+9tr3QXGK17Y8Tjj1VuKEaibAFgJyPMiqml3L1JtPVupr8571En6dWOhOmKja6PF24en9ZKB
8feK4ACbqLKG2BpmWQvk7lmthIwYz/5sf89E/VU05CP226RTCAHOuDw1P/71TVrka90huZiiXNub
phe5nkBntVXWmshSiWyL5QSoJIY8zBTrQt0Rdgnk7za6x2bdDwhHoNzLPOHw5rxpsCQv/GnytHUf
f9BDCYnwUAn5hDPYRyUz7NPIyTb1lcKR35RlCukdNz4LA2y6f2a69Poud72tglPpFjUgAH53nTLv
9exX7kFSa0Zwst+ho/yOuyqKN5SdrxxCxWMrubi5mvyeyzVQghCRfTHPrdPQPCD2TJ3iam3eVQK2
D81vAxMxhSWwQ3Mnjz9GxUPO3EFdwFwV7RQkwDPOAqekG5W+VUn210KR5yOWvyLMb4CpJR1ztMBu
5drt+rRAiveRGh2KymtFGTxaDcMD8oF25F+0+UrevV29cae3mAUwG2qxPg+QuP5QfxTnBYzvQ3nN
2rDevrhSJ/uHxffdKE7qJwIlF+pQSTFcaGX2TqRszNVM6v/Miny45lDqvWzIFc8W4W+Ksia7YvF1
gNXBY/jA7hNQ08NpfQpk6ycOCERFq81/acMXkrrawtrjSGdFe0dRSGSFWaF1F47xhgiS9EUXGhJ2
BPZ0ioJbjN61IewZa+fKknnIUyyoJCFHUmfc3t6OtsaDhvMDElBcPPykOuRuAhB8y0dlX1/Sjq7z
zrJYtsW/2HCByx4TM8Rep/3t039ZUg7ZYMpTNA9+pYqFe+UMP5qNEyB+iQrjircDDUwysEAO9y6Q
pUABcP0lfT+5JByIekl/XuD2UAH0jGS+90JsVIYl9IeiIPEAlJhkg2UcCU4l6X0ywRWk7BYSoeIS
fQSmka8rvPCNaI9Vcd33Xj4CpBwf/EHN8WZbRduJtdrCaZ5c1EQY4LJJrpc9CwNDVlve1VYrvrU9
Kxb6OW8dquY7JAUJ8CI7KWct6ulpF3ZMQab+YDqQmGQGLoqQkScgRq60v3zPHYEordulMlVPhHZo
aKay9NPI75/GPwEgU72r/UOAdzDu1Apan43BUFX3fm+0DxcnioEVEZ0AW2sm1oYzwGRLjQhDQ3nW
2/vBITDaNNGv03tyro8MtH8usthCxQ5L9qkBq5bouBWqrQpBwKuDRHZ8+WkCzeQThBXDRtMBnZbI
b6e7Og6np6I4aylG0xDogAo3UV2OFk+A69XOjLXYyMx6/aTN5B3vYp6qGoHCTSMv0ET5eH9tlfTk
wukuv1eKxkofBaGspIEKvAgyasC2j3ef1ee5IAFOU10tMli5IYtBG570rPZqSsueSt0sx6O5S8A0
MCYTeUj4dDp7Q2KpXdaCMoEWGtSWd3pkeEkHE5ArEaDiG8JkyxBRtO/RFDqErXZlwYMBp1ce2Xx+
hFZQ2Abbcqoj+b5KF57jTZtGQLGUSDt333qT/gloamgXVfK/qY7Lc7D1f+9iIabR85+BdaSdxHFs
pWP6weEjStbSPu2MnFPiLz3+Wj2D2v2edsbuwE6cWu4pBj832XYrJeOhgioMnlCmbRm8DNEyIK9e
l8jfy8LCbH9yNTq2zJdkaYDi8e0x19kp06rTO7uXmrYHhZ3VkaSxh/5iRTHcWsW2DTBiLV1p/sRe
gX7Q9RKUS4QsniXKHe7Epmu3Y2Yu8LSH2lMyL2U2jmsCpFNfD695aQ8BHUApM9CXWIFYzwMZS7f8
Lo1NJy4siaOGrKrO0gVwJFbqExKk+BeqDs+FdnHzSHfLDffc7++Xgn3VAtSdHuThbaY7w6Kwz8sS
rCUKvD73GaV9hQatY5Up3tNhvuZOMSkvzFASa4vaVPBoCRNb/+HarzM0dOpJaGCLb8LumUlwF8x6
ajXgsS4KYUTW6qKHDqYHkRKutP0pXFnDqo2wza75nob5HerLqotxUEKxzH05TKBmWbYoWsWPikkf
i7GnPYcosNg5mXj7MUgnk8Qb3smdBUwRPDS04vPCfCil/ahIidlmMIO3geZshVE8wsr6xSKekR43
Cdhl/2XcrGZe3xz+yTx7LLz1Jw7g10Kb6xPufDU+Ms9qufknWlTvCDp7+4VRULXNdjIt1/gkWIrM
gbgPHie1ibqTUqbKo2uH7j58/QsxC+OIBuXkPiOoqwJ2kt+7B5VGLETwX5q+j8WA5RjjZbpH/dHL
48phISWVp0rZXK/ATLDIZ9p7uqDCsaifo3S/sk2/ZqsfVze+luCKK/ApqB8wZaBD6M/mfXxTZHXa
bBe9j1kvt6Sn/74JVOrBkr/ymBLsaDik761TUJk0WZ/Eu4bjs7ejEIbomNf72TenJW9aG+0ggIoD
V7cFAwb1S5S+16wLglzu/HfOxpiH3KFKD8820DP7a8Anba1rcmELNfXxUXFztilbiymFIHggUDWE
pK30kqccmXoau65Zes/AUiI4m3I4EyHCh3HvKXxunk+rxFfEXynBWsGKMEp6FKtjWf/TZmxA0jAb
ziu+//1/UKXHgsg/YoG4cRPw2mynNntBN45uar38mj4zhBucrjAeMF59l1iMn4nlwQbvxjBXGJEc
DptQmUowkxkmg/mAkJl2u4W/8CKKopRn4Zss+CapPWoanT3LOHp3/uL0bE5Beg3UrU4rUOesNruT
E/x/LMd7gqwNJXHqn4Uc1j9y7sS4igDz3j8Pz3D6BlU8bvZ7LOAMdg55hE5ayTpbrVix8j4GvjRW
/hC7u1kL+4eAYes4iABn2E4VbeGPgbD9OlKboHgHq4mj91uejr9fNZA49X4vejclfiJcayOrBcBy
H83cCmgyx8D86ny9GkUh64UhjD0davgNdPjX10WXmt8T00KRGQUEvOhWHcMTpBJ30N8/VAYeKTYv
u4SLLbwXNjm5EjgTEEULhsoGZyjCCwPOxA/IytBz45WSTcWeJ/4iHyZ4SuXliXTmyZ3S1Vqu27Vx
U9R2DZ8HPwPiSJ/PEhcAH3rlhAANBrESeMIeAd5nB3APgo8032fpNLgLa31KIAfG00xJoWwTkkCg
GjOfceykoLGPFCQwDiq8MaHLv9vOa4/P0VykZKgZ24iLsDuxp8V/5aFXLnvz3sGZoaGRptKNLbO/
gmkwO+DV6dGOfH3jyJYO9iosVLFKScHK2pjq97l0fDA+K7ws3ZfDm0gZm5/ObP+Sf6fdJSBqpii6
8WFtpEdg5cULnuXhT+3zztBZNLYucok/uo3CzMfWrEuy7evMRbbMOVxNkF3hv4gpuJ1M3iJEmsly
J2b0A1sZjj8iJ7ziXKJ8mAIiu36fhQvIWlBJLEBn8Zueaqq52yui/mD8T/pmGbPT+0peXVmoYKdn
NbkXX3paQ2toZYksa9iPZ5SLY6d0JwMcfkdPBP/g49smQI7neV4YwSQPJy3tauyNrd8CmC58UnLT
cnJs8M/cPmOouyfXs2ToBpZyDXXQAJUDDrJdRqwmnE3fp3MYchmdnJi9G3//YGwd5iGLYutwYPEF
TH7dFGd1Tc683qxMFdEVUNKO7rDtFr9V9DJfTwrwqyEZe1f3B3NeskC/bB/vgHz3IkIXqRgZq/LQ
2N2nfvQz6Pr1nDBXG4Kven5+beNAjVstHSSr3zEhvhG7YuGLKsq+bls64SGTZzWsYVb1ouBjZO3t
08h2/34FHgIWxTL4vE6amsDhTuk2a5XzoLgUz4t8sPSg7+mRuEKCIyDwDyhfpsD0sFUw3M2oBh7y
fgPt4tPw+AZhxyt98iQjc4zaYgn2PfFj5EleBeRXTYGGgcFUwcwYpl0n2X87Qjag91ZBvRPJcU5V
RMayLUdBPth6+oTUiwQRfFdrrAuPqryf2b5ntfN82BkolnSUmDGSNtLUeiQGxCqsLCcU5C8M+jHA
iUD55rY65om19fCLAtpJ13lJ8KKtKZHIhtnAXKQ8qw6yiETNnqGlrXC2yYzAoSBc7+S5XiIWo47S
GgvN4gdh1V9DCO8sH0VA6ShFxNI25QxMF5U5q2lDn/Wy0qJmotMjfDoU1qjx02vZzxbYyaFhE9w5
Cvrz2BBcSMpWssbTmOaMakb79mZeoysMR5laaJmD6GZf9ryzLfzdk8frXoWIg9sWnYsctqb7KM4x
6qbo5Njv7gqVXxE1YMq57x+HoUGipyjcpZ//xIxBFcWEdptJN3EpJBoid+cjFgv5fdkCD8p59qJn
gtJFKIRYfBmEge5e5MJyGKBVwUSoNJYLoMDiGx0MoZHZxQvS4s8KoxyLcdz+xaem9IlyATcZI9pM
CIhbAbnxfGBb2mfReV08TAar+iL6DQRI65oxiO7h5ZlBKlX7aXcMnU097xYMBJFhMLhTTbO26elq
+yTpqZRoeqOpTuoP4doMQz1pSOHLtKgPj49luMk7/kewHaUAzrrsqn8nmVWl4Nk1n1+msoeYqa1i
ChO0QoA7Q6IdEon/YRYQAhCIXK08EJPq9T1bvBz5h0T+H+hgO+gyJnOAQPYtCeUTZtMTg0VADNC1
4ZHgxmCfE6JwnUbZkqugd0XVUqY+SO59rzG8KervWIO/iL5Yj7bjO2gNBJiQco4MAgAQUsSp9VS2
HpW7uWdHpd7GR6K7vestuFDGxmo+RJv6c8w/xil9RCETOdCajDRLDeuSpXdxKyANok5Pb7rJXdFa
t0zp5I4axeIpps9MvUQSWvOFvpytLxUyx24Ia16CtTkJWDzhoIrkpyYtcpIrgcqOJIIRc2U2+4Wc
IGKOfVZ8wvrGieFdH9TK25bqDgEBs1WpkmTr+uAOPB1ZxpC/hEKgzhEA8nF5b/tDw3bfeHG/3Pgb
d3fPnq5x2R2Kn101aQbAksIPU+RzWsHpRqtcnyiq50elg8cwEneUoL8N1gKwiJMJ0r/r0/0GWEK9
28PrWXI6LXFahIS7RA163Zaf2c6WKsSvkOsYnKLR2yrWoFVQL+uOB/o2OaBqTbe+tPws1EZezHjw
m+axS+CWXZ2zlgnXd3ek1PlGJgjCd1can1PLI2RM9Uq1muhDf2A554pEHF+Dka5mav6Bfpijc+44
FHuJgw21dfaX3PvMQTFciMNneSaTcFKaLd+z1NGnDyJnp2kbTjO/OcXx/0ybZnJQLouzzwyrgBEi
iXYdf092kUOlifWIoZX3C+9RsU9hjJbu+kumHYd+lBEDaU+EigATWuBx5da+j0F/z7+SbyUx14Ki
JH7EdqkuILPDDTATbcnQb/o/qM1231hrbN22SzOPTwFjHP2lWw2BjWcdbiWCOIXA2CzZ1vMrY/NU
TtW5RDFIS8TuSeSQDUpmdp6OekJ9/MdXf633c+9+tOzjmIognXcGo0mxawTlo3d1BNE3AV4MzJqS
RDbdoM4ARYfyo09iUOFiHXB7vEvHOH+ZJoQPDCfYdGONDUJ7b2UV875cfc3HJ726anYU9MSq6ISY
Rl5snKFMkhW7Smx4+ZT81Sny0Hz1jJPh3ZH04StSuh0t1Wzkqq/IYkGz0QK6dRjYOBJphXYVGczq
5pfvivtBRIB6yQFi9JBha9Sas2Mm0w7Db9/dGpr+I8Tnl9DWuAnLxwgy7ADSOZdZ31N+aJPykeiw
RXjyrct/qj5f5/OX1Juk15/mtjIIZi4/qgZA0P3wLv85f14y9nwjSxhrZOsLcjeOr35D3N3q/NhV
oYe2pttzLV3wNwKBzDoVWbZBO9KoljewrEouNsHr7dAjpwMrnrT+Fx1qbw5eLoeSkBf5fFtgnWMQ
nBa3afSl6hv3M4xD5f7umzAIJf7Z0HBt3u1R5u7a4w+Xj17Z/ziVns2SnAZr2xADIeZBF501dsoa
j6azwxj0zm0x+o4pYGfD6JtXXHNkePBKGqHl1bHrO5LN8xw2FnWl/5noi9nFBn21pN18iYxGaj76
KJABPOmLYZGkc2E0JvdjHSrVP5VpRIfscFmDwWhfBSX84U/tjTjCGpMiPx4p5tKg/lndxQu7B3on
bQvaO5OEEf7C8uVMsMF3tbHw4JuXYgJPrUVGXLme1509nvwk+56yiLL7zPNCAfs0ASteETEVpVIG
Bcu5yxanuG03Gn8A6XTNU9rphEzzn8JosFWcFsQ2kJcXm7supJXL5p9qDQo8QOcdicJa2ggDODDs
2GuVkU25WvXEkDCAF9MvY+3hIGMoxeghpVRsMYDWzOUUUIpQgC+v5shNaCVKaTWXJsD/sFBg9ocY
YZr5xIHSmPPC0OQly5iR0nqvJuQUi1L87k/BSBO5VLNSL7Bl+oc1lwNaw1eSYGyq3FmCnpEdv1vH
nZ6SbOEEJYuYLdsHw12A2nhxP6NF70sOPs64vGLkr29QvDFTakrgBRy8Qm2JJ0wwWbeV+lKPD/ra
YzL8OylJTwU53Dnf6EfyUgunZ0T1VSJ4jSI9WRE2875gt6Pd6z2ZI1hla0Saug7mdqoZ/qlnw47M
IgGRnY3D/jmqiEzlbR03AI+ngATqXxjffeFTOR2kTiEjnMK4NaM5NRDZw1lhL+DoFocLC7ISmpJT
r6o1BNu9/pHZOqFK6Fpv5fRtPh6Db18lt4CJMRzuTvUuDJ4OMSa1EShItqv2kKKgRIqJzOk8Hhvg
T3OteJiphqgDRfoFrkMOYWcmqA9yLio0pM9UNrteNU44iUR9xzWHMwVE6y8wkm2clv3W1WYAWVjb
mylYPqmb+MfOd1lFrFVEpBUSDmOnf6AVlBl0Z62R1w7diyK6vyzdTSrT7IRz1g42eDX5NCGBQ05l
3jEy3SFp3YisYZxV8ZgXmJDWZx0es60nkjido8tPBu/qE8svVVyt1GvwWexw+GlPWB/BCBSkkLSt
MEFEKRvaWDtSgJD2NgPZi+ElMotH8Upf7Nw94Ce3bHI3ZkXq0OT4xi7t5p1hASqyz+XdbMIHlNLk
9PMnNIqbWwTsD7jJ7Wt5UK70lhdwhcLAFKBdoAqbih5L+lbMtdM1y+MUB9v+mB9PnYVfprcKIkW2
x2oNRA7z6J504ukNb3VXvMEQfi4OhXg2/5r0W26+bDCp2DK3wd6IVjJnOqmp3FmuZn7QV/JAn/5P
3lGcEnqJ5yDAeRcyHJi2z/1uSr9oKVms3KVAFSs71WS8N3JW1LmVeOKDd9dFLwlmo5XW+k+5sAOf
aqOKVROeeHz8q8FqiHJ0FZfEUA8GqmaMkcNmTBBb2OQD++sRok4lVsDYpE1W1XFKa5cs8usf4xKe
F8u4bZ/bTN4SQ3H3DLZ6U80BtAzSH369/CI8uqCcwGwDh6PBcAO+SPn74omLZlsc6l7eDQCc81wq
oL8pBKsW/KfXh/WJe3WIGHfHV4yJ6P9tN4znkstkeT0+mD1U+nROL2EIqKLB8eTEZZ5De90l4yc8
tAa/5IgQoxgtCAhuGQqZcI0j/N5pZgPPai5efvtXlmG4yGtRDsGgh/deRTGg6+jHd0kCI8yxv7o5
UT/TmIBUmjLr4TvgXUQYjJkFutIei2qv1wYMxGDeUNXImrksoZn/Y0Po/1wWwabPlBWzqYar1Vsa
geUXSSBA3CSbFxsbb0DDkzQv41qt/IjRKycidSg3yTHND8oaxV8hbeAVOeKWJjU7PIo6E84E4Q8+
xlJpbhf5EXrhRULJQ2I8mWvl1UImhEhOImiN4hoyu2SN+rX1pHeQ41IX794O6ysETMb7hbkKM56i
D6Ot99z1+Xwu/wyWDUIplgjPsDU110ayenyF6HkDiLm7zlXsztQlXu2XH4nYwpePDn3vMhbqqSUN
vIkRWLgpHBHTPufweyFqxxrIMcmfZJ56yQTHJgy6a4mmINzIqxGCLSvvHZP4mISU77Xk2XFDaCNw
x4HkCOuyJAlK7MP1C3bNxuOxl7frV0ofRgC/yghD2uw67777doa5eLFZ9cn6Xa2lDj3r/24omOXY
q5n9wVP7xN3u8BBavpC/AttifmmgBwI1iAlFbtGK0K3WJsDcHAf8uAEWocoIXCBFbqbgVGNZBxUd
jz7yzTrgFaWadK2mQKpBL+5KvUY2LoNDJL/CQNkV51TTaWWjm5F+LWzj7hsv6AATe294sILZGdp3
0SnQQN41LmQXgDYAIh2qNOxy+MdVsoyWJITuzl34fvQaGkRiPP91jZUPctkZNbGhUOQbV3xWHeMj
iaHzXqj8JNQMYk+kLFbZVHZJk6U/8O7rQ6WAY6FF+qG2Kc4If+LaRRySUZEUCkTuzZXCdsx0Tvk6
PUArlu50f9AHGM49a4dKoGrW+DWKVNLj3FjOzkjsHPmtoALJdmpEo2CDzkNIaWAgUr6Rf34iw06q
aF1xn0qDrQx8K01C7XyBpQXPLU0txnI7EEAe9gHBiwUEAqlK74rY+ER+AUfaVXxthm3oaP3t+MfQ
QutnOLeISD5L+qAmtdvvz4BTfYeEJC2acyBuwqkti7wwUziFQNW8Bu188MIA2Yu0SI8mF19bWvfZ
OsOJVY+3Cvm6iZCqK/7J1xB02lcKLzmpIQlNsql/46c4Pp18nlfGZjdGbBCSlOvvFrKNIVLKmafg
sygL3Rief03Uj2PYPWT07iA1rBVWTvqm5M841Dg6HgVqPOQSnPQ8JgUZP3VCBP56lhRs+VRFQqnA
oIbfRQ7vEpZpusFiIKqKEguLXXFhaL0cDBRRy8vF4HE8r4f5O0i9eY8LZ+fvvlK2ZCBQti7N2Q11
dFIZ10yDJAzZQWMKnpjk/1cdHX3A2fu56Gcn/+yFFJjQIroquEsiH7s+mQ0p84hCya/I16rS2Aes
W1szzhqV8a8fQbeOdiMllwSow6JveCnIvvaBjooS49k9+oVns6ljVHz7b7zQZhxRS+Dn7hK5Hq8V
AiZRS5ISZCSIPnp/oct4nqLYCSeUK85ypsbnCVYuvWc507dactIIY3XCjAOV6PqRwfC55d6i4wqK
vmISuWSIHw+9X+oDdcDS14HBIYkcTk2KrifDg/iUwUyUIg499WKgdujue/XBLc+RVr0PKL00ckGO
RB2DaMDaDKWznXEtL+ug7mNmbwuUm25/1AFk1Pivsj8jmg21Eg3K4slVylj4+K8Z7OE+mz8VAs3y
qtftUxXjTKygzBeYVwmh7owWBSELpy488LOCrEU6RfZxKtSkt8IRCTO5qKJYsOjYxnovMgAVrLM3
rdfV/Ud9EqdMbNYoDAl9AkFoqHXgWawjF8drtGUNxUMElK0bcu7G6Xpgs5NDGdFZyEWjKljihpO7
6+P17NgFVwC1+PwPXTy7yjqiJiyur+XamBojoHPa7Kx7J4EyAqFQzveVJ9coNUQHkkJlFf2vpe0j
KNfDx2LvQw9ANGwOKWJvDQ+Zb3jMl8C15IwpUGdCOx/8Qp2lsAjDX/6GmSI5xXOJNd2YliA3N/lP
PFwuBrl5/jqsutWvNhGHV3dY0xB79cQQZblSddNpjEqrzi2oLsHHaoGQKsJQeTWMtF9Td2mpT69x
dUNmrlsyW2yQzWGBkh40+5u8vct9t2kuC+YFfeMRjxclr7JQvd6A0mZ3+XHSdUoGsetRfnrsPmaE
fbOYKuuQhtzRsS6COaNfyTzBYoFAHlNtnNJ8gy/hcKFzrQiMqXxUjLgMGxzen50YdIniTAFa6gsr
O/71zxs36P/3TfcQeYvfNgctFowLS79RjROp7OaU7Ovb7v6HneVb4qUm6zoeoNm26H6Uw15MD4cc
kmXlZ6GnifmNM2L9tcCQkrIFcM0V9j43ceH6kWtNgtbeeReegkpouSaXawLDtxapDJIEy3f1RGmr
sdLw8Nw06h+QB2NAzFDPZzIvGwdS+Cd4LT/mfBXTje0+DCAFk71kINUolyNRXeBLOUsKWNh1tb0R
fWMa4xPZ5eb/rx93yD5cSW6CmAwAiUwVVLK2ZeQhn44uojjWwXAxwFIWHSD8vvVWi/ZZFHyKFSvi
prrSq2NV5qMAyBEtD7+6pammBKK+Cii3yh10MOabK9CFOyRR7IykMxZ17aUgWfMakPV3UXTeKBcm
h2a93bDqVHP9Rf+zM7OgRd/mJckKlNrebJrWbnS1zA8dRs9wRc+A1qJ2W2rmwiP92QrqOmDTEwdJ
U0QBJJggRo3bxw2idKiq/x7bK4fcWGbeh3MgUJLPVisB7MZvAlzLCm/Z7u1CHwu3CLXxHSxp4khj
lcspXCCRzZoNlP9GAqbw6u8CSKbEiM/G4MSdxuADGCOJ1slBEwNrQRQVFKEuRG4EsJ4q4hMLyaB9
t64AvRfhgMsAABbku4PmrfRNrC+/TXa49UKtoDkdlHX8sWzzAW1kt8lq8x2M2CK/W+OrfVQQkSzR
3pxpl3RCkQj3jSoVKsmOnrq4oc2GIMrbe0Ivot1shtcYgJUR8CUcQJOgdiycAdee1MRmUEA4o5qj
V9TANyee9sPcS7QqhFkkaRhvZH+j3B6ziUsYDRHur2YFJRrYFSEyDAeGolNVhW6NQTIkWgNNSNJo
/HfVWnhJtuvEvJUQJNjE4A8dCP0/d3dhkG8UQju8+3lNgrkEBlq3zV5UfY0/4yUfNVY9SEldDQYV
7DTn8ePSXJRrzrGfhZvoDGn9ZxmLIR4plgKw6m29c/fdXcmyIRn+m1A2UF86nLbDw/RJY6xjMyHB
7fIc5LT94+uct+eYcBNItQX/bCneh8LqFXxcmYbiuNPjZti1GGC9uti6U86oER9YaWf+1SWm1jjw
7tcIDzxniHQpOqef5IqaBWUi1q9KmBDwsyv7ebokgMHYrx7A1d/5Z0J4UTojw6aFZ4HeNd8WxUWU
cexGiWg/4nzSPaEi9zme6udqPG6NtGFDKwu1MZdx8T6+M/Hd/RS+zoZREXysPrzZqngo1iPn3NOq
A34nDu1oZGRlofo6LHLM78q95bzpAMduwokXv+ZrwAjrgM8+81ceguMoY4gTMmQtp6E6fEoNKEco
6GwGlZ3WbDmbidtj9HFpMJ5ihITJICX6HmOFOBDIulHz7j5aL8RKEbyfh1kQHb7AY3E5czHPVQ7z
iNhCGmD3R6mexPfGEyOAJX+kEjBaX3KrpMYf0cKFcuDqylqMrF2rMNyKENlFfoHWoOgxoZ+Cb9uT
Ns+U72r8Yap2A2BID4lsuD0rkwxtYsEaq/yJDSEhv6nqqyzvct7IeBcsx6bcB1qb4eCdohg/eWP9
qATBr2nVlK2S5HXa+NEkt1tk4n/1GANQvv5mW/DbzoHESCzT/zjEku5+plytDuB+GLyy4ysWN550
VRtyBwWiEwIs00bdww46f3kBXg9yKKH+IFjFFY/LBh0ivK5z1STK8pl5YtAo0UVJXrJ6P3Z6wzKB
JLXBJUVKQWWFtP0zTvwt+bUpCG3w2kbAZGfXdVXcFrSEe0yOniPpyavhyw8U4Xf45fv4pCuRN94x
8yS/GPSfRo4LdA+kTV+kg2vESxnY0cLmaWSrKCek1npysq/kOM5M+q1eSeN1LBF2hz5Bbb5KRvZT
ABz2umiKxI8gOb8Cll8aE9R31K42Ynh6aEgMF5wBHWOh3jgM6aY7j2S4vTTx7nEV8CHs8DM1TP5H
o9kE3bVVXy9iFS0D7vwtrTvTwPtqOREiD+/x1bsLrdty8ZX0YP9Aa86eaFO7zjho3KZw2iGDL/wx
MeNiNDp75bbvKb5euHPHGnsfEYr63NuzvQOtxYKhRbsDRkor37xS8V8FD8hBp8+HDrfXbKJQbNf2
dZep2jVtzo8bLuCPSSo4aijwVBTUxJQ74iXm9hjjvZoAGCmeE+rF+Z7peN+dfGd2QckKrDTtqy3D
FY+GOed7Tv73LhNECkC7uNro/h2d4qVGU5gyQj5g+Y2NAuEgNrsx0lnFVKefQ4lBST3QnouN3Gwl
5pI/hE1FAf3/++6f8Wo6oluUi3tmqq0d7Fbn/FzmVFhVX784NTnbDmplNmkdSoQpN54968YVBZ2p
+uAqbUOc1KsS1pt0JqtXdWi40HlUmSXyDinFvSzarTWhaS3vaQ0Xi/O5MF/NQeG4tqTMxflEQ8AM
0vQnc9jzLvihOGtR1Y9p/RraARttnmbUpzuBX551XvlVNld/kAK/3l9U3Nqvvce3Ou3gfAYFwyey
lkBw7Q5N3T2sCA9UhWLpNfYn01iHGooVDawvL3RopZ59ozY1vfV3cdLbAlxDIONzrZV3Vv638ZaM
9TffE8E2aO9puy7ibk9/QbcM6CnvXoSfypUFYFomNa1HHU2lCQ+D6+1pTKU0tnHun71zk4y8Ck+S
8li6Fvx8M1IZpeMQFyp3g/dIkrOTLZKEWWZpRWa8O/Rb4YRe5eU+Di9UgcoxjKNmKAfmGTz2Uzpn
eM7TUGnTbzPt79GpVImaxfKPxSUZBnvqT3qGb1Q89DOf2l2V3jXW33LDtsh7feT19yq47xvgnrU6
gD82WyfWgPo3+cJMaT/Y8aEBpp5ZRTiV5/piYjgqGwDzj8mgG/qt9tU4uiAV7N8OZ3RJ5vZpWGvK
txYmypZry7IUH+QSpgcynd+WsfxbUWzLRqXc+zsqHTmiBn7qn+UsjRPDfustn+ghMLPXuKJilaZW
dmRSx6NeRIhYwlqwSjXtaIKnkMrXfzQI94/tkdAddIeYCSfVQFZbsOjXOTKxaX8HXkAijIw2q6LB
kbMeu2tWSfVHbvsvzioOhHPRgKuIjbSbn79YjtOiMQOJRQNh9ZuUqGOv0gdloRkzQAlLtBy52C+W
VQfOQ40DXpHzGa7jLdQbdI3l3jK2W94EsNSCgW+UizZT7ctokCj4D5+cxDUvgnExRtmABcQCPrPB
Arcs7XeMjb4KmC1Y+PtOGr8xfOxJE/YQwLF40xP/RYPDknarCTmKNUfr0VQhVaFAb+CMasw6ucyA
Nu2HaXNe7GTRYqr6wEyW6/X3eccBBFeTQKkf0SEOLXBfH9mQz4vOtWKIUFrbLlOU3AEDxkiEl1pF
1N7oyN2pZUapHAsr5D6Ccx1rMSSHr0ddbQBLOpPWSnTDQ5om8+uXDOlncpv2tnscJNncg7QnfSZw
bW4gEmR/5YapSfyOouj8FUopJFjg9nQi4XQ09vaZEbCSpPpvJ3R+W+rE9bF+n5L8+YBPZKT0DMGe
KoAtd3JYfDtbwae+fKkQaY3hrS/sS9F/bbWqt2TSwdacJ/xeTs13Xuc4Uo8KO/oP6v/19jGjTK37
wxyWm0Kt/4HAvklqXe7rLubmmQu8AKnt9yv5Jdp/m7shPD+JJko7MTKXK3mr0sDmLFHGwNMGJyGW
2y/EBgBWhrUWTUAGa6x6k3eq69lrqaIKJyj7rra4FKlFAhWYU2cJ8skrwvzXz+mH75UMYQYeiS6B
2UvO2EgZdTQnjzLDxNCdUp43UlNiFVwi0vVINsx4DgfKO8DkN1XVu4Gq+fd7p8JWdxD2q5VJlD6H
7Bzy26cwErwozJw/FWyEjYcmE4FBkS+1LR6V/KDyBUfJJZCxcLHeiILKVsQ/KrhKRbW11J5fJTID
1T2xNSZA+0MfPOGkIk69U6DzC5ZetI6e8vEnc84SyZYCxW/eO1Whbrl+vn6KkD3b99cpNCzAd+oh
Z+i30stqr52hipcE/Uc3cFXtfn7i0qLLk1y90TTcxsBwvvQB4zds5HG4aEtdsQDW1NyvgQoLwzmL
lX3Xu1y5dN62tIJ16kot1kYA1m+aF4OKKmF7kKfFGsqKQLDDLGrgp64H9FCPqKUxt7sEdGtrASmW
w3DBD05al+Yn+uZ1mjesnM+tKKHJ3q1BRO9oE8IJctJzFZphY3NKKcAu1IBnRiLKwJWNwrGoeZoz
M+bF94XLTQWPuqmNHoXIpefu1W1Ir2TkJ1aCadakiUhSM7FjYyGYE4zwGNk4eySsR7s3qFg2XcjM
dw1vNyQaGxnu1MpVmrSod9kMiPPbrneJvvsSAgxKeEFGFC6bSy7m5bnjtmJ/Pp5qtmXkBBSdfZV5
2IQKrHiiOJgS/3uX84Uc3Il+7Rhn9eJV1S5aJ/wToyRyQnog8h2WrFrNhqWMxblZxlUb2eT5xiFz
oviGGPwbxawTBfgbOczsVxmUAtLEzALFTXwO4zESFalF3JMZRMf5dIxQjs8XjcCn7yasIT7VXYWL
uOsqv14+yWh56p2AxN+AK69QlMjmQVWV1MiGXjv9TfYbs04OM+jL5d9p63NCFFcEhuq41NDCYfNM
WicYc7QawKKG3WZlM+vE78rbp+gtfiJTjPS50dMrj5ut+7dCeXF7r3g3wiIosCY3fyaRKxk4hsCW
aupVXdRFpw7V/UyWzqu8BXEf4jBpLn/doyVQVhxYibt2VdX0seM9PXbB+7OQ8sWqTSK0aUs6w+4I
yUZdrCs+Slq5yZWFOeKMUm+a0qgsXAiJuelHbi5sOdRIUd6VNvuTJd7NxX3+7gGbZOFhdLd362kz
edluoE1M/dMGrS43zVo7QuQnDYRULp3DOWTf3SEG3cunF/HWUqnlrmWkAsHzxlwIyo396XzlE4hT
w9UuscS0vtnhTjMSsVmN3RxgwFt5taL3//0LkFavQ1rDNfI8xEg6IAKoFUku+mXOs61WKi0E/5+e
w/EJjmON9rGcC/0CwhEfmv5o+bHd/farIop6/9i21yrhz2RZSasRr64YaY/LSbpVH9LM9Bw+mRYk
uN8d9d6tHtT0EF213MlWBIqbvlCEz5x10kW4UvLfD04NTkpJlcg6Xb4Ak5A19MSbGKyxWBOxW4JO
k8MDGCE7nabRUBX0oAL5/Dvtn76ogcJcnQ3iOCYx0F4hxzsXYM+ZiIzrwyWdApX8wkvikp/ozMIl
Qkpaog+jRsUUHPH7w6hUx1A5yImcvkpcxd3eNYvlBDJD57Y6lt1A7AOv/kFYmf6Wkj+GOemmcHmV
TzHQK1duvz8qaxrjjD6O66Xh1lKgSLYAb01AmcqSLOQSPJtrvYFGCMMWYDmHCr6UCscJnPHVEJ22
FAXyP1qGxR/9BINaH40YK8R/kRIvCVwNJAOK2UbPyOwoehR1aKiYmt2WRTy2D5gwc9sHC30I9D0t
ocYjkOFPdaqimV4SwsxOy2vFPG/ktCgmWGGHsdIjP5RmkVKb+9MCFDK05ch9VlH5nxJvNCYAH/cr
t7KJXy8YIxciKLAzA08RgVIE9wASo7PXfJ9Z+Dve+cKfsdXWCbLwR4QPYHVu39+vizBJTgLrK3pw
HHTSn2JS/uFCYaUFOUc3NNhL1tZiE3MJWpfvnNkc75jf3zo+QNgd2gSuuG202HvG2i8m7FmuiNtY
5BnXyt75wuj6vc2arWQH7No0LkhVMpgY1ElPJmb5ntv11KFX60oMA/Am6HpnwdT5Gcrljl6WJ2qB
pxvnIGQT3KJqnhfbpQ8hLoYxbDLeTwwwRiLNZkNvbEty13bc9fCnBjoC88dWlxPx4ZMVppi/R4BU
XPFHwzTVyLgyzj7rr4SpFCre2eWY6Ed5zgENrnpfwGIbspWUK35LrZjQfe4Vis+kk4WjZIXAHT1Y
BgpVc5YGNG4vf8SHXdmituX3DEJOmcua7qHYbKoc+GOCXML6+l3R2GauWoR9Ir2ovn2PMr2AQGpZ
ERFooA9yKVbPDC7pi4RITeIIEKtEeqECDmiNigVldI3Zlz0/lHaoqxPJBnJjXaE4ea8a8Z5AgaLt
pXawCgYFBONtkSUCXkeGvmg37rlea6URInzybyxFilOf3Q46QiZgDeM0DagHRnER+fHWHh/hNx0e
x66jDPNZv116cechV3tGEhimWDVLPTrA+UkAeQ3Ncv4z6zn6/3lj9WI7zG2z9o+yUYBYb2uokP66
8T4hZQzxQI3inP0lz+jiTl9xGchMYAS0jWi2+zHWFc8K9d1+Q8DJFhiIoBANxupX3UvBcU1F1A7G
yfhZvSJfy3NSA3FvLx+joqSFtVaEmeWqYL4jTggjKgjcoyDfe7ISJ9LZs87xeTbl9gksVKytGMv1
DIuJj8ZVhn5BhN3BNV9gmLyHc29jbJar/KixNPFROTpOBpnlLobENYXeDYN0KEyQE8f4/p3lKZoA
Bzvt/Q8IpP0dIKzGdGTvQw9OcDLO819Pfkq9vBfokjkJts6paqTjBeBJnponMeQXpUcAkouZdRNt
3Cx1Xgafw4CoxM0k5jxBq3rj0Oep7YeYyAJxqO9fhtMZ+esUsJAKPTv/iuFJOQcnIBXYFKmV5zqW
/1qZSLmyQJSYWdWRvJP3MpAWKpmHc6mr/lMa+wO1Bugs9m+zCr1UcTWXRKu1KShbUfSD3IMynD37
nJlp883wxZi1PomAXrK2cr3BM6XpzAwBsctgLfdZG2oaq5CTTuz4AaFbSgwTRE49hXhdwnCftglk
ZqsCUA359W3+SHb9bMm29oRVLffTywsXUtpASg+OPiiu6Cfo4ZI4nEKdSd8z4Jq1WPy2cSqzSDbB
hJnPpgunmadMU2OEhtAj3ZdrbX8GgbRjt0HukP5xCh2bOnp9t9zHReeFdGqtys3ZWscehne9f/z6
tMXCDGwkK/vQnGkVtS7xFD38NTVyz5lopNPTbeilsoXk2mdKKtOQGZUYgrF7dhmvyIxSwHleOyLk
rPtBujBnUzaZ50R0oWIJcjAHgLS7/JxPFgx+oej/PfrEN6ylHl/ZJnIwwNlvsAA9/5OUb1eqRmqF
6wTMQe6RqPk653mXaPUFPBe4C6/AOESuXndsDw0tHGImnvVcguehRrF5m5yU7ThbXfJrTuqin2+I
VX3XtgwsVBkRDF7BhOu+FGIj2HPP7cAXa9KN+hAQFjPDd9GpI8iGutcrYYPHlNmYN0p5F3SmaYTR
RCeEMOYmrBk0fp8m6/eqZgl13Rqe5cxoNJvd/vC2Ch4rZTpeh9s+XYdLXsQtC7rT5NwagHiwR/3D
+yCLSKToa0dxJzv5BiisKgzEkur4dnanAfLcZyKldVsXss9OJqbhbvmecBpJWzy6LJdX7n3GtkjP
DfYm/oQ43jfJ+Gnxi1nSpSh2gtsgloBykyzdWsy2yGa16DBquI1/2bucshEjWwH4yaHplAjXdiVE
3VHPVluaRU44aUPnfUEJJX/NpgL6AcrZ2c7K3hTxEN26l8kUoAqaQOM5xN8ryJHpn3sqAuxZX/+k
Flk9xo3OId5mtC9FlN7f+QNxp6Jr7z9yCLabjFdjo34maDhMXf2iZOwrbf00jWn/W5TN4eHGLsob
VhUHmzA1MgT6XI1jeef4Yq2quiisadlZ29Oca2r9PzjRN0Q01ZqNM207STrXWLKuv9X8CqXcfWCF
667djQN6tbM8GiShnEnpc74r/a2HjKHCpSFACqYJrehZykcDLjiahCe8yKNsxrLV6QGBMvw4wO5l
U366MK3j1nVnATIY/r8+VsNYYedVKadU2QRx/MtnYPSqI2bRmpKnsPzBJuGdf1dwOf/7a5u+mZK/
www1afeRi4ezBMa7Fm8zJxIGMxDgpsulaCoBXlulVU/3Kygfm0sAlANtfAqWPc6o9Q7CsY6bBNiz
WaP7eRVwrejHN0m7Qxu2lwcrllR6ntKCTT0aVvpNDdhQSAGzVk2JLvRpi0pBa2Gv0N7q6EiJeYhS
v1EF4eMdpAY0BhioiicSHm9MufeTrWnBafVeW5XOsgsD5mCwjigXCUEtOLwynSmXHAGkg7csOUnh
q0TPKlWoxN6XaPYCvZaUpEmoo/qxz3zd+dBhiFZlHlkKCaYzHylkyr8XYZnVT/MKnZX/ZRhvbKOK
Dg4z2EFFLCBGG+ghukg+x/K1uYj/KIdcCUmpC/qjs6PnsUMx91HG01nLn051T5eezfeapvuV6j8u
tz2KySnmHuhIDRnesnkYoqUGv2juIrMC6+ev/qzbGHK8XHgQDHf/BwzKfH9I/y2/o0ffS/HgYDut
qjiqXNmURpQnwNoO4EwDuVopGH6on22eiTvY4uwoFSH34mKCi72I4OmMzZX+c8Z1UAD+k1Le1354
jcSL2jp8UuU2sYxMU4XLi3HPmMdh7jmula2yPLLGlqCdBuVXYLV3ZRDSPIPfWDZpXvGzpuU/2QSe
dbrulJnAtX1yqcy+2BbxC47n3ksk+awWRzsBimoUeySde1PZSY0b6muIm1/Ie82IX1D0/HjzLgRC
66i5FBlQPLQKSrPeyZqtCixWy+XjqT+B27tByQMux+QB8gaSH2i0TpMFvb0oq+3h4opf+3sGpr6l
LGyLP0v2jVdxdhfl4rZjvPzY0T2B2VCf64pbQnPHc74Tmflsk0IoJ1TUg+oGqrKqZKqdUlAON2i8
H2zvvd6iRQVNxFz7Eveqngy//nTwqdV7/gq3AzEr4wYnUGW1jMw+DCE9QIuzLIFHkD0xVt0J6Vp/
wjjh0Ag06a2HSl7YmBEFyaQxdYuEx6bZD3AYSuhGF3ZRUJBxQasEfd701yr+0OmYsWMAh9adsAT2
Q+WCb0OPFGc6727jPWWGvxKLMMzb1E0+rc1WqfHp4PcB1+ESQR0SO9iCSH4a1OAVGffjwVujwWss
/IIDCsVz4WQkYROZxaTmeYZ97700T7nP5WZSzg/8fP3LTw9L51flPo2LSPHHpbR1N9IiRVEs5YOU
tN7N6lkAPGOSuIP4oEqNXyu9hfh9XjVtrLaf1gwoEHiVo9spqnZ4WDASSxydoyvja2Mz/Iv+gg2T
gjdLjdkQqVDQz+ruVs4Cd9i6t2Qx4gJNbcF0UGeVefPtScGK0T8phIdt3S2YnSVX3we1bSuCMegF
ht7QL8zVL53ZrO0+rczc4mAi9TXlzGG7nAhZB89N4bTHI8khvA8GzRmFCq/uICGFx1T7UdZQj0YP
pWclWtTnwtJ41XYetSTJMxpBn4bN3BN2B6nCMD1TXeSZXwA/diqXFMeThhEv6HVg5lCW9b7jFfHq
yLWlSdv+FyoxE9WpyPe4ISdxE5+VissLyXH2ZNOGSqzY43IWIE6/tDlQfUX24I6WFU3wow5lQBTP
dYzd0hk5hqhdckkgv/7HUXFZ6gNC5+5FlW/td2JqRPcr4HYBmehSMFmJoNcEP6rP8DOzDZEU0KPU
AEM9jDU0chIqRc12cDxlaPsxeruOjSqmmmW+zWkoxB78mCpBad34xlJsEAU4gqj0WkTghyfV7v1V
glkFGtdvpEUyZ2enbQVZXV0r3YOQXmtIqIh7NGbO90RE8whcQxTclffX0wV25RSCnb/K1Mk6bfer
bSf1+FHPL/4/z1A808pMMof1BryfCyyY5keKYha58trxlYIqj/PS+JHeqPRoz+fd2VmcGNzywby1
HC+Lt7XWBHJsevKNWJ0kkLP9pNH/htzZ1KjTtYGrErjUQ2cDA/U9yqp34J+MRp5JAZixhtteXPbQ
TEaPkvzFwzxl4xxxNoqBv/S6Dja0LV73dov6s7evgxuX57/CflTpP7jKbHZ5CB8yGwCDFSNMSqni
LJCLkwbAIwGdCh0X7SsaZqnfu/bCIE6qqZ7VwXh29nQC7GV7QVx/DeMPPqaknNETcN4nc0A0ufX7
EFbJbQGTwTyIBK7qJw7UV7a7nxtanptu8hRNjWdPTgfnBsDj0UcH41WT8Q/WPCvhW0450Zj6aQLW
/TF5TySILZK0xhEI6xKKcgx/uFBANtCQD7+DQJv7D++yRSfHPOeb7/2ZQZ1BBXNn7rEpRcyLUohE
5vkIlRcVKM3XfAU7R0Yp5/KFK7AGS5cIjK6DZakyF+W8CSc6C+pQ7uXwQeuJDUGL465Ax4F3rJwo
6Eb4n/G3noNGlFzK1gl25dUixVTe9v2tzaW9usQuwtNUGwZj/qHHIZSjyBSqURjovZpOLNHtx0YU
Hs6kID6kmPs/uu0W/1z5yqLp+8q++JVmCjLEKC2PBXsDOxK0hKsmuieXOuMw6NDtFRPr0qYtxxwM
rNFv2mxY9gx6askN0SDvASKSMQdiLjOxFpXc2qRTBBh0Lmf67FSfgKJLgOQd3SncnUcDHx/cd5/I
VScJgiSzK2rS76p1a7ZHEzXzwKleeQxx4DXnBcELuPa8I+/z0JHOYhyTCjFIb56oio/z5XethEzi
FvfD4yYJx32+osS7jrKnEvWBlVourWyKNEfTnVVduyQrMpvXAwAkh+WXDjQa2tWgJQCjOrBXJi/7
DHIxQS0xJM1RH9GISQNclutY4+4y04rt5HzcFu8xKuV1gMVBZE3PfQRVlB6RioWfXtu9RWCeFMGx
Mh3DjZhIbfImvnrYJ10pdOIgRir/XpCbwZlcrxh0M0tSj1Y/jhvpTwPd5KlqAYrEDpiNzK1YJ+Vc
dsZ/6nV86TxKdc8CQsHDxkXVlHvfoyaAbZA6mKn4SID9BLJOp+IllpfbOQH2Y2acfiBS74wDjqHi
H5W9axsgjFN6EbOYlgpfUhmgqpDUHaDIakPfQQubeus3B1q9WPE61rduZkiJBBX4W3UpR3CiLY5Q
LUtkazi8gCr/ytjPHHeIfuKdifL8lYCYfI/w7p6HTZdtmHaJqENjOQ/p5yhjSNTLcgCL5GDNepZl
EG8+vIrxv3we6abY4XeH9MjqVUr8QXkMXKB9Pw/oWz41XCVcans9YCVHBN2M8k8hM5SlHQf13tUC
KWfC+gh/nKwt9OBoRLJl5ulkbwA5A4dYRtuVlnQt67o59zmkbCOrqansEU6lhw729lCw9JoajLOg
85nMKD5xWFeU+X4hbkfsvfXdulCLyu00GsdULpXHVgqeDgIvLUGmYGb+OHihwMs3PksISS6oeuT7
NjtPKLwvDtkUEIacbIHmXgmohlZ7QnZ4B3YQwcwj5HueZTRLSyA5cFypFM69E1Xu0O2+4G5G3Iyl
vyHtPnbqmniChIGkG5PmWZI6fEDgWKJJspA4HnLvOF6fAKt1kGLQvhenQyN5xcr5xa2F5l3fJaB9
Do6VtdHAQ+e5/AE2V3TwQpxGuQGUqA6+sr2uQIwJkg81rjeAuT55EdV4HZtU/VMlWAE31Yhu4pcG
e6MO+WfLLAOTqqJlCKFSRnihhdku5KhWQo5gHFkwzpWOJIISjwLlIhJFbaIOGEgsAJbuH2pUGe8F
o41Fx03t/nyJ5h0hnjtY741xAXtHVJN3IWu6XU38I5aJ011KQTVzU/BGsQ1k7m4itgSOD31UvOPc
SmsrmzwLEs9X97Ncupfn+jbuavvITAHfwOP4Px9nhpxWd6M1943k8TzBMm4DuW8FilPlQ4eO4Ykg
pztiC3mm2FCy5v55hv2vgq7K7QgWahmNtQ522IR1Vtk2UpTttx/r84+ysgA2DOYBBo0gOQImd2I9
obvGoSUQvbqj3nMv3jdKED8kQij5CRYQKS58W/IMebuTjcRlWvu5Rt7ASG7y1xUpejZn9IkU4UJi
OHtok7Q7pZTRrM0AiOiuzqDeisWuW2qsb6RbmvkPngCLqEn0/PEyIibN4qWsyXTO36ZQ5XMiXhjm
Saw+oxqSH17bVrduz3eQFOMVazDaIhx4P0gVU1f7BvQ2seZ7v3damVak8d1Xr1FYDp0iP700gjf7
f5hB5hW/eSm4YDgLpDwvmAzXE2KM5REoNMrYiX8s85njG7mrRtaFgzd8daDBY4ipr/03RmmGfIm4
Ul/NsMhi0iiPbRlbpzqWEAGt+heoxYarmVJzrjD2zSxV4mvRcSGamxJBjgtUzFTa9C8ItHzevPpA
sRf9BLbHTU9RJz+C3icogc24BOQdF1VbyOyJEq8gDE1m4HNStCELDsfqBuSzKkOJDjbHTVrBVwuq
i9UQGQ6PzfYkkXhn33yxgD91Lz6GUbOPoH6iy65LrEa/apBnXcJzti5a7Z3wQDNgL1U5uqjx1Hfj
X2dyGckXR21rG9MKFPjCRhfELtkmm44srTEZ/e0g3AC11ggoXamorN8CquyWjNhgv3jdXlUWuN0F
bW8jSO28El9R3Htyg11yh3R9XjOpEKDVCLDroWzYKr4OVwCAVyjWvLQxFqG2CJVyHcHuluSBXJwy
boMIuYWN+oKHEtwuo3Wuj2VTwnxLPbWWl+6+aZCowzd+fjwix2/E19oyAReQ6ltIXDm0I4fB5pku
uElyDRjdgnlMK7eS7um4F2MWSqQkEv6PCP0yIBlkSrbtZi0stgraOhJjYEshATAV4GE60AepaqzI
l7QmVPm/PEdLZ+w8RsGqhucTt8RWwLYa5i8vOfX+5D9NzXonlMozI15cEgclQq5IzXjcOfcba4H5
rLhTfB2XYhSSi9H5iTo6nxSij4J+yHfNOLx8oeVuJEgbAZBd9hDCKYkqwiWZ0kJg1g7AwIjuA1Rl
105kFGVR5TKjhiWW9sIUqQigGOuFJLqbwE3Y3NcYdYAdCivzOvJKHIPqIfFtYkZtdFOjzbPXPJ5k
V1+u/bILZ8JC6HequAF98Gc66V/HdTx0yrFrLMqKKs1O5zWDC8flkpkPUiXn3YDkVV6Ni6M0h9sR
RinP/fbgqEufF6h7HU/ycg5+xa7zO/DYVPML8V0fpi0lnke7CW46NSa3JGm6/lpiNVwlBDyxwJg6
BASlYnxJjQ4Fsh5qFQjwPfCLZmEecaioryLsZ/sSjYsdvgT/4sGvKTu5et5f85CSfz5fBHnAojtT
8tEBRDgtqIMLbk+77PEzGTI06K3zEvKWDliWH6bQUPoMQfPgB3dcSdcZ3OXSUo99wgJ3rC3WnhR0
bmmSlMfHK4mh9G0+NqWePUuQ2Na0J4/REq4QUVIJHvoHSkZMhxb5jomd8qw4i5gRf1JEpBJo20a/
4sY8lF5mDNuP4KT7iilS0hjWDJ3xXQAzvJhjnFHyoBARBNCZTCOoQVHCAlmdbtchjSm+e0N8iedP
oeKPEdgRGuxTwLSwR8rgd/j8+itj/1DpiCyShop8vOkOWknzflTUHaI9TH+DCSZPbozoIbKlOY+T
dNh0PJU2qEuvXbkXFTd603gVsB988oKJw8up7xL/RgtW861ebuBYZE4aLTYp5psuzDyA2cf9PQYX
lYboL7z3IbP2Obm+RlJQzGzjkvlRZV1X3S/qIX7I0phLXQ1FKjecBYIYGwXJERWU+MxWFMLP1l5m
n1uaf8nkiVn2DUqPL1GPZ9a297bfp7S9WsozIs2o7EZ3+3BtivuTTlFAvwTLGIfQwgf12GdI9AA+
JqjUmdvoyIJxMILyVhTg/2gZ5BzoIiX4UzPlFYgveOWn5hDRqpUMK3bChRFmf+SbsCJLacZwb2ay
JUZyysK+ak06QCoOghMo4z3kEGsY/GBxLX3fNIz2LQcKyvr6ioPCNRBrdFMxOblvvtp9DVGTRDpO
Jlq2C+hFUi9fGfxxve6YFquiPVnjyM8EwA4y5tztDYJyu+HilAVqJBD4SOhW2AA/VMb1Ynjp3cOD
umRu3xBJE3VruWCn9o46B825NX6uEQcsBBFjy+pYYLZDDHfgVVFzyx0KgLg6eRgpQMfpKWhC6VmZ
vGGRMhW9i1zpdF3r2RPqSu3YXNas7vtqKxQAjWAHXeir273aW0VUISEvVTToLZj5kfxiwYSx8ycw
9yf+SXqiltSptHNiCG4n9VnBN0t3j6A9vTtk6doWUQgV8XVzdsMvq/rwk4TxvcLIk4JCJCe6/A2h
CEycJ86hiyiyrpCRm8NPGT0j5bB1enSe4kx/vQ5G+IChnsuRZldcHScCc6bDK7V578MVDB39B4kD
irQ/YWC0ouhkYzPudtfC3jS7upnOvvuB4NtEPxZtgiZrCtHO+KSw+9OZt+0a84iET6l+x97M2pGt
YSWgVDxhJyyWmW36kF6bm/mYEJ7nWRoTiQFNo0incgp2F11P0xWrqwwOC2S9ok8HcCmVaQ4BMgz6
9exV9ndIPhIaKf4xB98MrchChP7g5h7sqKsdnSO3OVBuRYT57QahJlyg09SN7JqMN6pjl4MPEIRi
/UPHmkfpsMkwuTx983Bwgk00A7jsIz2eLxMC8gMXJsFdnW1osFK3pZRgHQrart0XmrYUUN7XxXmR
H+9mWsRZiXpfqlc7zBAaR3Khfd8/XnPncmQ41jcQ/BScBJWE8qkGRX3iOHnYpbtKjaHD35mURpgt
2EuwccxG9Kfi+MpBH4YpZacHhUKT+iffmPZgau1qnf0Fch2AOIemOFFik/ceq6ic7EAT5NePPIml
NEAQvDobUVxQYkULzoMazuYV5lSfdBtJAFTcn6l4p5MCDPP0ba799/M4/UemPzC5H4uyHDMOfFsQ
Bi2WVovtB+GsJRxrRS0X1P5gVWuGaS2GoCNs36o2/9grW08HsZluPZ+1nKONilBmtM5fWh88x2D8
xUsU/AJzNl+oFoPno4OuI7JRfrAP1uCMqMwWY2t2TBcq8djr2vyVlxnTmp652E1VqiJUsIz58L2W
ZL0d0ntGRnoNy1Ks3APYO2vFhbT9ZwchlxSXhTRlkEajMOk9W2FCM+cOE2Smy1qtgy8yx9GYzu1o
LyBJuLvJCi3pa8NjI3FNrJSeNBNVsZkMGQfqUwJNMKTY2sRp2Pb/OMs347xtWGfJ7mH0hrFyD8Fi
f/3N0arGk8/YDF8iFgzyqt8bL5Yz2xlZcUjlP7nS6mlihh5lq4M+zBeUs0mnfXXXDgh47ekjxHD1
mafXjxn0qhEW1uQC7iHAiNQjUoM8qqvIGA9yD2RU0/RxCwZirBZydZ2MVYCC8UrAcnbZ+WCaYGFD
PDRkKzQP/ntDgMVyI7ZGKkmJu3V4wnIZhiYX30z6rXRevp6pVCwBa6mg/H2ixyPukgzHI4GCGHWN
/ehm9dhdMeH7r5BpVl1Uc1EPWcGUDQ9CiVNK2dmfr+gi0KkyZPhOwqNhaONAZ8aNuUXk/Ko/Ija9
5Ac0b5Ci3+G7BmzCC7ZtCVG8+ju4iRtdN8zbnVLKhPubywtzlf4+dUhTfKtf3cj0SIa1t6h9okpF
hV7ZIzysIeD4BL9zT2PrrL+2CeYt1dVDDTjLobfbAoeFugMxQZcEOx8dLRrfvTKx44PsV5UnetTw
86dM+ZxFbSBYHKCuLHA7EyFh9zz9FSVO65G3HOAUPm5NU6owEg1DHpJmdl6smY5eO1gz7fJmTc/C
7jK16qc4Ta0+jEFVXeKLl+AAvJ2LuDpV5sTerdp0eNNsJ9Zi4asWRJLSqXFnicmjnanopmtTGDSv
Aq07rtR8KRN1zA/Dpc9SctNToZoH8E9bi9EACJv1a4KX7rpOcwyMWeEDQZNMkTE8I61DHUeV6QWM
ATkA/2W6c4ApQ13P3wZAsAMuLvO1wrILE+0U3sy6JRBrjzuxdBLUJV4ZKcjo6TqkcNLP2cOAuUqj
JmjQidu5AqxWEpV1z7ai1YHRhDMfBaMEEU15024BL9g8PS5DeQyuIhvJScB5cp1vemNoYJUQlDLu
OkxueSZpq8U5iUdCkriel+exUWvM0rgy19r8ljz5462RXz8+/Yll1URP3vOBdHxvaovea+J1FTGF
WEuXxSnvox4HCEJr4EW6+elK9dllAAk8aqx2Ufm+fCSVlY3wdlTmewNLUKAKZdz0Gle0XynTWH4r
5nshDNu/K4xj15nGkm0pUl2bVn9ssVwIl0rIFfsJ+A52GaNHw2LKWo0OThGf5zjHqCA1evYfPtfK
zqOWy+IlWcUMF3xHzXftPJmQ5nDvThhk2xnFq/GyXcGVRF+dMZahOv/EYq6s3kZqXcUpqjOx5fGM
QPWCwW41kjXG7wIgqeOc8NdZGHR+yYKk72QOtfGHVUzYeP7y1WqsMSM6JwI8DOtI2zEsj37Ykl4Y
E3XoDFpDW6L4fo0JRD/vrMbvL2FhuxFxXP9ecj70re7ZM0omQ4u24f9X00spncpnyr8toYbCjUj3
nPlmjW9DpQ2pJ1PuqlU1wv4Zapip3gUeU6K4FfIRXY3ZPtut9obDdvzYChrOqgQC7OeQRpubm8ri
la0s7jWeoB12+yaih3waRD5rkw39oz73rmgH5WrN8z7asep6C+CYtmGD1J7nsCwC39zo1dKsZjNH
AtADjPeJFP9HYxpO5PQs6nNhA4gkqfNFxhXMGQ4p2dTN79EOnsDH71rCrEqqCXaEtq4Ujnn4IjVI
PxYZLO2IbtFjMy1Sip6TuUXZWya6XnVj8ym0ZA3vv6JWI0p1ukeuOs4nu573gf602nCTbkHjEZLm
/B/owg9WUbKl3xubuzJ+u7KcVlORXOwsQawJwgiEZZSPUcSVVRDcPQwE42ZT9vGKhZpXR9SULjm0
3rmUMBG3NlFblqnc8p8g5lMJzm8//ISu5WXpxarGeNV17dGRadWwAIFXuLsEeUqjREbeIyKJ94mc
/zPbn/Q/iqsunvRb7fUPUNBQ92BSj60J00kaIl8GR/a66zsHWRpc6dO+s2hEbIavt4AIY8LQjO/B
nlOXxaqkr0Vng3qfoYmbulQQ8lfAZVQiKVzG9kEwtUkddg+jOIMUOtHwCpy1wIRZ/0F/SlutDFNi
i/h32Czp2VqEaP+CgDd+0HjefPg3seJkAphAcTq0gYXfWb7aqNxGGKwgfhxDqjDbC5AxEHid+YYf
Jkf8e1ijxta/6iCUJBG4Br1lEnwmF0swHr+KiblQGiS8YTc9hLRt8o1InKSKToxTmhZxPD4OVjDI
2Va2FUAwTUzQZJtJyqbSuYS3TZpxiex8oN70zhcwUPgAnPQ3W/kciHc3L+d+dmM+8dv6vmcTKuc0
s6RB4AQiJAFfIGc4mfUyAWW9TacX2cV9l3ELWWk4K2UJEx6fkULMyTwpu3Gsi5r6TA/EqARIX0Ax
kaxg78qR9RATevt+hbx8dI5iuz0Nd+vavpi0xgAJ3FLkJaB72RudVLpwsn2ivNpcn/m+pD26Ol1r
GwT5BSw/4DfelTj80j88hDwghm3vflXvxMthfj/OHfgxOc913XWiYDshoqFXjk9j6nkXCHjjXHoO
R7MX9Znth9HyF9dyLEAJzoHUl7FsHtlHch0uJeVtNZ4fBE2Y0+kfHHxPPndlJtYzFUQRk4VtCX7S
ks23dSJPG+7b82lA+9jtFHY+w3oLpH84ROJ/RVAfgueXrtYmJPTXMtAdqtZmm87+zjrM2u/PD62a
nb+6/K8djlhtV5pCLenlCTB9KFilG/SbMk+ebZG1wWTnyYo+xygYuCV3d9D1x/0NfuhpO07jU4vO
x4QydJpoDx2hhiuRHzGcJN2UBuv4s6H9rmA2kMNPy21ugF2BV13DWZMQMxMWtJVOScp+AIhTYhkU
KYjdJ6C8SDpZRDnNlEwLRqe1UAEVkeQ5jMsXnitvd4NVIoNzzWZneGhOH4zjcY2VbFBT5AeQ/O2R
4+LbVYyOLNzlB6KV40jL4Rpw6YTeL6Tk+Q1dc6l0A4kZNlH5LdYC5uUAB1sp7TgUUZDcXVybbO9e
Zdmp2CuMJoUpy57LjpPgOwMVDfkjyQAII+wJrm7tgzZUuI3k3cymnqLwh46FD8tos5ZUBb5v+/DV
QA6KQXd+wUaElEmmp9VRrhdyFshMnfUl/OwCPuFNHrIMxsRRu4J6U1OYdAOqxACdUQoKpBkCK2O9
2AaklKJcv6NuND7H2ljK7AnuDp0Afdvs/vAmZyjRnGI/EZ1chAR1292giPrLlbwhQy1XYLJa7AUA
rOQTZYpKQUItrhGIyGUmKEx3bfdk6A0vgBYLzorxR6176Oim5hkO9p0TjWqeZ6eARf66wIcyA4Oc
RfjUBJHSV1NbTGk/DpmEZqWZatslnM7tbaFBHwrPYvCwECMn7fQLq8eQa1fsT+jPxpoZ0VBFWsye
rGhJ6rOBwn0wkpQM2fnWnVSF4YnkBsWvAZnatEMGDaOtnjuJZebeJ/vGFkfmd64ZaoVgEaKIwSZJ
iwTbjnVyeFIVa9QpAcBiargsfoHhkfNVlMW7oaLXTP20NtwLWf1w/kmOJIXV+eh9T9aqtTI48fQU
uvYP0loCzN2MSpXVZs6AQoKvJk+0/Xx+wNzMR7GDAaxMeyMsQD1CUqzUIQ+YGTEa66lrH5lqvKI0
0mrMe1zIaz5NocC5FyG9Z8+9U5ACvZahK7xvRjVLEp2Y8ib5IC5v1aUEXWedouu2/VwnduUtceGK
L/8tJAOqkd4UW+WnShhqE4l6Mo+tAa9PD1h4A2PqYWImrUvsUZnYHEylFkWE6Xi295lE3RP4qXzZ
T8EYHhKbs01WZp+OpU+mJs+yhptUscCk1vw0RUK5qLveXJ1O14Z95mdKPXgl/WlJQ0bfkfFoKn1r
mpKxyB3EJIfYzJAlnzhBAUwomVPw1+qilWscU4jWKaEthT2A+QFCuf7BhVJ4zLnEoMsCdEhKUb6H
w3X0+oEjyUxeqbOZlz3mJHMOGZGSWBrt7S0Grw5vP7cbMfJGckp1JSU8ZTSIRrNuFnwitRWr2M26
MpJmlpACp7x6yNKmz5jukWTepoi//jW+n0X3bT+YpwJw1lm6uK938fPdMtBLQGZp11OnXIrfdDkI
voJxytRVe5WREYAHOJTTmZ+V1p2uT8kqzkz8+asB+opIPq4rgLFuAY1SogLS0SdCkTbVT7tph0uL
B+SHqZyXP1KRHkboWXhj4tauQoG4SuMOS4LwThHGvw4BlhF0YIR0L+HxrwPElxwZWf4FyJa6PJCt
dN7aqNkVghzxS1mcl3NvAZtqdpIFI5db0s9J+8W34lzZmyZyaW2+3jjlai2RSPS2h/slXRP0vGw9
zp0+FmVrjiF0C9hHiYiy0BkAE1CWtTogAiw3eM98Jb1zk1+atsGC7SkhKvQcI7nf4ZnURhA73yxt
kqUIwWN+ybzPiINv3Bu2DjH8G3j3KTtsjcCWplAxR62Ye94iM1XK1uTbfeMMcZlQ/5xVmqLx8UXh
OP3qy68JF/iH7NdGRidofFwhNoUgbA0L2KuSzJd2Av24oBQjYfr/dYjCHQJGUFSYSxOqkC9m0ilC
LKvgnhZGZeYZMvVxp9k0XGFvzHuCbxMss5Cikcb/ariwssN99f/JUwSzFox7arIc9u1gmxqEtomV
JP9cEyISgWMA4w9pkgC5zb1FdUcp1JrK2vHX43Q9+JNBZy7ltHTSxRyuC/JREtKNQZ/2tOiNs38D
mrx9wPDVUTJw36CV2uscIWBqpXytaXZftWucPHHnaL7XDWJEoQjpLV43b8Cqez2FG72LkuxQmFNy
ug3rgYhWs6q5cu+Ysc2WBFsodf7d5VIZEYK1G+lQBR+jbFQNDAGCCw6RP4yvmMonq2ydhctm5SGv
iwrJt60fcAA+VEMiarFacUuEwCQ5nIDgZ0ptzWz3gNLIe8GBiSNBuCxitCUkSq69spwRqVwHXQzH
l0wIo+q4cYVHDFR/kE7/DDC4q3Gm6TazO/I80tdXYytfqX6kK+aiThm3YCT8YeNtIDA9U1T3IR5f
VhtGtzzd2k+WcCNL931vlO/ioo9wG6ra1O04PR0Kv66xGUO7/aEIXxF1wCovOiTYP9rZ4VD9FKB6
QtxzU41CBDp27PVOY0aojEC2pzle6bDz9k6SS3d5BUSrG28G5Fr+Brr2PZoy77eiLQ8v+mZSz5tA
0nuN336NfHkrMrwhXmJ3bNEIy5RZDuZDHqtsDDx6ajQeKc0gOrprnbyYKxfAqWnlp2EVKcV78nuH
iJVzTVfizOWx+TyHBnsnM6gtB2Dk5yKVBIfOzHaGK6Y5Gz7enukDFU1/tCpmWr6PSKP96AKcheFq
XzHgnXlF+yubwP0XDdbc2HUzU80shdnrZ/C5FeQQi++swxUEFa17S/bzzVoosRcT78ir3bhkQKY+
yIMEHSWUM2Y217gtLylqFPj8ndNqlcsLVh+a3o5OmLP5rbxigXUJgC79KCMu/gTNZU9G2F6+u2Ai
KHc7Hrru1o9ZuFkbBkOzwxdG5LYz/BXObsx2OI97ByhJYF2r62c9FuuLpXa3+E+b0vPZgQXC8UfQ
gMMMHkvJNLgltqx2JZ618zxOugKhenlUKuSy/oi+aminf08d/7Tn5V5O9DAuCFYn1H0Ip3E+gzeo
0XyonevnC7SoWVEYrjyQgYQIcTV05Th7J20+I0WUL08NN23nJoNPXZ/Au4XLm4+ks3j/NrW/ga7P
H1t8zGWAU6F0AkdMZenD3awO+h6N+bsq9dK2PI46R8naZxkp5nqZtTtqxy/iMAdT1clt/v3YKqIo
V3afY9owioW8Erd1f3f2T0E+XLJO2OjDYY/TQgsTrmtams3iZet8UIe23e05po3oZBDfHWgHVh1/
bbmd8brHhyKlvjs6uWl0xEYWgjxT+Qpx8kAFw3mWBUk8u2p/kQdXsQEyd8yXoTVTyl2stSfiCqgZ
V30aVY2JVMyT0yawR2WTPMWXOn3njzWB+SobEdpjYn0uqUmDHguTaPXR+ndjIVFQ4BNahJ+mKB1w
Pk+8190+PzZEvpumjWe2uDPZVonKA8UkQ2movdHcvOd9v0gab863THZMxcLLITzzlgG7Rnem10KU
LlD5k5zQC7qaVo9DEdDslRG18lpN5yS67ZRO4ORRVwytU85W5z0b49adw15Zc3vr0zv75D90W9df
VwnKm9PplJ9m4zheExTbrD/DPjsxqm7g40btXeflJpNrshenrzJ1xys+jSJ1GXjQQneoYgdg4yWi
5R/VloUbegrLE987OL39EwHQIUbbdjDeLGvm0K41i2Z9ZnpDQKT2F+c84Xeoq8jTSu4Nwvnrw4Qq
BNA5ANu5Kz+Vnr3vJD6hmBhJYBXxdak4xJM1aG7zN+k+HzB9KsaCZ3rkIHgmxyeVA6iCAlgM9l63
I6mFyNlpBbRpwqHIPzRIV8KnH4o3Z222Aw/Cw7ONccCVujv5stRG1zl0YdiC9XWEgXVe9s6ZUt16
KUwAni1MvmUUkbKRuU90HaKHOBMOV5YxZzNJXC+beyhY7GNNYxI7vtk9xlu2PbaOe7JpRG5iURTP
KzyLixxElDtGVVZYtB2JiGNDQvGXicJUJjgpYRpYicqgYfP3Zf8sg8ep9e/HySLLvFxRDs/UZS/u
Y+2aq9ENx8yTAmC/20goc9op1/AbppaYRgR49gqsWW6cLbg0hfHndfvAYHDC0Tdb1DvGf3ipZI7m
rqsg2O/C0soK9fjLEOaSyL9otYe6ITHRaJpnKLvZY2oUXAZPXOMtdVEBjjPl/bcUJftAuAxpjCeo
wSFrnh+/hiEXlXECzBfuxvThkyzkRYn+fjl8uzjOLwyMTt/+FkZGRrHXrDrKaiLjwcjrgU7CWf+o
KQ1PmYMoSTyAePcKrJHvy5Ia9TUid1ZG3m41S2u8bILJiDov8qxGPviYK0IBWtVNsW4YsZutnNY5
MOMm2jCDyhhDJq2K71P+zQtROuN2Qk1JWjfeGY1FvTH2vikozQUPl1viuXkG/r2ifJfQh+w5KIr1
mJ+2VSoXDijXakhHs6oEVDloXLCUw6zS/1FcUt7hsIZKjKshZU6vbt9pFLDB4jL17qP3KSHvD3Fw
dhybM/sUf2tP7YaLHg9x0296n+2SpT5W+nOX/iKeM73oS3wUMx7nDKol+1RUN+MH//Oz4B7DxEQf
H8XwQ1GTI79UwgBXjVtb8ygxDPp3BUNZXP2tzYOP8fwqCk4MpOhdFtMgXH3iY0LwELZggiJF5k0U
S4NabAJiFRyqoyruiqPm7ytpM4QzRLK+vwla4MVR13pj94uKMfKs/Zb9maUugpUVMWZ4bR4QILG5
G+sulqdNho2Qy0eHKheest58L5ySHvAtHsIOjzR/9/bEfykCQoV+vlKXVvSF5uN7llgiR2/1NXW9
MN21FIj1rci+lNjiIaEsYBiFeEpVumu3uy8pua3MYsHG2zmx9SuAwIbMQ4lO62CDbHgPvsKVg9G7
8YJCc3ri8slouogWV/ooE/RPJZDfoPq6WClBxRO36Rm9N/SGE/NaNqtfwnwHzYxi5AI0bF/WTWep
NMbqqSD3nuaoSBP2faD821Kp50eUzuaL05CbDLnqteLfiH5COTc2Ib+f1ROoutazCxo9Q7DYmdgC
bPjjwzn5N6Sjs700Xm0h4SahTgAIy/+hO3/ywohCzjAtAS+xw8b1C8EzZ6lMajWJHyecAiZjrWP9
v3XL6M7bZdzlmo0qMI2cGJUUrmpeontpgyCY2SIGPvfJ0WiNu9pTi3YTYqKj+0fcoO1KG8W+814+
8eEyWRwupDnFDT7EfHzEgN9w4OtmAQ7j0lkRmfQmK6ZyCz4QwLsek5VRab9QWUFlDP3c2e91e6SW
T1aajUm4ZYRcaID+2Xw18tepQGT/12nP2bGPFQz7Sq6yWOyx9QcjsD/u8aIjJx8b6zKdaWZvu9G3
0owjJx7J0kt/TFLdNWeRP5I+ENf3hTBJzPCif1uANT8zhjqVoTnO5kKPE6gkt7vcKgUojaJMDMhT
12nXh6/O/Cd4yWURe1w9FYRCZIG6zxkGCx06Gzgmz0xVWZB9IRXfjH4yh1IfIQ6wIJzeGFOdVdIC
/VwaEzX7C2LW9lKv9gJZtXxIoKVvwJSuTPRmV2V0bawzxdFD49pR7Bv5E8HmNVIk7dVgnJnAhd17
VWF6w89s7mpzxLhRzfHNAY6qUibxkD/+qhN4lhebs4cIRFqOk5+6xEWPbGtXoIxtgd2sm1WZMRD0
GvwjE4rX7Nhfel9sHVNHk5jAMZ+xDDdq9yjp0oGT3k4W7xWmMHd9HmaV9Fgk3rMKwc4bhuCIvZV/
nDl/qqIwOYM2ccBzopgPejZSxjsZQIdC/JXPuptwa7ZSK3u+AB8hFFEB3EqC7WeSNdWfEdosBbu1
gLnvSQGk64CB83XrVWxac7LyleUuMt63qiwoyAjpK14dgnwF521y8N+qvPvrTGUliP1R5C0EImwG
2G80Cifol3qNxWWznrBLO3wKX0+2w/VV5qBkJoKzTUtyXJ+YUfx4k/pl+enI+EOFqutvRo15JCe4
ZxEUV2EuDTcFFNQy8dFEEFMnV22jdTx7ny6Y1Oqul7q291hqSu5Ju6JTkaGBHcCgFXGWxIQe8t22
+Q3xY48ofo/KnJatNxP3mvmentg2EtxWdDqCwIuxKrbQJPUPRhdPhrgnSeHtt8wpgmIvecbiqojb
eXEpBtJGPxowwSmbuw+NbvQNGHdi8y3CndDdDI9vORRyYsZklDimQ4N0jFyae7Mjv5k8ARVaI014
FUQhBUEAHM0XPcVqZ05PDGhCtF/+/D8RTemUOuHmHzQKG6Zo0DSoVvsnJTZJrsRnCFpwYTskvodZ
hlrGbXIzUIS5LnXM1VO6CuIPBTf2ERc4WqhHoWyH/DGtaleOHZmDawdutgXC5x774JVSq8juLwhx
Lr2c49JVpogV3bCzAHCpAan4VDGUxC8OOC2GpQZ39DqdLBnp4NJMBEtKsAdrunFGtZP4BGhzzFaI
Gu47Jv/zl1/MeiimmybPGhdHtlJXQUb98r9UH6Q+zzTabiMpqoVP07PyZKsQ4snAl1Jbnl1Pcl2Y
cRALSEwxdNiH9KHDLeg7sn6mbCihxaATTCJ+lOpK1O70ybyPyvx5C1vNUy4CcfA1XxSyUnBoy/dP
IyuE1PEjRr5YAslu+R2+asPcR92El1HrVWrNjbwNefvW4mvyOByhMHDyH5NwMcWbIXBSzS6nX/sx
JB3isy2UMZP9tkor/oxQC+Zo7AQ1v4XyfbCIHry9CK/uuK14PlGRhSzvz3wr1fmzXEm4LktSXod8
YFEjGlmIw2Kcm4iBHNIIQK4z6yL+/JRn50Pp1MaabUyCHxhMBltRP+JV2qG08V4WjQaoSrdwSdS9
l849qgSAGsi2gnAuuD//Q31N+PPDFvbNEfvWlFuVXMXQxLriOWqWHtPTxgu+KgwayfG6kqa6vH2g
gT3psnFyzbPU0jc8x56F1483Hi1hNTH8+0RS9FNqFRtOjBFKCzpXZ7FEbMYQrKfOVc0H/YVeNfO9
5cyhspAxPE6Bh0uZ0jQ/aMJyI4tPDXk4Ck4qgGngOaS8A+2m+i9u06/0ZYjx5iN6ta6D07l5l/vF
iJUAX1cTJlPZgIRoqIszyIhY9c90qoonDviTV3e8xqWlzyV2lgFaIAiRVaajaYUFBjSTxJ9ox1sQ
dlTILwoMtqx7rEoXG4jrrktLcYAsAbwnE1D3jYCPvLieRg4cjKUVMiSMq39KfaiJ96U9nu6JECUi
wJkWky8aXJxy0g3anm9Ug97BHpux5i6QnBPDpeunb3nRVDgR29QfvJKMJvTbUvoMEHjl7dSFXwbW
Mopmtjm4W6fvhSbHpuELG67F0fQnMdU79yJiIKR8dbv1J+rWN3slVzN6NKgUV199TweVdRHGgzZv
KTKFnQAuYupQJrGGM2FnS+QICqBQTnyCMm+CRpk+aPyq1HiLoqnYwSPhT9IHjTFckzdtbst3qnF/
izt43NB4FI9z85D5DPYmEx0sMq/FBtRF6wpwkcB46BazERyTW5taH5h1+11669Mald9L0t2IBaAl
rO4IV4txcIhMkgIrmlvTkGDKPGmdQ2XoOR5qDE5c5p3hLv1z3y55FhI0hq+ovw1nyaq/LrfdmaW4
4aZn8t1kh6+sTQ0BdEVMpeqi8bJ5wLgt7428EiMGWMbym6PIJIyjnkMTKMBZ9fbmvHPT9opWFZeH
U+6Gzerqaar9eRi/1efVY1vztFF9yvd/aW3roADKgtTxsIcLF2PvHER8jF7IAKC+GE3X4xFX+c3E
Dfa0RMfOWRBP5ARk62EHWlfaRcxfug9CXkg++j6BvnsrWud+WFctJ+Uq8FxniQBaOSM3r1IBJ04h
QRDHPF9L96A0ZJS/1q+5Qh88GzG5kBq2pTMY8j//0t3yCvmv+7eEAB5gMbFYnPKw7va4zccAFD8A
SZreOMboDz5fWV3xlmu+jmnA02FrTtmgjbzx1acWShDTKo5XPMwU5MAp9K81zbJuoEULsnKT+/FI
IdrU/CpRMx+CF3ZkeyD2p+h5HEyteBsuXW2i2kmv8C1rCKXZVbORT6P86pewasGUBd1VqkA64hLQ
lgPC4FLU2bEkFRndCzHxstIyBaubMa6zS/xjU5fH4UyIYAUB0RQ8mF30WH7JdcD5mrz6aX7LjOdq
VmK67g32bUDWgMc4n10kYH+/JOaNRhE4ElycEdM652yioo2pM0LAzh0bmYiZrj4Z7/vdXJDCHUkk
uAMdnFbi3GvYUHd9jQfeO5SVSMPivBLm7ij6qIMk1AanUHCP8WxntnNaWaJXk08eVmPENMol4Nkm
BuIKAOkmv0tMFAhoZ1aNXNKXIBq0wIWjLf/QQEcsC7Ua1m8edLzzlIFJ+FwI33vVFU+8zYNlLEnb
+BrVsq3XR7ING2mYovo9ryMIiEkzeEHN0BpL7iDClz6BBfzQsWoVeDjO0gcZehxXN5O4D0EbImE0
cug9GQiDKtY5H7DYp8Bu5oR2FMp7RyPJcX+8H4aH2UCkvFldf/tcQDIoVkP4N6SgWUS4XsTS0vnf
JmR3dAaytPh52/vhzWGCJ+KJbyojNlHYIWDIAE2Xif9rHhipZpDid225vz6rkkAwd4+37/iBQ8EC
vjlpsYwEidQYyJ7X3UT4UHARnNpOn97HhIZXXWkZ8P0l5l5hHod4cFwBtGD+3/QNEQjLtW1Q/RFo
95hyfVfzoqy7AoeIYmsNNCdFvuXIq7aQQ+lcTz53XpiNlKQhzAV9rYlkQDdmamo8xhTxBFQPoQct
AXz1kggAG2FksJFJodjh8Mx/Yr9VAEgLOChMxlHCil4UpRrvQMWDtW01XlutqWep+QhHH6/7enCf
01yzAfQyQbeAAHDNd3tB/X9cOo46oI472Y/sKnJfTb4aDmbeXHtl5m1dByuVCFOX4pGMqJxpRdvH
lzNUrZKBxbnpqNS3P/nDrIC2iamIVAVc7tP4cSSfinTVIhfVJgAjw1f0+tEEvnOQJNkBG50jLYFH
C2nN7sZIOJRH66DJO6qNolK/aHVMjg2Zn4glCI5wGm47y8SljZ7RbZAN6ZFz4PjUwdrdhyavFCfA
zVBO3ZHNLBIBMRE64o+NhCEAfgMCoVRhapti3ZK2q2AORmMxuewSisnrmU499MNLq1VBIHrN2Ciq
VhcXXDC7eQzP93UTt0FESdQHrDgsib8M4GEB7rboKu7vVAF0hObuGgMCUALXr0W/w7ct8Fsxuk+o
jsNEuAM7HLZzMYBS6NpIs+ncKflnkapZ/U4Nb+7VFkfvSruu0hIRgib9q0whNMIXn1Ay7BRjYwTe
RYloQGKwAA6ljOB4JXzyJMgZynGGZ81BoLaDO9k+mr710unE0x+AbIaUUsQ67mvEJyerr2/9m0/S
B/VsPSW+7PKKaTLQSc/E/o2wThF10N1UfONTEeLRj0A21z+C3WVljoJR2F7HhDvIsnAYa7WBp5ir
YGfO9gh5CwqGlsG/NmkotmsKXPbBxvr7JaVQSP+Eht9sQBxg8/q2ZvDjM70PK2wZdoNkUTJP5pLc
JY+ygddNbBffYFQUuaYsco/olFNpPtDxYjB1DOu1SeIo0b1lChHManYzQ0QNC3A+lKanpQOqCGqQ
9CGpkQDE/9RrMsEwYXMBBc37cjQGl6R4o+46N1bdIYtNXGiME+w1ueDwrQSs16noYXmKaohhpRdW
7wdartlbYBAcsyHUShxIyyBUZ1W1j4s9gJmu4ludowJl5JgffcDFoLWmJEM+pjHdFAvpof8fox/u
KeNcSANAjP8uX336kLv8jf9e2d4myZ2StpKrKh2L+pyEX7yaPa+XaDnUpJwtpw/g1kZJW2/ox2/3
DgJsMErWDdQcIj91VQuDGjufLCyt579E5+gVfClITcVJGiB9xh3jNZCHuYiyKyFvDxiWRxbEQ2wb
/B8PC7PnAEzrSkjtNh4Z+BPdf2PGhRxbTcWWNmzDVym0iUhDg6Ttu/ObMjlHLhEhPlbe0FgMEwEo
efsb2zns/xy8uAS96N5AN6+B+I/7R0TCRhdTsDgAJVfpFu6qx9PjWnAOk8nX4m7P7Vo7LirExCWZ
lOEsRizIoqVP/LYwoWNlR6sl9uzUGv5n9qS4xs7XLEWESy6PFFAteVM2awezFgsfRV6+eqYAPL4p
Ve/8v4QHs/c/zBJvyTRMOD4T2ZqqYmQqmX180AdkUqjCp5C5cZNCu7U0VM6QcXFGJxog7onBpzCl
ODqn2CCjgThBwWdZuFUiKjOaUnw2NDKJOpWsQSOROJnndJfbR88pIHAL0G9+pd4neNye62iO01xq
Rxh/G8EW3cpudIiPNTP3HyKyFOuxVW+PxRUQsg07LX6Ja4fJWW1MqSTgausRgGyFDvGmwcAHSJOq
hQRZFS58M0EMDyHrnFo1bTqhDtTeVepMyPSlMWgDpnYsvOc7etDJbMS5wrFlOMkzoBVYHZhZ0z/o
e7++pOYlXbrDAj+72R9ei9ubk/Qh5LRiiRUeOFPCqyJiT9CkcJGsXOkWby3E0ow/P1zjjtAwL7TR
UsmFi+ynN3iPv/CClRwfo1gVkqkxzukNq/l+qUdZ/9YrfgZS2vnWSqxCJOI9AdoKu+uKVyA84CPc
7iPtpvuta1xBTGC1y3uN3SWquY9mr1lx0+yPkvmiICm/SfOFN2FpnBuBsMAKWgF16i/ZqwcpW7Yc
mKuGkmvP5hzBl0Pm8YgdwcRMzx0p8RvtyggMlY9fahTYlzRHrUwifL0nPWEbr2liSFX6mXB5dg6E
/UKpD2RPJY1Sh8OSnNdIxNNX0XdwsXBV1sYCurBGNL00momONV73XNjBqBj5EZjNhLg9ojoWH8ot
0sy1mHFD3DH0f3PEUiMv4eb4+QGBlnMLYRGp/U+byVOCUFyXWbq3NFH+KJsgE1zsbfoPmRpNUP9X
w/uIi/0tn6i8oOgkELRz9cSxX3kK2I1Z6kP4wsdwE/RHCJn1y7iI8FZ7XEVvZlPVN2+18qGAaANY
DXo2NmB+yDy5xJok6vTtbyAm2aCs044lbk+9OfnU9Y6471pKTXSSWXEkFRDeoPpWOcjIEOJGUz5i
W34ZvNT6ExtKyev6zmrVZR/6mHIi+DJXvaBjUmsttA5xfdSRSeQ5wOREmr9KavxcK8dsKYQIMdxz
csLoCtwTgBXRbM4dMrvSMjdDQr+C+oNc8L3uVVOI3/N4+bgD+io3XJUtNmGbssHLPSeQbT4bRLfC
9+fWdOnfIQyY5baBVR10WeCEW7gR1/mzYjOy9CE1AQuKtPx0VqBvIQvCF4VO4dsGUXthX0IQg9e1
DjJ/Qv1PkggUI8C8GGmvZrKPGaz3u4yminD8iSi+fcyCUVDx37qAOMu8EsFRF5DAjAE8TdXpzNyq
kgyuytz/g/gE8TgAZTs4INEdOl38buNli/KiTOJg7iXmm+aklrMVvSIh63+d7p1oQcB1i7K4LvOy
sRI/dW2teJmbw8AjGb7lS47KEdjLNuYmDwXYp1kFaCIgY3FZf9SUhfYEBY9JyxZE2mMHKv9/Q8qU
nON1wMOQDt+67eIQR2gATrmsqOIufTg6b0h0P+xzapR+b+FUJEDU7XovLUKNz8sxmI1yaKoet8ZP
rzu3KwF6By7lvUG+Jk7jTwawcdSObhKgUePX3KHJSoDV7CZnyaQAiHF4+chzs/KKs1UE0s8ggr9V
hw7pUoDAE3zhqJl7MKHyTdI8E4GL735OkwLJzYgnYb/s7WVXhn7ItUSbv/Z1qyBCjytYFqUlHtr0
3m8bK0zcIhC3o1U3nxmZywQ2RUn/V8MhQYM/d4ZX4vtC+atCKX23sYLLh9uWfdUKGR0dOEN2hEW2
Y6WRnk7lPmS0P2tASOxwW0N28JjebcCTYC/2vdAwgJRhbcrQA3VWMm2MAJFU03RirpbYZdgV/M7N
HqOGQ1P/Ad6qTWbe/4E1JoU2J2yaOTPG51romXjS+41rg2pczhSyxyILZO7MIm1uQMrmTUfVOr8B
RIiK8WzSCQYV2s02cgB5xOw1MpdwDSleUZ8IGys0j77uIGHp5ov3nBbXqdAs6RcdokBr2x7O2FqT
X4DpqFwYimL4XQjCyPaSCqOM4u6rkxXM42WIUPzrItv5qVgbhh+0m6UYaT180iX3mrt9L8/cXmoy
WZ9aXS/xgjK4czkpb5jTr7A0h3F9mxTiGNYxjVfD1ZOsKXAL4WtPVsI3ZZZYEqxaOsbN1W5R1M6c
aSAIApTCszUjsIePz1pMI4nO/oQBxrFCBfPVADzbRfN9tk/61zQwWb3f3Etbx81l9zmhZLrRcnVZ
YYz1sH79p5BArldqMKIX8rmPYX04VUsuJMQvPd4n8p/KKE9gb7KwotWlliznNyMjs6dcy4hoV2Uq
lhcEaDBkmFCplebPMCCmfnQV6MYEcgIg/z71+OKAcc3Ta3EODD2/tbClabuZPl1uX4jwnbCbYXVL
q04m3fLabmIIxKQvIoXL3HZAnAxBWs3hHj8ze7kVBBJuQCqKhTySKsdcTTmgKyr46wef2w+zlPxW
yDOy3Ir9mECEuqUUxDk8+R9xA1p6eJLHp/TyNrt42ZZ8wST3LuVvG35VBKdYwsBu7T5RYuVe3LZz
9ujiX/EW/XRa/eDaWhZZ1FjElywxSd9EdfantCodTFDFFXIBHqYMq2PEyPEOJ67++bha56s61u03
+2QukrEkycheSa+c7Xr2Od7OBXjrMzxyhACyBrQMxaaC7w2Nd8DUNhTHDN1elu9QK6tVP8/j5gef
UTuHPUDycAq5coqRnkYTdBOIJsOi5MCf4ltTBvVfYXSYeQ73yHJJEU8ozyYLpGi4RPnh4ehbQxV0
jZTZbmAe64u71wWw8D/rLz6xXyAA2RyNFUs7YHjgZG2ulyrSZzVe/sK2DEk+3lB/bpmezZ4W1rkL
fBJvmA0fV8ThrT6/h3P4cFbvy9Y2HalKwAnINdemMZR7NuGN5H7bVfHyABnJDJxhEWluDAtab2/p
sOWT154BBlnqaxImqvPlfLmTFLMAYFvcQB+bsH9yAOxy03nPtclTTd3UMxofOnmWZ90yzPz7BSUn
Siy+9n/pNH+DUDzvwQULTVwPvUbYB5rj3ThCMmQYfwwcYZ8mTVLgv1ybeyi/JqdFSJws58ln7vPU
3y5G/qtBFj27R4vhSMIBo3iJcGS1uThOfUGc+7sGPzzuM4KpU3yq2Ot+7WZA0KwVqHgHCx+X3/vd
uZ/RiSHSp/Qufabs2GgvuIt4vx8hG/almj8K6BUNsuV2I6eCFSVozScedk90z2+4mjqdUkGmEZmP
zdGY/cHuzPV68J/mLgx8qEBOvTwBVrE40kQobfty2c47odgSfCHEAE9/h6zETcHb9za/6x0FBAFH
tbPMvqqMfehCb5ZeV0sx8qV+rM+hYUyuo656lTD4cAY+m5+oY/VrZYVCMQP7ZuGTrUI4rC/XDXBm
CvMusjodAqrsDPanV7C0VJv8Qasxaf74Hcaf+6lmjTIJtQaWDilYImQz+/QAvqoAkZc2tdfTty0U
+646xodlQqzgvyn7tkBVNKSCS0UFOHvHDwkMYX8nVKCJoe4UT9Nd53dum1EfmdSBiP+V1CVZS4Ox
TIumM+sxefD9b5ONC5P4NU9TwDPurumAO9M1j+FS3RkDd7zaTPsfTklUzAtA8dp3DZVKEbU8d+eG
AX+slnFYirQ02a6l4aGDUuiE7Q/gjebtl8W+SAfO7hdOkCU3gZthMx4iTINwXSMq3VFxu3MfUbWm
nbDoxWCNfWhxaTNocCLyhF60vX0o562i+nwUfqtSCqJ/JqbYIIjnN4FgalT2+UyhETW/D3RMnH4T
ayQl/AQLINohaJOc/6uzjtH0kz6h+Y+7JaugmKClZoga+aRfunr1qxbmBJIHTrWNv/NqmIndMeuq
W4IQCrOkroWSYI2Xvznz0+Kyo/9PC/t8Yz4ryk/cklqSumxMThvOMLmwcH7rrkbIGxEOVmb6T1Yd
/NP12+7LTwW6Yhh9D47+sL80JHX9iF56LbNu8gisZtmu6hpRewfC8ORqBkvweGYN+mSynbPMHSEE
BaLkT1tFpfeEjv5CCcAlIH/CpdoTPlyUv3wQKRD80AhBY1eWxTP+46ll7ocm14y8gc2DjeCHVqAi
rl5AYPlpM8MnvbbwKfXWKXE4vcni1fnehbWTDh1jMdpAulmo4COfvZDr62nkmAbvUxd5RKBt83lL
Qse1qGO1LMYjXLoAKskOVTZcEYyE8wCQlPNdsT89voXZ5CyngwrXsZBGA4F0hy1uKGbiVvOul23O
bXhVR2TSwfIFtQrZHkc3Z2kqtB61fgvvFr73EZ+Osuq8PaGBGahGT7aPvw643AH+UJxFUqwLLRmx
xbnXM6Sic6TRaQ1lNVAEDod15lFzB09kNSD4iU0SpOdV8dScHT/lrz2iZ8J81LeBDK4y8XqdgRjP
VoeOr8KhXztuobjifOGT3JX61WYJKLebgIkCq+I3VFq4kp76cMcO9u5u4sOfd5NwVG9Blv1oT4qU
WzoNt/1T7K/A/HsYCAEGW27O9/MQemwIel7BpyL8O7ODcLqpdV1D+rlLuxx4uX2v5KN20jLwquqF
aAMWlER1/IWZZZdY7tWccFDqX4te2GeTlUcqaHkJldOwxIRhYLa5k3oDsu6IVkHrs6OPCGTnlwFP
LuaNb5I3j9EaWtyeBR7BzjnU+jZQB0kWTnwIuW6KjAM1naaKQRhDM5V7x+jIWnE4bTZsazvwCq5v
0C097sC5NaGTPLhlr6z+ONfZIdYIh/zI+8tAow6nIpkXOE2kIdpK8tpTnox8BK5Rn4eriCWirbNd
GKIw4rYAiFEy5pB2R4kIl1Da1Pd/2yLVIzXkDE5tN9w9NP1Exo1oi1dXb++dYryTuQV/ukf2MhHC
IaV/ebfuRjCqJaAyY/fzgT0yh3JWz/2SVanD3HY6RsjOmk1u/3NkKKxaoL2uAA+aCPtL8miLeqlq
qVsGd2xmI3ZIXhjgYAcMbJePRlk3ui45OJo4JT6luVkyE94Am5Su17s188gDWor/Ax/Kra6virx6
v55jUODqxO3kmVDfqhlQAF/xmxtGH63DqBTIBTnBZrIrwQKKaOameNd5Yem4giZmEYsu6yB/NRtY
RoYFILPJK5hxeggEZTka53KOoobQedGWAU78+ppLhDzXoSqX7kKeIsF94tKLOvyhXcH22fyRpfnA
Vk88/iSCLGN2efFD6cmpO0z2ogjz+LEKqmt4Mc/IT5aR/H8d4WbErBLEJgd+5votmbeOe+43rcU5
ooxlE78rRAvRv2R6a6EY473g81sxEON8Nkc9n+OknhGW80zTt2pVt2jBDoJwgqk46UmbmFW66xWt
S6C+rtx85FDFOs9qZmL9SPYbDycfRnDIKtZrO6opgYo0IO3ZeBNRAkhslX1u0YV1C8R79EGC8EQA
4bEu7PiRTw/O9FBiZuosXrppDrlgEuYyDQZnJjGrgcjicQF3VBkkL7a2gj8/xP1/IKOUPcLH/hFr
iAdIQAJAlgFK9SGtzn7u45beuczJwvMZHscSSIyVp1ktS7+1WITYxVn+4tPFbRuYgHBfY7EgxXSo
JFPiUl0l+NbcrroFbigR3eoS+5KwuuzwFjPnm7+AsvN/JwgboND0diQtKLzKR+mBvnCohlROuF7p
wVI6rGJ4aW/B89W0wWtz898RBvDYYVYGXsNw8USHocnlx1XoNLwqt2xMukXk5hTtkK2Gk20ai09J
WNC5rbnw4i52gQkHRNkZUBRSqjyLxNl08n/6hD/t4q27Ff+vx4fjELbc5pA6weu1VVBDyACB4OMh
KLpmZnsWKXqViSU94CB9lLRvqVT2XQWOYkIhKyE/gWdiJ+5ns9qI1KTEy59/vORK1e0N6XDJFuli
WhGud7JclktXAomx2A/9qOPBzILFcboudbBfkpgJfctu6tJYhrEtNu69YNDOPloEPAdm0Q2cau4m
iS7YeEurITd1c7Vd5qGVf5WEJurAlT+/W9pWjX3x+c8nmQC9YZCYQzRxqfxI1bifnpLQKdTJzl4T
wc67yP5yx6zK+PATbda5LkqX47DmfI285IptlcxtdwRIigXsZdLpOKFiAJATdVM6EADK7I0U8R/0
r1qce+Cx9BqrVaMzeCeusBKobTqvTwa1FT52FpWab/YDlmmRcfbIk8e87m1ZLQAUC/4oIPGT6kbO
BNhb4XYa93rlVpBwGO8cS1UWpNFUGqZz8sfg293lE5oSY+1d1nHspRt3XfaLQLIlg1G9UZXBA9Om
azbsGwy3/o7Ma26r2GVcYsTWaRUCW0gLC9yqvNhuUsGktpej7wJurlrop74eNw8RfVdNnBm4gRgS
+Ha0D00ipbKFMXi9fmvXz7dpTpt7BjuEEIT2B0t3peu6qB6/w1sthSz2Qit16WgzvYphWo2r1Con
CFYSMQqnJ27gMvyBMBVkqyT3lbX7MT0MaZjM9a/zBqAIR/Nyt4IQRaLi3dpGuxNEcVNRAMNC6+5o
oRT83qfU7G7lTm9tgkjlklbqddxLVzvXt9vSPhQSMmo/e6F2GMcp7V4ylD903uGeVFTN9EeGBM2P
HOx+24Sc7Q3thy7Ubj6bfejDA88unH0hemfsPA7ZbhL4qtQSAZslGS8ldv/9qWnm07iksea0hFF8
RSCmwfAMbhZX+Zv0imppEwKEOyxvmPvSxbikoCyebITTLcrwehW/a2q+UFBKOvPk3Z1IP2cjTip4
n88EOpgBn9n3/TzwYYsW8+Ala23cUjQddz8RjEjC1fQAlqVnhEVRnMTqal3zb35tgUAueQ4p+kSt
tg/DRTZnS+NtVo90UXh7feOArXDJ5iN1n0q83x580BIxKQsJvrZUpluvsToIiB1m4VgAmgkwA4e7
cSDSOKPQdjFAjNzJfXZSlrBP41ikJ+o4HNaykZqdp2AMsr8hwPsSB8BC0eu6RY3fdUZ1aJVAXPBU
6kMFWMC0ogKNMVUMc+7HQgau5IAOCUepQrH6inzwyAd8ZE1YJYw/Q5bkVyT/JhiNoR6Qyhjc0Ryy
cj1gMCAVfUY7BBIwL/QHWiQlJTQNtHIqYsfr/jPky5rAbul6Yg6hCizuFJ7fLWWcUVzlaKUR81JD
dILNNsbsQaGgcNtF1qSZ1ATJN7SNIq7GYPtOnbLTgPdBmOP/79nlpPdYv2jPHf1A98toMbwP0cPc
K0EJ38n/jZTcxzPGhJ40BhLXGG/p3ynfhRJyqRvv37Al8IR9jNLRIzcF+CdbLOIK3M/IVU7cikvT
/dHN+kCIeevsjRBTitq1DC/MCUREoQTIrb6mwtkTZU5SGCwqiLFWze66UryzCERITsV5XLQIpVpR
Oo1Uyz0qp/YT9lJpbgKpW1bL0vuqj2BreT13Jyskb5xn9gPDHr57e9wiewXsg0LMoIDlNrsnn0mt
KKnvBEwdhwbL0+bVY9acxXapbRTBVhNZ8G/9gxAEHBS8cLOkbQemOqFbYKJn2+VO/pmcWUFmTS6q
IKZJU605mNoaRuxFdzpEpn7yFpuCUb7nlxXATTWTSPArAFeJU3dFid6MLwtQt9eaRC9h54A42YlG
Vz+1Y4kzhfdDhyV9KYjGC9BbNGviIvMx/F0nR/oRpc2pBJ9CcbHraP81duGyonoObXlJF7hJbGEb
QO3L18NYByvVkaCtxn3GOAMLGaOl/TYaHE8od7t5s1AmQJJr/OpBv69RfQEckiaSgH2GGnLjg6P+
Uq+FT/SpN/pLkHHa7a7IXyGoxeRrpcJGQY+QL1PTYEEVk4FnfDKFMxLWNPzlCCspXQc426U+f0uo
eYskr2RZarC2vsv0KHNaAL7fX212F5n4bkyThA3xKkY2Yq5oFNatGgtYqlSAPvNjOW3/GSlJDRF3
Qy1FYNyduzDlxPPdwvf8AYB3oBZraaHVN4oIaBBQh5PU/vw+uGqaee7RtOCWzO9T8YWAGTpwjn7o
pdjX7JR5dvUe1hFzNYHZ2HayGFYuZ06JL4jXebJEe1MpEgCisTkpJnpmvGXruDL3P71PPz7bjKEZ
bbQA1V7TXJI2jLaTtnsvJb4ybvyY06erI+2tjW5D81270v1Xn/qjbPlTOyywuAjUAzV6lYy7d82A
M+6U+ZTUeUhmNmd0y7+SPBKDi3gxX/mfRbQUXfl/a9SueWqUhSprtuOB9HZmfYZiBsEvzM+WkeS2
tQ92spioUzAvP3rNWF66mTLb75V43JfF4EJDVrKdIgqtePVwO2b3G1bbkZqbHO/zhLRWuRQUUYVZ
7r4qDLG4vKxuX8yLhilY+oCHIzVp1kuxR7m1aJ3ZrWA1tNo6V8NflCssG25+fZgxRZ0RH/ybbca6
iHn2oGufzdH5kigcjEzQZ1yUugMgLBB3KQbtAikkU8UmLril4FP+8SVBWmWZ89Sjt69ErQvMsyVP
SuLhX8XpdG3uwWKoBD82Fx/fINS/2ksRbRj0W6/0Eh6Ri/YThjN63RUsLUaioqvf4MD+YINFWUEv
w/Q1i9nsVUMJMa38BRPK33zF3hoU+Z1K5izSEj9kkkMXMRQGOr/BuJG+Z8T9+xToeUhgVYWXxiNS
J3t1nsbNkkvRKXzczkYn+QEcT0C0PIKFCcUuizY9EJXTx2q2F97XR53aXq0zS5+e1BGaWwTjQnLp
t99K/PrRZOwSrQHFjbPHUH2ZTHyMzjFU4MmsG7tBJjAo8BpHjnNysBl/osFJzTGExfBL0Mxfilm2
5l7Hi8s1wX0FCsvL4VFfCn4bdQbFhwHcm9bceGhXaIqwvhNCLWfOJ1yiJDTBsD/az05ymuXkhEu4
Oc6gCakxNK7LtCCvnnOxCNEcubvh4tMxW4cnZsfzvEUQHbgCs9CCrNnCaC450HiVu+gCkSAYdK7F
94bCtZKTAew6jXSU5Vj/hHI0Nx/lVd2ZIPw3dWkZnco5tz1odTO5n6THoGFzGn9evw2f0cMPl6jo
qehvRI0QPEsVn7zBBjlpOWX+Rp8q/nrvLsKO/E3epT3icztK6N3oB9XWMnw3JP4ATfhsmtUSnHtd
zw5/MrKgYUz1aM+tQb/H/Wgb3J0RqH9lBvvtfAm2XrwkHZvgdxHCIkILI7BFJx5HZxHGIogCuNdd
M67TfQPYK+Q9QneDsD+3CQKY5Qn8YRiAYGaTFKnVM32ouP+Sz7n9tY+BLcncxabnfpWDVgdZ34wn
bxpQOjU040EWizqR+0knmtyE+Ng38v/xjVdkaSt52beTkZSu0snu1+QxsOON8pjcRPaniJy6/jq7
V1PpxQ/RZAQzMgWwzD1We6/PGlBLWoXZ2PbUC5sx8fj4XhZzppUBG4zDSYMGJDDpMaPmgTWUO6rO
LFgyD0ywjB/E6UeXLOLZF4hVRIyCDefcgmgU3/iWE4oW8RC0NUMdcT0lasW9JfryOtW3PKnYPk8A
ZGoU8b8s++gN3U5zcj53d8gO1n3L5smoBASgmwRhP/XYrDKtbjquOLX8uqaGJnh1S7J4vTuDQMO3
j6TjcF2oSBWWsGXrsUiR4E6NYP+cdXqRBlGT4JRP4TreGZpt+FFl29q9Dz0+D1mFTsJoK9h1Vijg
X/wx8R+1oXHA8dqFhPXrZHdBorMoDv7bSHMzDpk3sqayorq2lNnvj+qJzLvEEcPHYgnF6ySKwxgP
DV296HR5mY9QyP7TWEVh1IwcCxN0WOKR/HfC7OqPIpjfxmVbM6eMrPq5wWiTFhtE62VYHfNDBUYB
byn3lZy2Rxk+tELwZyf8Ra9d3JTB5EShOfAZf5nGC44oG+yixyp6WSQscGXDLF513QGEV80ZFLT8
JX/hLHxZWv8f2Qqq8O+pAb1KpDYYEDWzjyZdTJ1xJ50tKkThroXls5wg5OMtX2O2hQb4Xj2h5L3O
9booho4blsv2EclpzOgcBS9zR7MJ2yYuCPhI8JevNdJpjrJD0QJOKroteAhWS2pCcGrOvfasHiV4
LNAdzGHogiwLVck/hh4IjPl9qTJyysuOewf6DlwZh+tB26bCU+U5aMUZkFoHO6FRnMzA4AuBMlWp
wj0WFFgOP5cMia69J1zGjZYNRxK4WdYq0cmZQaOTF2QHy0zTway+csWCBZrk8AXd8buyFB+pkek7
97NwkaX/JuENlOAyAgwZUBxwwytg33z2FF3hFdKrJYRWJMDA90GKucrfewpkC84xMySl6PQbbHoa
1i5KpRa0LMrOAzh/ttj00nS3af4O5JdEdbQD/97x/3Z+OTtYmGNwxztZ+xHr7NcrWkyo14TEUeDP
ic3T6XVuP088A/kl8lzFonXGp/6sNkrr0OGSbPr8D6McmjkvZSQsaL2eASmJableGAfn8L1p8nsl
/rhIXAhtbjz7kyri8KlFOU7t15lJAAx3qxF3oeekYhlzmYyQg0MBRAhFE8FrFfMq6JqMzierYKiI
k3DZnuST70oS1FFklJQYyTZ5ibnIkKc0jorpQoPkGyytjKkE9XkXzLYeFcuigNx/NVbW5dmVxns0
BZo630PWxbkMQTewFv5kT5xRfDyDovP0ziEQTAEZrXrcapYW+/txOGYoBlHuwxaIsXYn1jCX7nLt
GOgd+c1VR+zBJVQRvlQls4BVRaqud63Egmx/mWRkAu3HmOWyRzGK3CnH+18UD/ua0afOVYBFFf1s
/BkPzUGb0doU7uwuZdLofPnR+SZHWhCmWFNcBMDXoX9ZQp3Yx0YordnaiSiyPpSHW02AI5/F8luz
czPKW80OlQKhYWlrT9ThXNo2udt4+oy/aOXD67ax7+mxmkpESv/oIoYhbZsFHq6bCk780Dr4l2RQ
+PwFX7R5/smrNNt2LSJfDboo7mTk1lGpdSdAM8rCn2rK76LFzvda+ICbPeMsU6HRpUJsKnKil1sW
AbkIgmqmDUig4jgje9uadaABJaeRpiH1CQo4wXep1bGNjbJE73FbJ5VnbLxfA1r2CrQat4Rg6Vik
oyhmd5PDdFBUdVkCCia85l0mPigdWmsM2fe6K3dwUG1XSoK9N4OWjyrOOuUcw+mxK34VOFGn7WMz
cJZrtkWC/DP/LNRYeKBTzpSBPEAxH0BrH9lt8v6u7HBQCRl46dFgo+OmBitt502FKpMsbsg7tTiK
nCtzN9B6tcMXYQqCpKimBq+JF30upS9djrSLFoD3iAdHZR3ltjooD8lZGOoSLn2/ji4NtvOy3jE6
mxzVxRw9G8DCJNKY0MjSDdVUxOBksfYfz/NNww+w1PEUPqcqa2fCvO1EFurVICaqVe40MyM5NLvL
ob41VC1Y8LE5kkLJ+fxjHKPdWYeIp8dK+8sWxt1p25woSFfOSb9fbC/dwnaLDeOQPl42X6iu1OZX
SOncHGdE0LPPCZnBou6ftrLcwSTbfa2dZZU5PkNVeKUt6uzts8jzRCvRuFfnpG1zqreR4pPv6t81
WM2XD8RXYG4NcjB93kke8y/XqUnfio6qT+LsKpHCxaDuLuMFpwPhog81QdNKBwMPy3wOruzcxiH5
IxJONlQi+ehl4Jyv4WqroU+VAQNe72cyeNhZOIWUYs4tOvzitylGr9CHeD6RfaeJe4PBfQcKG5Hb
xCu812AZtNowiZR73C0yWJ5K627wi6EbZ3mEiW9CTmQbhvn0T6xsX4Lzqw6whn2H9Nf6Eml9pXVX
LfHuiCv+b0JISSHWBa0IGFdIYYgkHV/4ojmdfmkNxgwJU0A9dM89Vdwyn+muPYBkTQ53DbwpBL7u
WMzoZqWmd2R4B0InF9g61jNwFzxNadLDC1LeRK9WjnkVygD3QZzo8WNB5VpKfxxmLKLd2VDXpQdg
1M6l9/HIlxsPXXV2jji24O1zsY8X4uw9Yp3c9GEKp4hG29ViS/Q1i+aSw8GS0XlSl/VYXUxi4ejO
DCof5uWRMWBOhT09i9Mh8QRdLoniI3fjx7MpeLtzbZAQ3au0USH14qJKqfPGWbOxKgT7NfuDQoI2
Eu+5N3pVXTadd2aLUkEIgym+S3u7fYTQwIXwFS8e6v7q+tykrAQE9BcufK0oSIbixoNX+NU3WSI/
miTkX26Oflmmy/XbA0hcz+t3JJMnCjoCEd4JAJWgbQUPP0sXn+hGkiTDMp/n/tbb8DSe8VAW8Nml
frY9i5/gX1VM4NG2nxnzcrdQoZB7H+lYnZYoSMgFXP++6Bu9LIvYLknPbQDlWLYa2db0zvBGsrst
+oVB9UpCGYMA/j9GP6CeJFAQv5+e1ZP0ARqtYmp8kIFGdJDFN5vBEd8ttOE/I85ZFopHxmBpHeZi
DGFmbclOb/EZppwasi5b/Q7QK48TrVsCwxLiLxllBwSefqnI0+3sXN4TVZZf6Eose40HdaiUiEjW
gx3IscZIK1QXex4WzCSoXlz/WtTvYpDFla615tyltZnRyRndhYF7UXAVx6DsSJGh1oUC1XS+pc1Z
VuXGjhalQd4Jq/q7u47KHPXcMnTPjEEwhPCM+ZiEbqedUf0nz4/NudCkpQMQZ3yNuVnQDykLnyR/
TCy8xKh2FQ2b+TXaunrx9q42J0ZLr0QEZsZWNXj+TroHM4djzAiaMOHj31lUWydgwd3siJO09cek
vxafzZDJ/d9h2hjflp9rPSP5y+x5nAJAhPzomWoIsog9EZq0Tj4yjBkcAtYT2WUV3O87bnMwdjoT
PUovZOg49d3n9OazDWMgoLq/nV0zlDdXuvrwFwg8c8RAkd2aXBVW0fkZsKrsO/Q0b32IwDcmsE9C
1w0AM/CeBmJWPsSJqFrSXPyX8VA7TMbxj/JW+8GqNQlaHuMjI28ucryvKdD5+CEy3jEcbRAp+/xe
PCJ2JwHYzP4/UnaBOyGHACK0hvkOFD2d0nrGejQJSlC9rO2syDlgZYProhvk0DJCFjkzlK3gu6Az
kJQ9Am8q1WldpHu1BcPErdJVwdF9dEwmmbkhg6Vpq37gwqDXAkCZtq5a/zAqKFjw8RvZstuilIQZ
4B3XuMlezeIahW/VhQDXVkn9JssB++ykMNbqpAbtWnHMyQ6PXwJ6nOEuRM3KMGuWAnS8STSLGOQk
UzidQPSGSXJ2c6nNumBJP1QwXaof61g0JQwiNcHQC8S6QA7sfReyV89xop7tyUmDM7ONVS2baGhM
sOzhPT8qWPvxZltzVeFlU8jbyjLj+rnqfFQCNNZ1SuLem5YPypjS+KKTcA/tvTLtWA/qmaDa5kD4
wNNSqx64oJpmLeN1M6jvm3uMsLDEQkln/VGwy2eLqNfmfC6j2OFtNplReDfiXo/xSEMwFh6bNtFV
uQvlWBZg28p5jz8DZtBoB5z6CWkZjy+7nWImLbfUJ96hMC4F4sUUnPDcohQuPMOrSRwS9IYI3Xwz
hY+6E/XHrbwDsy9qTygKYUCWpkyKUcR4p0pEUGpgIWSFm+7Lk8h+O3Bvr6nvNkkuuAGONs2PNN4q
eyXXlw9Cb5IkZL4+pTYDSsuJGy0NzbxwlUY52EDy5buMrDQ0QtW0pJeWeVlPtzW/Dk4TUIaOxBAV
lS4I6r8nesphjNukrTow1B9vZD85pXIEA4t7uAlEvMBJh/hrDalynzKbstAlgEHA80mSMk2p9dkY
KXC48OAYEzgbU/v2AgGH6O2+7KpTFKgPIl+yM5eQUt380J+17Y5Slj0nm+VMtdFVx4tOwP6Q51dX
4vYqye7Yezwmb8Q8ZoyRgTz9Bu6j0vaUWIW8G3E9RZ6Nxe8M887myRAJ5PmNvfv0J4NMvejwexzD
+0qNcx2+LRtC+DCv5nfSwWCLneur4pAcEjpBeSLdx9IRsStCLKHCEnFM4cDDbm91VRyrkOKEeqrp
NLo75uKUBmXhUrQ2UTiaAquHvXW3Q8L7q6DODcumue66NJ8H4QB+WnRQkr4y/JBbCpK/KkBbpaBB
NBKz7m3/AHBhq5xeUC+VQ6D0dw5TjhFpijX5mFSsxBkEeF/CBnDuhwxW+Hihy12eoQ+w1q4vxpxp
bIPGltEWfX4ckkZo4IadIjHFGGBQTlo1VVHQMKsNMPD/VAwyWCd9OsPZWFU/XN0wj826CnzR19oR
O7ZsxMXF52DtxRCGI/xcurt7OFFBrG5Hjlo6PrT8LO1ja7cF+FqPSQcdmoZUObpD+KUIQoglzjfu
XRN+TRxHQgVSYpDGvdQRMBRJnfJ1MkVRzvuWP/7++FZ6CPsK+u4KqL6doxRbs5i/X9O4a59fO0zn
1sJ3CMdIyoAccYOmiKzBRmVf5wnaXJfU1p4HgksYE/cfF5S3LLiuFl3oXvWxFLyethfWML7BVwJ/
Pyzrn58VP8k/j1/sGtGoVNagCiU8ziKbYsudhd/BqymFOHYlrQUEy+b/ikPjByXOnUU/LX48sR4F
LP/XF7xUZAU/6KDLT4f22xZSUdMO/rUDw4yGar6Mcn2IybclL0bGJW+L0BuiYQcYgco/gqZYl4qv
DoTyk7+KOGb/bXI+B2YgXZJsgS9P4zYU0qTSXsx/rwunHeXS5aAkGjXytfl5GoG9vARaRoOaoG0t
KrRv3zkZUAHSpLuAuAktbR8Pfs8hfMWsahyI/JLPJmTZjPVH4gsircVtj8mkVybJcG7/kIWS+sye
inUZgQmMWMEeIqpAh7tbX5sOEygCv7Yl/sM5+t5m62OzPuLnYiD9GtTK+FphIIMf5LgOeB6l7TvY
2qFkwrZfqU122zHNkw+L1qHTQ6qsMwwCq851DT/CsMAceIiVoQTZmsB76afNrzjsbskMkeIwkvI5
XyDYsLHJB/ccDMShOD6gUf/4mxsYE5qZPJPS+fm8lTplkNWQfhtf5BPQgmS6c5rkulRh9SS7B6RT
ECwerLlWDkmAtpvwCBj0xuyC4cvbxpucXSvubdnTARxzoJNGW302Het5cYX53TiG4vyBcN+H/L6w
UP6cEkCGdux5Za+khQld5Ty6kfQbhm976UvqBsC8AVjIuesMvY2AzTuhMhBa0r/eizkn629sgj2S
8xxBrGuxWGCATldFv6YhPKqhMKscVSrwZhaCuRjYuYjBcYsea+aeqg6JWuBD3as47Epx7aOsJDx3
g0T5WDI+FCXC9hRMRdWb7muBwyZqxM1CBRIqBfOOY8jfI/eYHlGjKIgGKXQz9KBEWOtbagkGZzZA
o5rM0LlkymgHU0jZmD06WvPMft+ysEXPMyvn787JiOpHG4yew665PlGFjg2vHWsyvJs6sQ6Zn/sW
lz/kthA5rXVg3HmukQ5hWmUi0BFfbPehft9OfubLYoTqJhGwiLU0wgrxYbyzbzkVArGotf0zKxhc
HJ7Cxvr6o7+vvT497x9NFh1sdgqI658lTsFCladjd55NAjMcdDpAKPuQ94e5h57NuLw9rgjzsvyW
hvj4fo1N+LillyzvGftsadtFmoz57SRDJW7YHTjASUbYVbj13zyFTV2k1M3LjyOjZsELCS7zrtwi
dXGhr7vfjl97dPK/Oo5NL3osnzfjl2D23jc+rqoM3dCC9RBSVq0ZyRW/N9SRMDqiWdSnnz+M96LX
5VRxN1wHkpvkgeHDSgMZc/Oe1VbyPRcLg5GFHABIKOssYDjtkTNfkxbP8+elWfM0uBsjpyHrwCIo
xzL0cLd2M7eRcjh8F/vxMouXegdBolcE2By40vc5AycESrQCrWokAufsbDhwLFG48K6hKOgVrqGc
urZK3UriDYpC1ZnPYZc813CsU7iPd8IEf3ZGlfG9t6eXV6Ew9gJ/WFb4Dz09VLB5RdqcLCbeJPgp
VIILEl3JYYbI7VrfvewSer7a1AwsmyDGilOaTUtfsbFutVvQFsRfdcI89PNJQIC4ok/hCrd6XTeX
Se01NKGEO5F+BiRjUZoS9VzFxagKkmj8cLVWSyCIb2h/7poxLWnscIsMwe07Md+AMqry+ujZWjoK
3sTKfBq31tDfg+HXG9SsU4VKE91EnFO9Rs2IXEEH3IS+8FFXO7IS37g4NZBnL6bcqGo8Gvt8RhYV
v9pFcMlYMgcbLXfcWjixQhtmAijPckhkNj8oTGawoA8NIYVpuj2B/qi8kqt0T4tENeScyEeMeBP1
yljHCrAD4dsZJbboewTQcHPy3pLg1hwQ4n+BImtlCCawUbPKSEtLHQ4/GjnJcy9tM0VppMUAQ4FB
MNxJkS2XLEmCczMj8BB3UJ8Fd09iCql4gb4xTWkZ2J2DRuNw2PG9mVuu1gn807jmK5Em2Fyl/Onq
hzZ4TVQF/7LIdDJarmsJ1mTjCmQLtg7LOYLQ35mDs1KFLzEIa7/DMN/xUH4mYGhhkXRhmGbNBfbn
pMOejS0tK+3U1rclaughO/W+uhf6UUDW0D8Ah/RUhJbCUUkV0RFiFwrEh0gF3TkrZ8LfJ35Y0chA
/2BE9jDzk6Xp1DaZKfy4jP8VLs9bQl9ijy/cR6oVJmaf2swLmBEXrKq5VcVInyOWrMDm4ATFmjg9
tt7H0iH11TS6TpLUEqGjtI61uItrHGlm09Tj7MAHwnF2aeZIZxtThVyld9+UzJ6en6jm97eC/K/9
ZJhQXdz25PDQTLgvDA/H4UH3fP2OAmGMsZGn79YHYDDUF5SswN/StktNs2mqz7fOFh1MCT6wsauf
WpKBj2jUp7P9Vl9MJs60xCRQgxCzj/4WhxnZTF9unZ6xgPDVQ2cOoWGZtjyvHzvjvJMgfX6zJxlr
1abBtlGkMn+r4nNIVoz2jgubDfFRDswrakyPdGuu+pl7gc3NjqlpMq2x1deLJ+ew0B/kRaVOOL3S
FPylRky1/bmZga06IUDltRlZU0JubQb4dMOk5YloIdQmIAmGkZd5WCwJvNU5zyFnh6ULVtgDkt6t
go/qMtXUup76rED/Shz9S+WDDJUOwlbzCHj7U7T5SnzvoGjEdyZy9ddNDJGaDkRMQSzSG7FE2iBZ
Ts8nOBLnzjtRPsNJe/nkMlqzwsInQ9rAorNDUhG/HEA4KOLXdldV0weqHyOLrKJEeBTDR18BQBKt
XNvLWVOSYGumsJgC8zHJ0hZDnBIIclRtuijbExL3zNtbBtTsjncV90I4ZsPhGY8dya0/t57jki36
pOWKfkN0rFKjuECZbb9tMytLrEVlxasJ9Xv7QOBtKx69N2oMIRMawuG7JQDIWOZgw01ukRUi6Fmj
2JY7f699gaCixgp7gp5F52ZUg5jz3FOS9LDuquQQtxQPbiUvWX2D6bKVPlFCx3UOR0koXAcZbpxU
Al1eJPuMa4cVmbGkz/pEGTg62udTyjTHugSsknysz1bRzC4IFkKthrK2hMx2PA0/pfDD0VkCVnc5
WkP8m4tJWjFwu5WAUa2eX72GTRtK1I+AhfmpFRVV1BJjya7NdAoFM9RCT63qdleLUnlmP+JbUhVX
cXCKfWFOooBgd1KEh0zzK9eunecYRBzJWOxxwZJYhCGnDGFTHWsbqjJ5V/NGg+SbWbyxK2ws19SV
GAqd7gwIlcWxQoQtsLLPlAIY/h8DJqASKTa2ffPmv9H0MDByoBM0AF5YuorUPqM2U5sqyP36lFf9
bnovmckFWb+tDNoxVEUdRDxDgV22DFMfGlbKH1AVfu/hQ9ABhM+GmhAA2RnNC89ep1cSzNM/5fPg
tka5ycmuLW7MBNQ7GptsF+5gW+EUiCIlkHCxG8hhY1tGOFBNHFayGbsg5dXRLxKxp00pOnjhBdfm
TKzyl3cxIsVO4jg/5NO83CzkPKYqBCUPkhdMBsNS5ZUkg9iDNy2/Ikc997/CVTiTnLqGjhDsP0pg
1d9i3f7ByIx9xMjLIoiOvyLIk/V2QQ4pfr1lfvzjjm/o/4hbX/RnRLrTTmNlXMeJJDm0c45zFTI6
DU9N2sPQ8509vV5GxQXe0WpssMVOSob86rpukco8Tm5fUPkfPRfGbrzrdQrVxjuSB7bhY9a4drOh
YhJze5HifjIO3OHEwx7vaQyZ0V+mH8WqOTpPD7pCTw3wGfumd9Q6S9lNS7QmRGm4R6bJ6XSvoR8c
XhorL4kulxSdpRql8WBvD2GTq5zWxox9qgfu0xBg/b7WmABJ809BvPcWdvAp+5i4EjE3w2OVpc/R
imqKvh8QltxQNquchYtpkoG8Vd/pRQOUErUaAFCHdVvLmt3xcaLm1730Z7K5GhglkhU3qp37acYb
s/RfxFm2WE5KzzmMJz2YcDi82WNpfSA82ZuwXjqAn3DEyQDSn4DT3GYmD8fqgtZrWSvyugfx6abO
lGCN38tJPG6QHwThGvCJH1tdq6rBc0Gn5wLlLCXeT+I4S/r2TMLcDXzh/SzM8MDRJ54d9PY3+45H
cGg+0aEfYkz9++dWuxHvGrzhHIwqxXIN7mHl7o9WHx5VltoDffG9sUWX+yw6bxCQyrpUGXvg9/+b
MRt69tzyivwUUJ0h1ZpdeqNale57ITehQVjpqQJ1OLgdNXGrthewbgCZ4fY7MfEVgf023nCn7sC8
jwW3WlY9NZVy3KEHOFCsB30LL05Nae2uGqpZse7AwGpG8Xsi5bRMOcywu2PWzpyuChOlPkwtUp8B
xFqw3qsridDXsgJown+zrYL/DvZzfc48o+x8/PvMhhhrxU86knVxtRlpydOxuGS+KAhqycjYkYty
1IOaM1FxbYYQWdZGlQlefFHv8tD+M++LA1HSvOVg32pNgW7uXsdOJ1G4Beoo/eHMvaVQvJlEe1fy
8PTlXR8hVUpdWaIjDL9tyymbT1iAGKGSbySB4/JMQsIRkkNeD9qjLijVpTHxIhHD+FpsoJzVuO6y
UIkcbjnK4FdtuN5fi3vlhPt8jzfoabimZg+3olTjKxND4AgAnCfbJrchjqdIZu3w+sg2/sxSOI/0
hKD1pv5BtvWBaM1gjV/0/sqZsGL4ZwxiEWaZ+5k4g2WE3uBc6YJ4e67i3DKGnwgWnOVS3+7tvU9s
wF5XIZKVP4gttcme8E4hEJW3yllWjgeNKvYd2AEs438oMPyoYutwpMwNfcfTfxHlO2vPUgEf2dGL
5OTwoQ1p+Ts5/IC3Limk+D8oCO6ZiEGEN3in7+Dr6e5qLacrcTPJcGYqbKbwVKGxDSEPWOkLwPCK
bkq0beMMSUw+UiRMeDEcwWmXR+XKxtSp4mK680jkdhUH31gYBb+W8e7r46pFRcQUxYSWlNF8sZL6
YFXi23Y1bDESj3m5XwPI0REfCMemldpYAv6oNmsgKKkz1ymrL3yrCxRqHG4ktyDHHm0dvK/cd8/h
/uB0wIvh7tBdc9DmMtYvN0NI/eo4a9ZKWq36gqgpM9Ery8iuEP5IY91oLHMGYJSwQelfkl3gkiRS
ilz9Vo+vHLfzM59xErDFZpJIiSYRR14EZJ36+eLFmvrWT+NtAqlMuBEmVBaz+IwwLZ1EXTbp2qPw
DXI7RoIfpRMMlyAFhvrVGdIl4v/iUE9PJ9S7niutZSC+saC/Qyv68ex8tZ71qK7w5+jq0n4qVxPy
bsZzCcReAmhpxbUqQJA4D1frIC+Q+jkmRDIGe+kG3UOFMO5ywpGqkZE/YLs2kJ8YGuHe9wM8JTTD
gPgVA2XOv4sj/LCAiiVBEbkcKOwDA8341tKX8SL2qEIhMpQRL3VDqd7bXlAvHLwxbcecfljbKCff
nNihfp9jrYNgvmDaAzck63oWAyU+75brOeAMLqdloUV94CPaum1zetNyqW7fNBZa8jAX8GVgq3uy
ksw0WRz57H0iWVdg3oy4t5XjuFGFvTExDvURrrHJNcNB1xnJogGP5YGxNz8XIVM+Psi9dloMyd1e
oVIvXGYP+5Yh1MVR0woY5O2vBabxKSYcqclMWnwBXd3do+ufUOJv+GOjzv2NBth4F1dAePXny+sG
oHRUFgCwBYh0/W1LjpWQ4RlM0ZVXO9A9qSzEMtxm4MZm8JUFJ3Jik3qFGVmXRKPYrZMiKI0ovaC1
nqkK9JP/JAChquwOM7MOwbzNoU0kLyJ/JB3/z/AAN1n7elHLyGlF8uP+Ha0+EIN4Qctqh9l7rxoX
p2cWozdyEOBEhcCRQ5PwCw1XyZQlMOWNQ8rQ26tqLID7tlUEGRLdSQLxi+Fa4MtJivZP4o65yytg
OclE30qSKVd7KWh6iEAtNWhYCqiL+1au1UeV9ly7kPkq9JRwQEeCIqeK8mITiX8J96UiAzqvhK8j
6Y0oUQacA+k/1ucy/DbqhcpaGNyjSUKf0q0BJZ6rUq9L1lDbMzW0gkGKdUXMqkSt/I3Y1uKPpZCh
pWeKpPLhLSJeesP+DyJGn7+2bWfC+9PiKodKh1jclBrSiNqXGPO0mxDd76FF0UAXu06J/RSFimtw
l7AmaO/G0u72HX2Jm71KT7b9nW6oFjWYtUlFV95btxh9W+ekh4+HOIZ35mBnFZKl9MyX0O6PCI6S
+qormAIeCcROo/03bBKTSE1Wf0+TrtEzVf0xwCqs3SyHwEF9NeFzy5uckCLSzeXmNtSIutUzS/5i
4L+faOcTiATMOQt0MZyc7QTcTMUS3WxKuJVtzFCiJbKMV5gwcVj53XEANq4EQ5APu966JsKevSGk
uWRV/qH3vHJXIZXdLhzN2DdJQDaRI+dFlLKxVaf3CdAhcU7IwNLIWxsD5qh6faaiBrVPOv3KJKUw
LO3LqDhOhyHqn7N7SUOU3ywJTOcymIcpToOipgn0l++lm63D9EKkx90mr4wmtM39BhlDQaq9t8sT
zk99QOrWkwALpi2BMCzmStBxIpsczxkMNUQRDJcR1oMFZhhswFpNKulBVtXRTzJGWT1e6j1FLF4M
8s9raH0gkH0oei7E05/azM2ld1ykXuBNuS0JUuy6hM9cmM907Q4sjj1Eh2gUc+Sflv5ipP8i23x+
9X2zSsvKrwtD3xQgb8WaAxfO4obRDM730MaqmjbtkANhEp8jKCYjDkUAU3ZB/Zlskb/wEiRTeiTa
6Wea6zQA39rM4QDLa5mHcL0BmpqSWHpFWkmucFgV6RiTxOFyXW7TguaLPhDN+NcJSAPUrUOwSOou
JQT1moL3pMewSjg6nz5pNResnJoeeT/x1wiH1LCPwesfOhov/CdOcjVSS6aRpw29tR7L9f5Blc/R
IaP9HJgI/5fYk/cQYsJj5A9AiESZU0JYKUwmfwv54iA+zGs7EzL3/vWXLtQJ+FElRNeRYHxaEsQA
LcTXZ1bpWa9cKaqHE6jAbJmlfkF72U6HoP/1dI/5P+ZdGBA0JnbpYZ6TEubK1OoeaGctTk1gaS9t
iGC4yj+tFzXKV0TQ0/B4LiA+GebesFUF2mVxpEh7KS4TyKwn3nZpvEgdCAJOzkul9+HBwH98logC
fEv/5E1aS0v1ejqrr5zSce9DJ2IS1KimQO112N19V5r1QDEKaZigXWpsGLpEYdf40Oqlppc4mZg0
IV0j0hiY3uGs6veOk7dsqV7+p/Qr4/4oADwVcyRj2toH5dw3XAGHYR/FnDucH2JDM0RWurxrp03g
RFWGN59XX6f5ymJx/uvxSvKFGUHLRIvH95LotGVDexHABj723sqlWslrxe5Nmmkg83Vl2HVVWGyN
D6vbhLfsqeP0Y24ta3WfaNjSjXNTOnUc/Xz2nJTkUg7xHhFN7BU0L0D5Rs4U37iT0iA0NPkmkgih
Q7s4MecNy2w7QZoex+4LC30KXGLVd1HfctWYsC59PnUQpFY3XRyMjMCMSZzGZN55/lWrTCPHuX92
KGl6t3A/nwefjupm8KMSFRJeiAwr8DLyoDC6iSw6y1vDRG/khFAltLN53rYehw9OEt9cp+gAM0E9
rjIXAdcDsnZqiXyK88jTSTQmaZsC2gqRwWpcly6F3J0gb+72umeki7bsK3HMDw6koaIa5ksESv6a
dO2Hkluv4/jGuScGpb0EghSi1kYr8XdXIHvkcl5Tjm1nYp8pf6krdceGjhySjj1OmZ0QvUJvUwmU
Go4yUrD8KaIvXFBO47FXpJEoPN86ao8aIh69klj0IGx1xrr1UhQ9WcgW2IH+UVUc3y3ceASm8Ej2
8jIDDVcexg1OAk0PlCvKO9Yh3EEVecdS+VNG2iksX+4lZP7//Xakw5ok646GSheCfacdAp8kbZ0o
N6+nM+foRiW4m/3E6f6rH+1EoM+0uZ7QBv3l1kgqhIgn0H6h1nRxWRxc0SEhyMHE1zZE9rFJjSZn
p81ZCHNuICh4ixS0rUP86GmBVG5Z9DMCvNkjRBW5fOb5bduV4ygVlHF8LJ0VLNEAZchH7GeB5nAV
ihrH7l0+0TnpSwZ/CuaCXBu6D1ZQK8rB/UCQHwwTHbh1huc6yzdYSq2Qkz0lZO2NE2sh2a2OgNXh
6iMo0xwaUOBiUSjJEJr7fLeORTt2elFUE+1EEl8+SQ4n0i8U1MCfzNvOMYSpl4W2EADX8RJXHjQx
cHDZuT+NzfQkL7QsJ5pTBZtKMgfkaxZ7vG+byP+kuK31gPFvYkrya9UnyMW+A2xI0NWRBNtWhN96
L9K4EJkBlfJV/+VMIRbUvvzKAEyaGR2eHzOVFihRSckPn7gE7n9iFfrJuT6jya9IPti+GhBstWew
zZwpL1OvisBzBr2kh5cIdzuGytyNs242g0f7qxKG5ZLwYCIEzKncK0pQtEey8XM+cw+XrVsfV63B
vjHwQ4LBj4yFX1DRS+Rf4PCF+d1JI9K2KVqlL7xWHdtkK4lcA4biNeu8hPNAo/oDMsNdV8Ye+SnQ
8NJ001rusmes9QAm3ExWRrnYmFpL6AZuyLHXl+l8pn0FuCgKDOYHnUWpS4vuu2q8GEH78otoJOiA
x2MY5qtFG0mGeZnH5iNTaOtZkacqBgjOlWGfF7846t2nstvJvW/wQHMdwA7C5RC4zDMVlLiseA0F
FWVEM3vpimVKd9NuFXeFcSiuj5THO6PjaewYj6BTVlx8UHGo/rUR8tGvvNZaB2hu/JvlIamN47ZB
0WVZEM6AFCCBGqZ0MMTAVN5WFC+yU8OVlooPmkJl5m/6dysTXRcDox56u2fW0U+elMj4ZQgYcBsT
YPA7LTCCxCc5xMaSimVW8jBeE/BbJWIHSZ3AmSy89gMDW0UQm94T5edpkss2Zj2jhtOoOT0DLxXZ
iZQTTzBhhF8z+9cqV3m69PElQAdoR3Hspg8MxQ1J1FASTRpyBv+Ru1odFtzJl6x/bANbH+RZg7DQ
cBHNfRKUWfsrdaz4FQP9y21f8hrMDRxQ9sKi56JQqyvCWXRmZC1bFYpZl9ScNM1DYZ1NeOVKYg0T
1WtZ0UmN+H2/hsCZ76rV9tmdRpljccfbTnjMupWIvDTaAPkcdRSch3bewprHGzheNtejrY97Gfsu
NnPfb/F7BjN2GQTj0A8vsMFLoeAujGAjDc2IBpdmwplhqb0yezyE44mH9g9PhPEJ7Uo5DOD6GnNZ
SaITlHKpjT5GsLFVRin2KNz+xWfoDba9lYJTQh4JUsFc6CooFyg4sn6wNbh64yzOWOfR1jTF92jZ
CdLO17mUpXtI2n+G5iVY6iMLV2LzB2IhU+20lfIWCjazkCz7/kMdtS5suJmV17WV1qFE+DRbXwiK
9evK7hjB96JAyUVeQUrpHD2B6aEuDHpqYJ6O1xxc8MXqpmv/TaYur/ORntM4AxQeQ+dpk9zgxJxx
FFhSy4F/7DWHbiCDMS/7gypq5u5tXZAoZ8D0s6/26X8d3zn1/PqhrQDohUe+W2ZF7pcpralVkp4x
0nBxR5H2CRaxar17Mt1FDk1vW02hMYiyfVJfbmIDI+obideoDsHZrw81++LVLRbQmfrfS5TckJ0G
DyiZG4hmnepVnPpEnZDg8OrPJHlZ/1iPSHjfyo7aLPTH51gPkAqdGOESoDIxV+Wmtt/8ajY9c26B
MnkCyILGn3DZ8086KeVtuwEdTd27I/vkMxtkROn/TH6zv/7/AmPjRATgJBWM+IDAhFGOZiJwbBj/
4HnmXsMeFSs0Ote80sfCpT8q08uQq57WQaRfrtcvOdQwId8wFem1/Dlzrke5rhre1HU53W+0Wyll
IgcXhfwd8/yqrTj13Oz7tvsH3TWM8oeGlBWRgp6fClc+Q5+6JAHMZMZrjkviKJQPRh4ae9kfHky7
AJm7p7uxMmNLsUUn372FcVuLDq7nr1V4kOz8ieSHh3gP3bAKH6czuD0eDcuOGlZbhZS4PhVZH2S/
E1n1caVdAqRI9eJhMwT88v+NgJsQd/khXiyjLCP5tLQP6tUO87APwGj+vMUOiFhoBPy634PnCBpI
riTCUgW6mWaNeqvicwpLO1+qFAWhXBfYcKYmwvaF+22dqiYsvbi6jCqT82pRvB6yDHwBTtTvyh+D
G6NRmy6LpOzCW7y7yc6LB9BmtiVEaQlFPPqD10kNLiE39OPz9+w9MlPjzCGgvyFwS/GA6uRmcofV
alLSlMI9Z62avxkvQdspmjpwN/Udv7E9WaSy4BInAVWC4bF19O0+VlFDTpK670REyYO2AKTrIoyM
o9d7pcCaa+ZIxIV0AaEtYc+vj4QKq31QAoo0/pjAQRc2z1eImv5fmVScE4RMO3Jhm8J8bLoSfQ4p
XQG8DtHea2hy+BIUdxuWKsVCc4j4A6H3u/60Z5tLPCKT6ur/KeQ+v/9URMC2G4sKUS3Mwbs2hgIb
yoES4XrcUZuksJhs+bcqsTwUQ/QoxhZmu6Hr1a3j5tXrRxjznYlix8+itDrKJBlZ0m93mMX+p4Ri
ThU7+/z3mK+4tTkF/dcbexKmYjTfDDUj+7/SY+4VDBkqJWbZxpyKaYr7gn67/SvRO1ksgUvyjQzo
cDYEeeFNY/mDQIo+PqXGE7yDrUJn7wlEW2NhrCheQV2FoFS2oi6gUaF7SVoSYGeagLZeBBTNhkDD
4rACxqQYEPAz0gYTuEuuRdGsfBaie1BUiQoyi9hm2nr9B7PP/ghICfhJLWEbUPABh79xOp66JllD
Ix49275koGvAYdX8o3Dh6x0eTUL0b8HgjE+0w1JFyaFKOvTdm9d6LbkQbbART8QG2Gj2E52iAvCl
ywc5ZBvFLcXb9TSzuYpJUlLC/BbwRYhop6hAoiG15IWm7xuYJtojBszV/cbkHrXO9Iwvrp7m0tdg
hgRrhWvqSdDVsfxFzXhZHO+g12ESRFW4aRsVzFolxQX8kJuCOQJFq3mtyFq0Hw2WuYIadrfaVatL
RE4WlVUE24yld8/Epw59oOe5dxNKVwUGxMNWiYuqIyDIaVZi6EFsY80kKsskE1dToRi5iCKGzpzj
VMTZRu3XJAE5CWDebNpHg464/aole+j+MyGzXBXEpAQDvlR7BOK8PuiZsOde+D8IF/h9DdcdDpSN
JadFBeotESxO2Ldar3n9juim4lbyJ5H3qRxbL8NJUfEzhNgQckC0zE//zF+9kxSk6/gj8WYrJfZB
7kwAAie8o6JG2958kQO/pXmMg2nQ1vmZIRy8U4RgnX3YjZ4BPdqjyIdbQfxVM4o32AyDslCXudW6
BNVC/zXbDNxRH9MCUu57Jp2EEAUjUk3Wa+RdTl2BhFNw1kl0+tNWRwi9WQTB9TuTc2WXICxz9NQz
QnfdOhl5jleLZQ6eQFqQ2nv7ShBYcpL9gSZ2KG0+3E7p2d+coprbk3sv7DeQynDjRFVJLQgpkvHf
ckBb+ogCineozAo9J+ZzEkg7NVzkXdzNW4vS3qUURu3wNoNQ7sgjKcCluzBcSP2spG4anUbFPp5p
2mFmdq/5Y2ghwaDM3Lef6XEqd43BkBuSsO9DqMkw06o72JqJ4qPSDBDUjS4DWhtqK7r5plnY0Abz
lXCSo18Bo0Qo1s1u7l8qlSx1HZ8T7Qf/UO7bCE7I3IWWiy/rymgltiDNabdwr+Ordw4bFo36Zi3s
DhyIrxtjlMPRBhbU98bNcHU1AqCa5p42Qq2eB4sVMi3fHcV15Gp+VRNv2TMFWELM8fPNK50J+z7b
qjklNaEMB+XDKyxvUqNzHffR26j15c6Vu0Tyeigil2BBsN3SN1kGK1GXaj7XLPoMI6eepe5l/uS/
2+imP25VWSR/mWVp1HcI+diLwMXZFP00JG5+q3T33KOBWCsLtC950i2m9DweMclwiDlRnRSz8csm
ekTYCVKC1UpSs79ZUBy25bJbAsyVdt+qXYIrWFWcRSGmq/7XeZAKOn1G5s37Sfx4MGvV0QcE7wJT
5xeyBT8JjEIfTYNvddS8QRfhsCaudC9PEXh+qh1L7eC5Ve5t5xjJUvHGknttWnQVPPBnd1grJRJ4
omSsBCg34POBmmyU5AT8p7x9uEpJvuGLvHqpuifcRSIEoEebIXDHwMoB8f7KME+STWfynCdicJut
3IEwzVw39iuuNUn0Ll6uMOPWjBMybZeqSPdE1b25r/IgA67gkbWyCfxhZdtgbZTvkO2LlLTxIARX
k2BYdTAb/uBDykRwkInQmNPJ2jh+GxcKOI475LmfpFOveNCC2rty0mjh9yuUDG90D4a42W1K0XzX
3eWr/jpgyaf7on5GYisp9QXepYPMtCbiWOxcTfxWJAnpTiGiKun6PFZqtvie8jogqctulF4QKLZm
7kb6m2UEpws7qR/Mk8fuO6RuqcpcswtYomzqo0k/pygSgd4HLe1HgHKp4rz9t/RfjmLPY/xwP0kJ
ghqbeoo1oOXF+wiNLe7YOg3g7ZIPY5n1aSthL2D6F499VYanVf1TwWTWxIWb37Xq9fbZtNxVueYU
H/wo3igMPILkevwVYVZRawBcjegx+cgAZh5072cjeBcij8USYRc5s10hxa1qLNdhDI4Acu3DwYml
n306/QzaALCMSdEm6aN8JIarBV1bCYGtH6W+NskHcasnqralBu4CAnC86E/s56/SMNm8VaOnGEZ7
0bnoDr56SuKzPhIkxWzyMXNqraT46wJoJVadLYyhi9kJR5kctn/aJCibk9N5zcYW0u45JFRlHExC
/6Xv0/zYkWtCKk24gXBl+xKxFy5h+8kWv/hgonVbmJg+kGYnnd/XzDpN7fXTPoP6utNwZxkGfWWZ
skdOolduC2tdNe/GJLkAMC82mwenz5upchmeVmRXbIzgIzUY7JZRlMirAyRujDyIq4tvddRIka/5
J+2PVbUxFFSGiDOSVxAi8PUKF3uCrGzygQYDXE72ToA5YHtTgCMQRr6pQv7h0AhDpxvhjrZXcpdH
uk9TWTZ0mhnkeQCB9W81aat0IpoBotP5qA01nCCeuMqrCmQV2GYmFJ8rcevmLyxePNbdJBphwFOx
97E8zTkhOQxh6yn0UmK5m6roPqNfICcyzJOP619OCXztA9yiluXQz4V+425/8Z9u11iUpcO1ddTM
vssk9sKOSzi4CX9F4j7b/ynZIhxwNaOob5m78HllzRmnW8/HrDB47OVwPbm7INCMYgqxNqrBY0g0
syxgeflE3XP0RQgLXmK42U93x5cwiUiH1/Ao/YtjPD/NWEhPlReb+oyuQxNaAJv08gLPOOkbYXEA
y/TprWDvTS1wnwqyES31DvI7IBtbSrErWB5f1Az1Zwu9mNecleUt7Nr7Cp3Jb6nmn+sAVnceAchN
uLaxgkaQAS/+R3PyUdmHxJ7VHxv+GyxajzUSuD9zgJAAhmlbi+WMJ42QAsqW9WccVLI8Ehvz1KJM
r2hH4LzLPTT0Ew2TAcWvTd/01u6/pGQ6WEOZH6026+ztabahuc5gz2r9mBixjdcHq8cfgEp729Tl
KmxstIA6DYm48PSyH62BLKRcs2w3w4zkxJLLbkqxSt5rVHH+g2zav7HbQx8E3kdnhhG+tp3+c9Po
VfSaYZKXEEfrBEpomMCuUmNwR9quNiUKFmchFATSd0+dScjz2GrTdYAbfmwrgxqaUgstBjlSLlW4
eYhK/o+dW1oMmJxxurLyWu6Vtk10IiaS9/FrA9MzdMDtH8JYuIYK89GznmxLMapQ0iuF80NbCO1s
4zQy/jy4Oq9IG0Lsw+PCYm8cYx/1DNBEiurFON3xec7QjVqtI7ZtpoRnWQjpzScG0fA+6NNVtGdT
b5p4g2KfNGDBENAs+52qFll16zOmnFlshEUnAiG4pbbmbslWymtCh2AX+ojBidQkfYcXMu7eCDFq
gXJI73l7+7oqwJGrJecs73321/U8bf9Pi9+wJisko9BKrX22pG98ZlC5GpcVoge157LiL+hf4GQu
kgadVFJ4uHrG9E4N1gvKss+IA4LOg/hYQUxs10juuUKF+38N/36aH7CpRYYYN5HZ5+I2Fqqhe4Ti
icDyDOEH4O8X2Oh2zUmSqUtn3Tld43UB0hCwxr2rmxeD/IEoekniC57jx+8khC9JpyQeXi7PaXBU
8nhagwl0o/eguBaCnMzA9j8xWaZmD10ZBPgJj+EEuAU+15nkpI1JNzlYtz6cDntSBqefvLFmpGH1
dwiAJZqsAehCLsMITJupwMOM3yQSEGQRW3e1k7oz1ie6aadDsL/4XGUt9Eb3LGdv9HxxPGFpEZzt
zB7hAF3GWxZCGwedW0okBl5m1TBAeoRAICuMSF3y90xEl1a+clgSG9ci8b7tqJNuB1dAL8vnRoD9
xL8/xx+GBmp6ljWnNooObu3Fy9vpY9zEkmG8nsMIFOy7q6YRMb3XTQODwMMTlwnF5TNzF9RC0zb/
GFjLlOXlUPNX1mAUCEz7VrH7mzA22vxRmERxG/eEoq0Nmt4SCq8FkB15Gx+Z+x6ho51PAfnRgtSH
lhj/q8VtyqB4j0u1xICIveMsejhxkzZNf/8VtW9pZX8WTKcNBuw+MNsN7TP3JsYLh30qik2r9kHw
G6cDCWqK5z3Y72Vc7cu+jitp2d4UjpMkon/iH8KY1aVZGu9BN0coryt19XvI2Ya0N/1BoPCIstJ+
Gvt+OsPmBv9+84yDhe2iLJIyrW2gL0R3nIFArQ2maG3WHirn0wxnYfvX/55W3IufqEMHeGwE547g
zexZ9s7Iekht1vVTW7bpPKb0RLAk5B23FEnA1qk34NanTMu7Un1YawuAnE2vezBIJDUn9NiUkpGJ
EUNLLxkzzKtQAYiS4VL8s4QUsKQgLvM4+vx6uOUG4dQm9O0D37rmCjx/yFfz8fjKwWNNZKJPsnRO
u4uaWq8kO/QLfDoPrk82JcwJP/AZpkCcXQ1H7hOjblq9pGg0IyExiIYSPThJJ+9HksHOiJFmJb94
D8fNNGnEMRIApit/eIOiJhxroUDsEiDMTMR67xGAmIXLpJ2BZUNi40F4It5bd7aNY7Jzo0EyN4Ag
hc7aNl3+Pd8p07LKzvGr8ftfDcvYKsty8h1upziB6j/tYfnXcQrMAJYGXidtljHjZXFh7weY5vr2
fKiIMwjkDnEzhMIN/+QqAvP7srBbWIMXoIKBx8tRXBwS2klrFsETB65F2TlGDp3IyIBAKCsdgkBQ
w9xZH8JGXZGXTTXYHCGKi48Ub0gUM5yuK+TRhhxIO8klPndE72UOrQ+05eLRIVH22qB82l3rKIyB
Q9Id30x2wIl/Q3BMwLgtowdHHlYWt7wVmZeDMiBtAu7gTSUxqhKc4uxtIxMJ7g7bvTUSa+m+S5EX
SPB6bjh8zPpU0Fd+rQx6WhHB0iZ+17xkK/ocWiGp4GdFY6wBFwvjrzPOYSaIKYhUaOPFJnFASQw3
t0FQ6gpeZneXE0F9gjjemxlvopW952qRO5m4iN0uAeLx95afKtP62eWZbEhk2eiebF3gfNSrkBt7
up47Lk0huoB/BIIurcx9ty21QhHPPOgEAjr72iNVm6elKGOF2ITLUmU/rqbX0rLWC8j9aI0FhpSM
4M1Q286OMq+dzQzhTgyzf9M6P+RVtf2j8UCHrR97o0NuKRb3uOLQ84bixmCnaRGpQ9SUaVQjciR2
JCS0Q4YFBsFxNCC6EseHLVMkdGxXqhZGohD6ZdjxRzLjTKo+HPfaM8Zlfg7REEr7cVxagsWSoWdd
75rKbO434/ZPSBXY8zbBnm1CQxWi8FiPMvU8TPzVJYdrQcEzNL/3Pk3QMHMdZt7vhUU5OpX20+I0
XKeGQUDSY86Ni56BynoEOkf6YPICZ188YRaOm1wX8NvDO45RaQyJZU3utuvXm/idf0/1wdVv+610
8UdvpostbGEamnMZ9MsxKYyampOxharmE2wFIqu/zV0i70k2UwEQAUpPuln5etUCPAV2SblMJSJf
UVKqJCgSxu4o4hjjHvo7dPHLuAeWYDNNN0tcWunrJ0BjFYguqAdwVGKAyCqQdLGyck9nEKwOVRKG
+tzGlOIGvcSfsEc7uPi5UYxvg9vss6Y9pF8CJAVW/LpL0JT1+iyVH76QByaf6cNv/Qd07hsJ6HxO
NsfEFr20p1N0RCURzItLJzDArqIg+NlYQPK3Ie8G7vPGVRmdA+F1VxAn2ZAJgC91bfFROmYQhWHB
er2HskIItzo6Tgl3BzjCaQNGfwitIB39jyp542ngj27c7B49kIHSM55x89hQO/W0fpmRJv6ky9Kb
8cskuDNzYVIKY1vVsyQnhlCdEJ5pXdwyovVTsO3h2FdhxfEsn7VPArOyVTQAMCqgtfwTJ2r68k2g
zuL2QxO2qTEGuLRQ7tNXIWgNJjTrCN5YOaUdH1zR4/KiKRLOS+3idopruU0H3XihwRxMq2OemJuI
0BNutVjmsOJ4v8foAmDR0QXoiq6VSJg2/JU1pINA5Z0XlNAbnrh4kUxlXKPzk34bX509TAnyzO86
59x8QPMMFwmuHZOFjZ16a3zNd0qRTHWvZh9lgJGl4zCJaDrsCnlrjbNEboPeaBE3Z5ECHuNwOQNB
5mrt6NPKBT8Hzzz6Xum5m92Zjp921dbrdf3r1pnFnXYHZBBYSfzFuT8N8OxSp4RhVYRm0Y1BtA4j
VWjiI3GTo95RtYl0IABU9236Q0nd3YKnE50DkFY3De1p5D0UONQLRnYbdzKxIkLu/Tot/9yGpD3k
HN2p6ll7J8LjBryy/WxOpO1dRDCi8Hqe+f7r3bVv1Nx1I1xhJqsgdjaQ+MXBVJlg+CxoIXzEsaKd
4MzXjCLbhceEOMjoBsOVj2MMJLelEoBv4WL3VoWkXDKe1BqSpnoQd9aPDwddSyqdfdsiKpydsl5x
VttXy7Zrt3RqK5FTEdf/K2Jh7chRo9slgMF3uMqOU3m6PZFLHgB3vILmalMd7WUWiVCp2WRU/TAO
vnDpJmXKrZh19TaVc4NciQG6JjPgg+CNJ3qVRnxQJu5k0lzTiNby0HNSyZVvRK/LPUXi8i4HPOFu
sIYDhrnOVRekVO9x34pzAF1V86ODh1jO6xigMR3Z34S/+ed6woXNQ+ThoOqMUf7umeUKDZgFTDpO
jqfNJxpgP6lb85/cq6gT+9hCHwaPV2klKlVxgg5WzOQ/Swb1fdcdakyN/U5kU3IADNff1IG2SnZx
0AAHNEu9CPjOyiWTdqI2zSOD8JvkgqOKfMVGZ8qycwQEFHJn7n3SD9wctMuBCe1GN78w8EXNxcQm
3Kild8LTF7kIe4MlwY6DmAR313Hj58CeriOCXPEjetjbh5mFb/IQZSYuWza76iJlN/daX5ZT63XK
SilP58lJhpk0h1Ns54EXxfoihRBOfUFi3A+ZcFrUaeeZnUgULkUXpaqlIn7dbYbdVcr9eTJ/hck/
MgYF4tib8ss/4N5LghcKvUQulgGg3Z89qmLsA4NiPuip3tX5uIdO+fsB7j2oDjk1c+Zxz9nf4J+W
G9ojR3DtyB/ice51hBKDVn+oznHcBSpWq0eWnWgJU8XbmAj6uIsvTi2KLagmdedbXvVMa2A/FQHF
2YbnVf/vfFmOipTOP6KojVBr4FSPDe4RxTIy7LTopxzTlnLewVEKnT3oLW5QVzxD7tK+BYb3pa3x
gx2Qpk+Bx3oD0m/Bo0A9OMGIE4lGGXLrOfk+37YhWeSWomdvBqzTe169l38SVjqtY6kjxPUDTNM6
+vkXVKDkBr6RQgzCMpQ47mqOnYYGVKaTl0nnMH/CcHy4I5xrFHwSNBYpXIwluHPPF+YL/Qycpe+w
IaLBS1Vlb1nk6+jvdUJLTRdItoL6pVRLx0grhYXnlLgOXUTjmdYE96zrE3LJwpoSKVwja7Cl39xA
7U09Zc86+jTTB7DctHnDLAZsjjJHu1/YMR6soqFa2aGVdZXmj3d+A+lLztKCL0NuG4Mr5Xqks+5q
Sj0lL+XSW3A0dCDs18HUYoB0ccS33A5KO7ihvZ2zKPsph7DTB+O0d5T/GqU3kKhCJ0zRNBMx8ysy
lDfRpjYpGuWshz8XjidoIb/f/O1f/22HrndhrwL0IqNn9E4rIY4laXEJTd9fKp9RA5FaPFGS3wmR
RWFFIoxr/6j7lEDmFalm16da6sPWGQxZseWLffMz8ai7Jnce9AgsapSXta7E0NAfLQOKo2IS+OOg
ZQfE5Ile02wUI7+XtwNURM1+tuBxhuqLJt4iDbgT3+KhC0dnBAGjo3QrV8HJfYT3Trk2CKMFvS47
qaTviIrX+1Xu8+gJJ9I2/M+n5Fweu8Bb22r8EqsBXSaNLbdKmn9yhm37Z18vKGe3qq6MBtu96VcC
kMWk/LzdXtReSJtJTPamB7fMPSae4/OXPzJVfZK3llNXqbw+vuNykNFBGhGO5ecD2XPw9wRysAhS
KYLd14wMo3iF2+o6WdsGgNU92rsTmVZOyyUu8teGiKmUeeDVa6g33Ufow6ikId1dnvu3Bhqugisg
uCNp91zE9KH7V1XVc9dSufMAk2M3xckcpmk0QE4G5mGysrFgk5q2BVV7THDo7WpqCyOb6LxYwDYZ
HiDC5+7v99Pu+rJUb5jO1/4Zk9IoKbOtaCrlx7x7iS52oSJBew05oidwbx/WG6EG2YR0Y61KQAfG
qYQLRYmivadQnhEEpMvmKklabUi52xoaH3rOOkvann3a2gff68+3oGBao666QL3FSyonN8DwCz/H
jdUeEoGnWY9Mwivrh81jM4NOZV5OglCBbrbi5xz2kNlt2VcJ/48XNqYktC8U6QN1KcaDbMzO4a2T
edbH9l5Qsye8nQAAgTMwTiRkte3bDd3/z8FvsTItHpy/n6X0dKqlz1TIbk9X+7ieMNKaRgviG3g3
omC0TbfJWaWok+xsAehRMBzAGQ74kA63Y4SoftcBjPfT1PG8jLDwhoC5jH5MUqUxzAG00Ql/ABzv
HW4plQMBog1+mpvJs3IvrHwINsh0etc8UdxK07M9rZlDOhg/p5dbnxIe5DfBZ3JRUEnpiPieUMa7
xN/XtN0NqwBcJhKtjPYXQAlgBW96+6Qyh+pP5x0E33m+6Eujl9MAo/gDJgj7DP7KQ5PuAKzoZINx
UqHN50pQp3mGP/rbkgWGR1I9Z3tcalVpzcBlISCf5ODplO0x3rjTAYEKpq+afHoQRBtH+A3D4ZAV
9fuUuJCFyRCJUYOyB3rYgQ2z7aJSdREb2A0yUQLSqxG2pqRKHmBBbm5c10oJkdIH1nQRrpAPVpTk
md/eBnqvoZz8YWUfEHIx1eb37Q8PkEcgCnSdce0uufvafVxuiL7pTUTAX/AbmOmtMcSimr6b+S0H
Ufo7vXk5Vt2gUpsTqIb5XZkwafwSMgTcToV/JWbzQSUqxXOOEWvyNbj9T2H2ebmoM2MjIfqcswgt
yJItsUOc1uE/o+EA4uyeDH1Q3ixhM0yqy9syroy2g2xBsZygwxrbm+UDic05Yq9HqzjFna3o5APH
LZ1O/TxSFP+ZCqyj5uwOctJqbAlIoB35lxsx9P5N2Q2S5bINqcy25lPgOw9b0m/Ziq7cYaFWNZET
j9X35B3AR3JG3WhfgvsJAUEp0SJhMXqFhm3PJMVy2hhhIEAt3a0mqSyQBuXdc97l76MZIy0xKJRz
8mb2pZRZ/KR0+g1rR5aoWbFuf2E480uqMMDLOavuGpFIQmeRX/w8n4xbgBXGEC5P7UeRNRbP8j4N
kYotgHz/OC8K7d5SZwLW136jNPZxEfgq8vEpNDFvO3q3pOFkt2ilk1hD/rbt61AjD2BV6wBn9NH6
oO2nYi/uAk6pSelkYBqEDhdAMeDS/stEPQ/JH2jR8cRhBmcuaD53QTEopzlYrIJnyRx6nbLlbNe8
0A0z7SOs/sm+L0Imzv6mfBBr8djWLHBTbGBUx86anME4zJmnjOjuhvLIPp2r+rkoc0qS/Yttc7zW
zHN2aHYPcUg3Uo5Ubgzayg3SVgbP0h7v8IaE6tgyRTgh7Ed5pq+EKtdvOEXgOdJS4l6EQNXbYuD4
0th1AIfb2cL5wLmB0ER3qN1aBm+lV1unny3FanSfXpLiIdsTalvuI3Pqx2xEjb93OoywkdHDm98/
F2PwQi6tep3o3h5YSof4HDUGpaqrgseSbl9jJUVk3coSAgIOLOX2MkcrO5TnMqUFspieqsJZXAz7
Zg9tOFd2ICzcxLSa2ckHO4mfLU7c/1QwOw0zbuUjgRbHGfx21VyuoBpaK9qoU6iFwzsrjigFRTBW
Nurv2BsPKm+e+xidlZQYGxfIi8glmM9vf19EyfwD6NEibsLWV8Iv19GuFRkmL4TBBUXSUCZ7RtRE
K3DQyFmkL397EaTw3EbVy5OVz0nU3uanRt9GBdqeicdeBKgZadIUdrUfa4nvFt54lQj0Wbb1L0pq
hDQOvXoY6blR5sMRu6YZ+b5u5OsGm4TzMjchZ9wowKegHPvsE//HgAOig0AhYc2rT6blC6zArZIZ
/1s8pUlO7EfQj140VR6+VGn9Px3gkTC3Zy012fQW5vjXZOa511PPz61WwDspvwXnzHiiKY0c1ysm
YjfQSEw+8hapofOQFbjws1TEM5x8l9CfiEHwn8aIpUaKPKEOc7PBEUUIUR1D9OrV4/NbW/yOGzH/
P+Nx+VqcTV0Lr+MoazeTYSfeNN69xXvOYWo5GyAkws0sOt/LVuf8Cgt1DZWwCG0fyWqJTEc1Zg8T
3oQyPxcdpAAAeYfW9TZnfMoFSWmtwBsOfE9OLIX5/1C+C6tvx5bWhKCJLxOykuL1n6Pxu2/o7s+J
I+yzb0NNg0MMjn+Db67TNh5AJnrqD5uPJpH38Z+/Z406bBox65u+nOfh5zq4Nxy48NaifIRkmLsB
yn2077Y4Z4lUSJ/M801w2m1MWAWkixXbZCycywk8L805ghzxJXCAx4OUz7xckLxVwNWP4ssE6gMK
Jhig9Ta5FyW1pR2VE0yOjqe7wib/wlVEGcJLrRyiiv2AZ+wQqy02PueOVoLMf2KNsmVWfSteKgLB
9M03Nbo5WgnVjRDU8QTD9zzEPOnan7BCtGHfGQCNWgnumNl6fb24iuOzryZPVbiAZdGYJejbokAR
MY5hOFiqSTU/MZIzuDiJMPg/hwVF6sAVbVNuaaAf87X8CMRAEvYFaw0q6/dgVmWlYhlHhwptC2nA
hIHmT2wYf1HKjyk4YLy4HoABf3zZ4ea/N/vF0K6LLfHTfdlwh8HVANgWTUVPUZ5epa3J1oNN3KaC
tpb+S8gy+IZB+Q7WY+6sUzsCgXZGuTD3DLFHIkvsgw3PWdD1GMaAeUH80SFuB98niBX6PTGXGIac
vkPzOwizWTNV1ZvexBW0P4RZNa/063s/m/bORk5UriJ5N1kQYBkmP4sEg6k/9Y6jyS6MA1Ro/PRh
Z4RQu+Gu+5yMgu2fXG1mAMi/oRla8c7e2abm8xNB+zeStuvILVtFytOpUX53tE2FkLCO3+9alFEC
owVpPG/ZeAmPydHlylWIS1u29sZgBtc5JASmOx6uQhDBwYOwEoxXx0q4ctjLjKPsqTdSBAfeKxP7
0Wz6GT03FbdMJK3+MsZBiGUWwROEV0UMcF/0nxsSFcj76uxOLCf87dVrKWrivKzGb9I4qoFiQPkn
PX8pTjHH11lu7wVhsWgIl6dMDKWB1M5edRS0UDxh/+dbWhYGcI8u6C2RRtkqX/oAsrQs1y1tQMyj
7da52M/9eok3prJoStglPpEMJfwNzyBnkG2o2AU7gCw63YBqvjihbRzfJdFM1xIf0Yaw/1/lXJQn
KjENRjwowDataVUQ7jZeienLbY5H/cpN/wexHqAimCtFQp5MSpQcHYyoPU9P4kVsILbKnf2Ccbm5
8Qr0uS5X7PrVP5SAxVFEyVHFLLGU+8cfLUOyC1IVThYioO7lPplM1TCFRfguqABP0CUbMeFqjrAK
NW3aZuHfcUOZogYLcpJhLXQm/tfE5KgErzoNjgx8npqLmxAQkeUk1tZgLDMDaDkQqLjNho2yFf62
lZ8Tw0I1FpJqpZATAvytoK2BxRExXpAcApqovErSQiV99Qh2PYfOtxxpEMZDdJ/d6NMqGLqG9FFG
Q/phsYqBk3Y/1XYteLbwEC+89eLetCpoNZ8M5GSztcoQ3/WJ0WZcmW51Af5JE0qFQPVK0FAD+TXk
y2ay3FqZMhJ2coTPRSn/C8dwYEDMaX7ZjJG3CQEZvrQXi9jVHSeXTwHWFck2xtj6RZrw0Lu2NY3u
17TmjTiiySosu86QqFDcLOEY/qQE+RkW/dK1P+8Am/SfZ0a/UnCoBCajiNYYOeFpWbG4LlKHn5CX
1HbrSoWSMtymv1EmbRiSfDrkt1urBPxtzoQQ1oaqWFyA1SA5Ay3egGw7UWSUA4N18OmIhBmYeCV6
Fps+nf7xyfF5UUp2SzALc39jfXp44RGGvSKjv8o43EMWLvETO18YQqP0EoMyDId7QxN3aocEthK+
aIk1AViofXO8ROQB3gfuFs/B5hqgcIeBClmF/8NV2Ee1QCLsaIYsSKlb3mJrA/NisgoPsrc+yXY7
d7nDR+7wMmUaGvrj3Da154FUTapblwEVg+ubkpYLdMuZ5Lhr4Jhw9Ucvcu8v3Be1n961jyXvDq/d
aOtz2f575gGfhW9G8+26saxbI9L8sCUnnBBrycyXHZzGckUHdCEia+TxfZd1fuYDmYdKFlMZNjO7
27wpl5HMDtfiRzEUFfxfxzuhtRQwqOIi/u8OoV0Vd37851qBe8NVpBgy5adWrJs53cAN/na6ggvh
wrzqO56A+DauuMwBObuSAtShCGkLbfLfINmg7p0O7+WQDFGu4gBFE+6h067+ifQRhiof6azjlPZW
+NbOBff0letOz7phFTmQOV5iEScf6QG4Q2Nnbted9gwd8jmZm0VZrnp8Dsu692mktjoNW69Kkev/
95O05RGusOoChfNjbt6FVNzTe1SjdJzTvcJvx/mG9mP01YTADgsbG4M7fWjcOJU7/HD/yxobNo3a
VPZxyYmT7YInFGlXlM5hi0seRVzwKlqvNbyksIA8EcSIMbfG0g19YwlKKRTvHiYcWHCHzrF/cMGZ
3iIvfkIvQi8FwZ002ORaNny3wuWjBQgoN+IIAYl4ricPEWtH3I68jdK95T7U+76B9VyWaLeooQh1
EhCcBs7E74bXo5efvnKzaV4q0nvBBLQoFGtlLEeIjA4M4c/wn7bGdS0Yak0qcU1r8ZJYmXkPMKOv
sOPHFg4tLJebs4XzHXNFiyQ6ES28/jBatYdFEynF6pIOCR7pEvo449SxeMCwsQZcDL5u8JbptadK
9b860lVXGdeWVgfxzoWHhjo0FYp87ezpp0ZfRR5mF3vfbq2XqZgwSOAHMtcyoqqYDS7Cyz309HIU
ytBU6XWYHNV/SJQmJkGoh2D+54GqA6qreV/p4k5gtgjVha32yVXwzT/PVje9WTwGjk1Eqs2ppRaJ
iBDE1UXUKjCP1JTIYThLRRvTfgpS9SFiFDSXLT5AyBT3GMp1xbKeKtv5Sh00j/GwemSzvf8fzL9y
yxng3ouJmw8hyW6Cb2OpsAFIbO3UqWenlNK2wotYeV7y9G/8zhztscZL/k7bOQ5hToJbX7eO5CcM
B8Ozx5+A70YIMWgGTSaUT2UcM/EJfR5CieafLt7+3qbsZIWHw124Ljy1RcZ4nDt8I4iSbEKitjve
UECxbwRfHxBeGlNpYOQp7xxixHoUJgWjgqZf333GJJ3LW1Sm1tK1YHz0yRAyEVxcgwY3k8+Lkpdi
sFIplBt7n6bjkev+XRJbyqlvuACNVZ4Lrr7GfyxDSZ2ItKOvDmol/NKltX+SV7fRr/uDJUT6cIJd
PnM1dZXm6dBNBJLs4QY6aEtsXjjaKuneBv4xWR7BFmjoy/Y2XkPHvMqYwpZcLNj9fEszllfsgF1p
zHM6SUlfuqWnmEudWhY42RdgZWN9OGXvkbeXwiqOyiXzH53hfY+esH1cDFttKGmz05ztp/0k5UN2
ORxqbFYlC0qoV85rXpF9uenssnbPp9jkSQvMAxA7LK6tMGV8qZU1QItum9AwxoObsT2UnQ/LTIbc
qZfQwiuzPl5VfpzDIKVgyjhb2q2bQMsdpcoolRJfyvJEhpGhbx194X95jnzwtmZjYScIqe2Qnmmh
PcKS79dtB29bpjjQ9sdUsdUifWZq6jPpCKabki9ES5W4fy821OSj8YKCvhk7mhkFQoco7wIqjjmV
4OL2UvKaw570FSW4cGAt6eH7NeoKdbxeR0wd35laV+i2blpZ+BALMkH8V67kdE0r1LfDZHBRHQm+
zeQHC7+WuT43Rc371he3ihSCc0eDu3p0WzjSuzvOoopF9ycXBFa02/dWaboPwOXyVZ7yVbbgK0nq
VDBuIlDN42vu9yehGzxU8YfRL9oD5EczjPePd2LoXwlqB2T8EY+yxv0lr0KW2vSgGX5VwZp0wERA
XFAcBdnsflNQf0ZrtKXOobSkABNhKSCuRxll/JzlYnzcPdTtyQHA7t3Sbk5CWxvFtFmIjyEVC3r7
pSy8gVvJC3seZWxR9swn1WayECHc9nkAT5c0uMAJzzc++dS0Uoi8SUwUxUONwc79v9ccYxlV9cmV
c4PV6bQOvm3qvUBjPXU1iQbrmVWmiyqKHO33oy/cD8xGP4+azZBp2bynabIN/YNsbnTQWyMMbO66
+xwt57LMR+n1om32kKOQBh2HxCuMqiBYvzznL7j8KMhVYrrCGtdDLJIfcbVJSmKgzXw4e5I4/wvc
IseEBsERW+D8WycudPrb4dVM7VijiitFWvRZ//SdNslQoDzpJDWuUxyOg8RiqLjKxHvlKHBTw1dz
7iW2XeLtIo2m2fkSTr6/V0E1Y5Ylk44AC3sTxRwQyR0xPmxk0JopPTfdX3wrwWNxBj9LQIChosBL
8M+cpWdPhFA0bX4wKGk/2z4EfNNz5ZjWFF+NYmxbsH/AVRt4Up9jbBRvMt6BhWCvS3EG7uOFiX7E
8Y2khSvenCahx1pYd2f9ms6dzVla3lr3M5z7Eyif/Jy+yq6dPeLKsaBQhSgZ/c1nUoj0ngaO0lBx
vot1dEiOGZagOEjtWoG9zGu2xEDgxUO0Ugzi7fV4ILM0/kutpsnBg++MEPDje3RavsFf/6SBB7JF
6hI0wkyxTMrzlKlCgvb1l5grBhSOqGUIiHTfFcff4ELKtJ4TFrtCMypTNc9dOyNmI/ITq4qLEQED
W2JTeScDaCO6ts1wMRdstQIdx/KgDRlGjPWHZID2/3GDsgdS/TJlLvkMw+xJ9YXIBok5gEXjQUWR
mV4lL4uRcGUY9d2bTRC+/sB0+tjtCsnYFDCMa8x0oIHLvsXq+Qgz7qU5/eYtnKx39tqZFdMVCvaW
WVyu57Orn/GwC60uYTj6uloLnEZUCiic+IRS93kcfkTRKx1RSdBXWp7ObNeA/2VHtHilqJdjZnve
Q1xgc5hPqNT0rKy2lu+3HVGXtU+C8BJp5RqVgGjrfDmIneOpSjd1xKBAbpmv1SgqkW8g4ZNjFQ3a
JkkQUfGuGkq9x54q8FgMaUp/etrjsQWn72Vwj+xd4A7zhmq8WNxjO+rLl6AICLcpP3Na+0S7I+NI
ymczUeS6ds2BtSxF4O4+yjfdEtJ7YHk3IujCQknIQzy2IqaiuwWJr6JpXOvG7NClS9D7G6iejHQq
uXbWFA5UiEC4HfAe4/UL8YgNuez0dXNb6bd9UGWKcwRkwAtqbLd/mL4g1aMbBFIzWh/GKn3Viqu4
a3yyH7y9RbVEbCrxAPaqHkb3WOHzLTY2WgtnQD4iEHQRbmMeFh6l/jaFUx9j8OTfUd6n+cBuIUBS
kS70AbBgxCF4ppKZkHgdSPM7YaC3csusZdF+RuPmXvTLzk4TIudY/mbMSEGUccEOrh9DONtGtHjQ
MAVMNcweJVpjwOP9VrNM0CeIMP7LoeA7lT9q09Q626exoT1XZBv03tPxHgvul9RjdIdFc36xPU9Q
8qFqbRWWIfnB9gz4gTmGySFoBJPWuNgXaUbewtk6S688BqkZ/wvXHRKlHxaoklIXv1HRHZx7ky1M
0+++1Uqt2X5uW7PH5ILIKRdqVwGofjUg6m39CxWwXMMKD5o1OqBOO07xxllgMS2bIAChMznAi/+E
Qq4LyaYafl6gejH6VcgH5PUO0tOBOjdcsH4LejrYqmA3BSE3f6dAT0GLttJrAJeEm2sq7xDIXvHw
Hfl9RPmpWDP2+AqJvwfuaqeSF/MBpdJUQRKzm1IiVCEzZHM+4zGg0DNyAE4jJBysZV5EQs8IR/qp
iOIFI6sr6VN6xNRmms5HU8+8O06CREtvPWqNd3ipgujIovapl26A4aKGMJWO+XjpK8Fu3sFB8y9f
7qmZCYJpnMRJ9rTclOrC/6aObStXzpW7JC9cEu11pG/8LwbvwtmJLuQpiuQmvMsfieR5TGh995X/
uvfiMFzBnefwelmp6FzZwbXJYaDqf/PKpQd0U5lOooU1jW8LVkzSX6jXJQzLyTe5fOsUe6odObRd
zdiUugFGlXsKa9fu5uoJqD3ocA+3rdnh2kSCyEj7Xjv8Y2VNBj/35BHEYNAidnEQj19jn5JU0tHx
f3sSqrPZJx4tELfpl+NeUXUT34+5MRhCE4QnNDd08V/vo0L/3yx1nLQ9Y7oY//UJedHD82r5Lx95
e6LuBniIdtSohRp1GKhHiA/KPZduKluvU5FprHUBcmEEd0OmtyNbbDuJeeinKrbFostLR92s92pW
0+3SsuAZSKO5HX6sJG+98KP7tO1S18vB0/pQqPxJGwEPlazgUKepqDOxQtYFQUDaPGf8PGuag1sD
hQIwxS3hnbYJ1YkmxIoPXHbRfnAYwaTEqdNSlbVoRkWT/+jypPdqYVq7vTnsESrBRrm4S2GJokrw
TEjCsdoBg7OfOD8VdVxLHl8g1fCZxIl6lThtXW1fS/GTbRAzC0MuZgG9/68lTPwxJdOYpiNZo7VL
+tLocGeFPYMOlxvrB2S6NJvEXKZy+G/Vw3WM5X+HXPnv4Lks9m+B34c07w76UxG9koIA4HSSQn4v
rLvJvrYY1jB9rNJHbwhupwR39d05D/jgrccI4W096Xfz9iBiA+bTpWgOOjUo6/VnnT7RG7GD6JSR
AUbQyE6ijpugbLUAjedhLYt6Rljb+0LczAdUMLrKyNwuI1LxswpTViss1PHcv5sZMs59UBmrqMUX
kx/7viXmV63zpShqRi3V93IZC1q6RuC1YWUvuHpw5oKN0w6UYAdWz+ZvSLIAm2Ga6Q1tVjCopJIE
uRSTV0XK9EzQKV6wjQcsEXry+GZs4nhN/HtDQwlCC+uqAVJB3+Wyso7xuH1mLAz8iIXUZ/L7aE+j
gx08aDzXHa/qah3zuAF6hhnXfoeF+9gR7+oeOp02vF3LpVrGaKN4IIQLZGycoDTmhZL5eUWUUkSr
X2oMJvbrRawF0pmSJuiwR+QPuIEwUiDxdeKiixOzVU/3sV62uZNiYPzMr/w8gkmKolpkgcMqoY+T
1D6HNKgNl0vCG8KH6Euq0eAx8bWU55XencxVQRYKuOanPsBwer4IK8Sx9GqzH1IrD3CeEcOIK/4y
9iA4lqyiQBxhN6g4UqngPulYItoFodtniRu3py3djBr2FG35e2/CJGC7+gVbPKh+e8bkkBy4dlMi
8z4KzD4dLFzQjL0PYLOPbOvIxW51usXQ5jrn/FFneU9oIpArn/jS+BLd/3yb/WJpcH0qxt0p/9WQ
1TY0fnLU/Gt5Y7eFvqtKZgNRP9R8iXVP8XRYOhB1YhIa0txxFUM0Q/32eSehQU/dqriiMQxfDMpH
B44Bj0sarvJxsTz1Xg0v7+VcRYQQAGp0rbJ+N3w0ziXw8ElOQHOPSTyaV2AJVGPot6xS1e4E3Q+a
M2EdIeRMT+DB3bPUjdU/Fl5mHIPZIjlRaK6LBxCChpPbh2fqJLKlgnNZOh1n6OHre6tZSaeFCwGe
LIf7oESKWe+qBMnd2LOs69vQ3T3Qb/vgT4KBh2StgBDaJP8Ns9ZkCroHO2h9qM8+F6MTMpiLwL30
3MNlntrylo/eJ/630jWJnMy+4QEBTSrsfdigP0njyD8DDeyrCnJ5KptFhhllnQTk+fM6Y6OeJqZq
arXlnUsZApaogBYcsw5pVU/H+/xke/eqMrnyETGffIgt7iU6pAGsngW3JbK/rtF1aJ+p7iqXuoRF
OyZsLX9mkKaOHrIphGWAAi+SGgAsuPAKjrggnIW99/VZQ2BZGfj7xI3YABYuLePCygXpuhE6suTr
jMCbL74KF3ZToD7C3QOhOzWF/ZircHtw2dY8cqxGACpA56/gOPDEX3S+Jd+nProIZvjChYSBjN5D
CNjSPs+66pcmvt5HVAj8FnEmPpkWA73pBu02OUxlTEBjw9+toeIeoqqLA494OgIZ79Y1wIbMYVkY
+mG8TUzA8UJT1z/iPIeqWNKkKMVpt4fxbN9Vs+A6hEso3mGBTzTKE55fG8PxuNSpdExZuN4O/Irb
e0xTwy5u0AdC1yMYrDsmAVtlANGduKQ7vqGGlxU61Q7JrnmqrU3iRoLIZ3Q0x8mARZP9ik5N5PJT
pzMp6Xyr0vgshZQ5uC14aUfDqJbUyzktsd2o+GZjnHYdzC2TDDLtIuF4UKllqo2DXkhmzcpgAHp/
kcuwA7V4U16h/h3jDJD8alGFponplPh2sbkgUaK7LTS1zAxdBwl2mvneBs+nh95WC2wOlisQR7Ud
oVIQXiBkFiZG8ITqRMfs8ixeUE5rJjznzsLEaDUQqmSvSZnXsFJKUL7JtsNtREaIiZp4nX4fCY9P
rddCShtWy5/Ontp7f+rQQUbEvEcrd5FgZTyhBID6Ch+2+dRG4pKCGngdL6F8SF2WsAnAKxhr+f22
/zv5HbLp34/TYTr3LDYba379CBHkiRq6WGZk9RPM9Re4hBItD6N/9wPyORAmEiToAlIiHSWUPCjp
gCqLID9lC6eQm1EKTUrYJ9p71sZBRsnnIQmg/8cISDQR69sPzZlpeFP/TAxBi4VP4ILe7ohKgq3x
ZzK9rp2y6+slHVil860Mrj/IWmH1SDi0iVg77M9JkAODWzmlh+BPspxq+pd1e8Rctq+K/tLBndxv
yDiu8wU1m44P+jXqaFA8csbkW39B6csymYS9mEjlAgyvZYOw55bUsowuA1hOKp5HS1vHzxAdsGnD
RBSfk1/tjg4yLz3Upzy/iPHfS+6BHhcJY0yZ57ThLbEBIm0AlG3KaGsQwN37uZDaJQkv/gDDybeZ
IiVkcgDLGjKxhDf6sid4YA5Pc3bwdJqlHkN5lY6jHaNK9Nkk2GnpVjMCriqs1kVcY55u5Ou3rsqf
kS/0i8eEz74jpBws6Dyy3NuUfACmrYSaBudqFXqYVDEQaWVcB6cP++/Her+waDqFEG/oHL8tc/Up
Pn4pWWv4o1XUTVidmxouj0g4rF/ErOCXHJNZK1hHZOpFk6XC0JAaQJ3pHtLfQ5z51T+BcrP50TnM
WrufvHIHD1wC+y9/CZR+MchP5x2LLTndiAZZwI0ub38Lgum2xRxAgvua/Yqr7dpIyXT/CQ+eHpfE
fxiukYJ0HK6Vbhts0WmyKLluvDKT6ZWG5Bn3q/qdglR2rj1utwwCrn5gSVbekDjQ2smXMGmfPe3+
qOrpAdv/fFWhEGwLOj1C5uc51IaDF6QaoMnHbeW3ZPbwDvYH9QvOleXjEwG4idTE9ZSd3gDVZuSu
8cw0ZH+X/FLi4GdYdqTsw2YvIkR+cE+hR1xOq/LC0zmH+vk1RV/bxJ5jhPja4WNhwh4RUuYvD0iA
A5d2DP8w7qH+wTS2ccaQRPKNPkC9ugTsJuu9JvAqtyw/YhiOF2mgiV0uks3zoSBErSHuF0YTO/+4
YCZ4gpxU/n1WyE8Yx5FAUvYF5tr20dUlXRJsqkHqtzRosqgLL3bvzqUvV3lkqCeTYu4DNeruXjgk
EU+OjH15ZK0Gwkne9NurdQ0pJPN0uMO71YZb22Y0JhaVbiyl+tqz9N0PDcNQHEDrr4bxF/n1yXRC
gmQlL+k2nC/89FsojXSrtY/SjYWEwkDEck7swTpR6iKSkktmeGeTRrQXxOFMGAhp2uW9k74Jj9zx
dp2ZbN3uONGENcDwTlzVZN49Tj8DAAHunA2rvITm/4CDsIf1fzo2QwvRuhvCbcNtC+RnV43tsPMy
cKQymEk3MkTvS1Cb/11+yDVvBJm3xVuBpsyqsfKbb4AfkfSmXCMKwIWZdo2e/pHyqNlRKKDpc9l3
zWckWBye6wDAGZUwgV3Iio49NG2+LQsXbbBU8t+cGRoF0BzpCtP3tpxv/yDc1lQOY+MicpKMX2Ds
uBFNuIySH7+pb3DNaJwnqbloNuYCBCWTa7QHP85eRHrTgt+jzhF3oZ7/3c+GZQ2fzCX4ISRTJgP6
BzwyamXjGTh9eWo9NeQWvQXaBn5weAWSBmpGfaomqGem1bF+iYq+OclVw5fZPJawkj1u1Uuyyp7j
bCO+23UIOR5d9tu1ow1L/uMdDCPDkGqYYUrVGLuw0ddjIH2EUR/SJRaA21ru8VGhibfViz8z1GnL
qmPdgZbUW5nwUkgRwFKG/Lf6g3YGJw42XyZuZWoQXrxNUXTG2/BWjYbTg7uLCtTVEMXq+x15EuZx
MqduSEAkd8yD7WSvckVf5JgzyCrSAJ2j6JDSOnzWssmA0isECdYRsMyjwus7V2fWpEmBBDguKly2
BTc9CEoewRMip8V/7K7+XF17XrXLdMs48Cb9JDBMUWWmHwueVFzRbpPO9VRpK3+gJTl0/EsrPqSJ
hMDbpJ8lI+/GT0GrKk8DsVHBQu4abdNaGzOugubYupXWUHvkOGd78ctmi6TZbsN3b8dvST1IXXgj
8ujA1REUSyHhLj+a/H5/67/inc2ZpOV+diTuBMy6J9w9lvtkNQJs6XSSnxCEKH/TVN/6VDLS1sf3
qane0yfXW42BVJeTKYHYSwd7MtHf3+QH1nABH06fO36OcombYurSr1IllMXCrDU6ZFcEoJWcdd5o
9+4B7auB2B/kb5QP3UPnfzBMcEHnd+Cveu2gsFI3wboPGOoSpwy1Sepp1KSO9sFRkRAZ8XmqLc1y
4CYcJDzaudEf6zHshgEGjeHT6pVxd+IrRWQ5ykq0DPflypTB0kYqm4QrtTj+IDPpJfR8qKoiCwAw
L5RRdUBw3/PP1ucFpriE83AfXJPuZCKnGtYeiOc2Gd0UCUQwGEKnZkvWzvre7Ic6XdJ90gjcoUsx
peJ+NvW1HnabZ3rfI+634AmjATHDe+AmtAs6l9CwoKhkCYFtol4Z/YF1/EUPuJVjeKLLXRjRO51s
h+GU73EvKPFg+XtQllx90g3hvDWTBD+sBuz0UgJFC5f2ii5jUtvOwuRfaIXg+ImqLqklYWmskBa7
X6gkbfK9omHeJefV2myMjCi6nGQViBQp71NI4mUVN9NsxlSra63Q9vgNRDf/9f3WikXTyjT+l0dS
9Pi9oWKRaag+7fUfA3OK1DDIF7yhnMEEYxJxSnDNfMVWux5WeBjVQplcVUDU8wBRxyi58j5/MJwu
lZROE7J4F60x4W26V/2m6vCKL9lLEAYS+PXGwDnx+Hd0myuoA3cZGgCQdE/LAfP6Ac5QHEm0hQhu
GE9LadHGPXum3HF7B8Yu+xGqEwnmtIDROo5FO6kEq9SWsqbLntTg5JdTi3VQgXstcwa4rhf1aJKW
0mWkLS6Fvw3V3wzASq6O9bH6N+70TdhwJzsxxUnpLxLbb1m/yvmMuD4Mfvv/8neLbjvckR2O49cY
Sv2uL36KySsidPzAdGdw4ePQrGspP1Fg0EB0v3jNivS0uLUEKjCeysKRyWlMn3SrsCGuR8CoxiQ7
JZ+urI/04a7VFtv9fcGSMz45x2xGqEQANw0DlPz6LkoliA/YIIUOYznxUO7nk65OX0ehVfSM1cLe
QO1mIqRkham8d0JEIhieip8KdNgJrRff5OaNJVpVjg+UxbPLUS85z+NYDEdy7myIuA7m/0JS/Jo1
2fo/GShHeyQvQrs/sYBKU+OxFpOlyoozKlu8ID6GTfZ9r3kpzsTEgyz11f5+NHYSwH8uphUNUCxi
HJuHHfvG4o91oftyH9WrVkdu8dezyFUCzKBJUOcmBodEZFI95LPDC847pIMXow7yzVfIjjorceMb
umEXt5jUf6d+o6TxbvSZ2DLIe/dYXeistX8Gf4i+c2SI4L0z5bkaxBnGmo4Y4MYiCdeEsn1k7qXy
etLIeljzUS+xH0pNLIRkPVcUK3rgBlQ49tc0OHngrCi/hn+TYnfH9mOYLlOvlyWmnXTIlwNPrrOk
zydcmB8dOnAs33MQVjZ3miHZQcRlVsXDd9z/rbfBCuSk7pEikIo0pRgzzVFpGVSZxxablua4XQeO
OrRRyn2OkOyauNhJDEeXpQR4qLFRK9HoOh6KbGFwLFrOMjsshWLfXAJpugcvLYEngchwTMbGN7v+
5x1K/nAYQh8tcMc2VYA0Syf28abwZGo1VKnJ1SniuxB4JyeZVOeBkqq5AymZ58GcXnc9zXOUFqFe
O03Oec4tkok3oh3PlAQesnmE/4jvLd3tt50tK86RJgFCur8HaHFhrvJHy18vj2fbigsf/oBDY+Cq
jBy3R6flDJi4ukdrUJekDEZI/14kLSz6isaPI5vi5ksHHD3peqM59S/m9IKe5UOMA9iGoo+PFIyt
r507HvLoQgRb1dCvlRZagS+DbzMl3tUrMe6RYycJA40NZXoXbsJzq5+GnuCqKgDoNkn0/3vg1E7V
rMZdb4Bh9N2vYOz6EmIfPA55pETtrz0KRpoDpOE0khNVMH/p8AC+aUh4ZbulhUxJ+aGD9Eg1qVo5
9OFtySVVISJZ1LE0sG726Fz/Cn6tT/kipp0y22ebmntOKBtMn9OdLEiMEBYpppQfWeOcagS86kJm
SAhmC+sJi2cuVVt5wIfkzHVtipF+eP9w0Acdb6yid6qzheB8G4EdQy1r5hK+UjicDmhvGyEJY7Ng
wBY+XApk3Y9Jdfpxbik57MdNDbk9A1CLBjjdyOmLIUfUw9o6k0iy+b+MlPLviScx3d78vH/peuFf
oImxeKSZwqb0TcLbEghhSliqmfRq2N2ZQmtdJVZWGvpkW/9s50kwRsLqacALXPS1VqqcaSCoSz4O
Zj0BOVdllNlDAzSX6SvtyJv8FidFsIUeOg3EKw7ewyrSzVTk0jOsVfYdG1oisS8MWC0tlv8/kxgi
w9L6W1V21bNVromVzUQ6sSUeKc7KjrrbI9YRK4a1rFDGDE5SQN3MzJgkW7/vykbnFe6AFhohbrIp
v5PSSUwRwMFDGHzki4D2X09Ilpv4qEckor6wnGfLBrrKJ7PO4eUoKJ6gfs4GBoczny6xQ4/El12r
6VVSHpu6av5rfbDwEIE8QJqHgwSKQFK/f+4YLt94mGq/EWeXw62WGVdgZGppEsD0hApxd3zkG6oY
ImPQa7MVLaIPVfjK7DxuwwACaGcSgmnOHQrXrcB+lpBcgnpQU9o4cnBgdEj3Ru6tK7iTXTZ60tcL
vAChMY8hIg3RniCwH08AwTtwFEHZii4V3BNG0ScgTxIvv0d8Z4GbE9oBnNL/fCxs3jgkvEgRTtmV
m6oGgFsyS5Cp6PA0LCRvweMC68FpIVsToeJq4cJwXv50JxoqcjonBUgkpNPRiFfQrqz60MaNqopR
9hIeFpEryUQXrCRO1yzm8CBt8+VCbGE5idSuPMMGE2uxZtchYs/WvctMTwpgv7V9ybiNrne5OCZb
5n0qAOAQV9xUs1pQY04yTfIff1IX1jOt2Ix2AKQEYQYsADLqUzAt00+OCMTmMTEViCU5W2Hcwtk+
9nZhdnryhtfI3Dsfrrjox89nMaz8FQsBfoGaUCMqZQqcK+q+1vxfsk2IlTYuelnXU8xwBV1riCR5
NJWq2Q2CJ046BWd0l85LRGBGDrhVrzuF2kDVjgABXLTwJbiFfwIVxffOzXU4wZepkC9rE/4tSMtJ
mYjAzeJ+5a7/3+geseY0ie8hg1WR14RcgbgGOaGddJcGBRlWLA11NanBZ8zfLdYPWX0NIbVhk8hG
WouCQeqrQo/38sHrZrCxicWt14y7uS1AncRn/pw7QtcrpPCrPGTzf8FjoUwqUVUgDlZNQNuc5pbp
GvbdrGT+7BnhJxNfXdgSkhiUWLnMOX6fstdcSwN3vRnW8daSeH+46/O/N4u+5nQF2CTOwWKGVfA0
IvBTiXDAzAmD9rtUikLz9jwlmBC52sQ+07NVAJbKzpl0M0S6dqkvxuPYpLxmyHoeSd910dKnllqS
0YyCQCp161OfBZCkrJwSXwQeL65gvXt0c3ItC+pyZ2QdpFPs73eNicb6jtshZrpw6eiFyPYBRVgj
mH2lQeW/GYTZXQELMjOZerhbUKJuxr6Y876bFEeW4jnwkryA3hkKy+k0nOESAr85qBIuFrd80DiV
U/hOFh6vsFMY89zbNunPPd2faGiVrImHca2MkJE37u3yjZlWKYA9dcNVXRNOa8kdaLDAJfV448wA
gJDQGgFW9tRnlkLUvKwW3p9wWLf/4mH1HTTfJFa2r3XHConfgUlfsD4nWzPL7ewG6G9tJvX39hCE
8S2AJh/pTNsx/vGJkqeFhnUmnGL/ME/MfxgrtyasKI3Z0BBqx9KxgAfX/hmlvdVmy8mw5rwagEW7
HGJ8tEVppmAuhTUrKqdUh3NLxnTSO2MuQA/2eDUeZsn7YXvCL+OKYJyCbYZlMFT+rJmyd5pbVzaC
mesj8HG0bgDVXKyVgnpLjhDiEOZ69X39I4jyLrnQO6BddMz1AOhTEqnS7aqk4JUyke2TgzaImSbQ
5/gl3//TFROlvsVQImpa9S1gaek/xFsistQja6aMggvPKTsPkJY8Jcq+qp5h6EeswHwyxLYeoPMF
LbUPkMMl0/7iTXSz0YCThVK2voX1fRoViv2kfTVcMTHKLlrKneUu3lmkm0lT6sr8mWvhqNRgH5B6
LXBctK7hpoVFJp1fctgoOGBxyMSXw1deOOa80S9HHwDPOLhNcYKU5ThRbh+Ji/mBJpnJCFGf8Qg5
U98ltHkbKUrlLxk+zH/jL4EFLWPOtNE7dBzO2LCmMsui5YBJWl48HUXBihXRL+k6SYY0+7ze2w+P
aaAdrGi+BCc1kMPwm6F3buUQnYVsHejASqlqwQG19ah3ld6+0RUwMEAgES45ctZpG5wMvutf/xzy
JJaXBfpJ5+GR+MdMMljPjFXt4rWtd+CsGKL/r5B7skP9Tcx5OmpWrHU/48rkQckRzqAfOUtmk60o
OBFb/SWW/cHy+6LP4/RMhtuCn0jji4EFBtUTWzurKlOee7jCAYK5DaEzxnNxhqrfNd4HAtPF3+Zk
sHrWCEyjnNmhyQrwb7/wj2B49yRnkrJKvlyMZ6yy3c9Y3z1H27N5cLTBvyEaVfa3aQemJFk7id6K
gdlNXwHX/x0r+LB237c5T6xsL/BOYOigTFHo/VT+w7rHFSwPL277TsGhseoPqI3LdkZCXIPqErja
JhV1mLHVDDDvHHAPJCFEmYH4IdfNPYzEf1vfxbASmVywSJlgiZ8urfLN/dpQtRI+RYPr7ninfa8z
Cj6N2yBdZ5vumxC1gvz13z3bCQOLGKT7qvuIsBboxH8R9ZjAtBiI65HA/B1vYthh9gxkrpwJebUa
n/GYG7r6/N5wPB5p5fTCRQX/gqajJhRJL1Tk3l3NjDy28tSgTEAXtizHiD4BL9WSiDKbfsohnWok
xPi002Vs9aeyYu0J9U69D/HCpIdmALdAl5/bji5ZulNA54nL/B6SLKP8ef3klZaTFlq04bopIzob
Fy6Mwj2JlsZUJuIwd4Ldfw62BNtIbM5AL/N7ewhmT1Qy3S9YweauTl52f56p3OeNmpKGe8ujj9bl
TafrZMjzTrdAqleEsYjR+8f3ylOdadQkcLiLFUvmoLaVKiRdctzuXiX9WDbuNSoW/rmrNMdYDUoF
GdF8nB7HTOQPJv2I3fbNf2eK+vcnAYOhMtOD24YnlF7ARV9fD/XEJtEzT2zf/5rb7tHKuOrkYz12
/1hh+Gs5rKbmPqQxvmRmWjwRB/gQdDQL3h+PhKDG2sIjzZhEo4uytw2gtMgWI3/AAR1rk/PbrpjP
fZjb8CMDpCGfHWH4QDxb3ZJuGsEQ4qcBGv5NMMKQGajZZ0Ah1VmAEe009roKFWeucSu9ToCUooTK
dLxFIQZqbqtBXWsSV7+KntvxvAkq3GHwCnypn6/XhW3Sc0MJvhmxxQ+z3rohCxH35WGufSQUiR53
ts8OTAD4PxxPswJ8iQyY0JrLL/tQKmNwtEe04QDZi58QHBcB2uYg5a7ld+SeaXJSM0luMXDtCUp/
oCA1wa+iDabG9PXgmZT0g+ffx1b7IJZQKXeUG0OfPf52URsZAQuTwLZ9VbHyyZAoXstXspbzKnYo
y4+np/kLOEnnqRvC4XLj753EXH86erwrIQHqf4N5vQLeu42tWoAa6kFVdBV2BpX8iRPz9mWujJBo
fDvj5pskvHgEBUWWEaFVI6ixInzeEKkxv7MfRTHN1sjyNMajwM+eayyfFv9tblPfyxHlvArneuNE
7sKijCLo0wtyZeCS7+AnMSGcoM7jOR6N2HgNHVf34ghnRHCZECjrhL6eTPlCzfgKIq6QP1d7eZuo
B9vGmJlW1kwCHoDrc3j2INPLfegzpO0d+OkUKYTL/aLFnddeHzQIOZNOLunpdgOwZmQwQuiLs3ox
4Y+pN8MJpS+ZU6fdL/ZKwsPETUakkSK77G/0bjQZzSORAVZmYyjUjGnH70h/E9VXRTyN7Q4eWXLk
u4LQx8No0cbZR163nsTSPQitWbAHI8pghRxENXFsbnka0GDOnzmYeqGyrrArvXrZGQL/RNPblM7v
XwqXEn8Oib7lnlwkS2REYRpi3mFw/PI6ja2D6hhVZLKICxmW6H1Ulc0r5HEekscexrJ6k/6GZcwa
Byikc1eilat8docCh6szwimLOLJVkT8VCXbEdW2diOc7Qtv6i0Kr8TnDAlFDG/x0EGNHtYYI3JUG
YmsKbYhMWT9RqTVHIRIQOyovgiIIvZLvdYVibpfdt6Yhuy8DF6sdLk/XkEltvwH7QDpNlCl8OOXg
w6rt162Mo2evHKX5sKDASE2UwMGbMmriTTWudNmuI0GI9DiHXw0p4FXazAlI3arRom/77vkzi56z
71qfamEGOFNny7pAnQnaS8BXYHmWniLdR4SNK7ofx77RwV0fMAkp2kp8P3F18QhInLFgYu57ZX/F
q+d6LK2L6F1FPckL2L8MnQ4cAPlRtFqmlI6eKAYxmfD8KaUn47bB6Co6uDj5W3/8jy21SaHpHHEy
682Y0gHgHrdGox4IEu67Kba6UNNRCcDPadIdxb4klE4NyuhzlQPXA/31voLnFH6c9I1Qht9sFVv4
3S394OJeVh7X3UjpqRRr2HIxuqhYMvAtOt1zdZKRTBqwss1F6ozRbNOdno6yd2lNtXDw6eVhRVPC
KdVL2L6LHKjibvAi9lK9iF73XPXjOK0Ee1dd0ESukaQjOSL5R6zJkFPmyrxSPd/AReQa2bzxev9d
Odh+JPHBbrI6N7FBc0XA9I7NMzs1pzhDUirUZLFpGSRzaEPfOa828PUbXpBPamYTCHTIezGYRkru
4kPSNpHbW8wpSzT256e7VP7LmIlpNce7zwoN7JFlFdCjSNA9jVuQWgEIA1rjvJXzTSlK7r8xF7Vy
a69Eky2AgarlzXHnemHV+Z5Q8L5nlidFGEiD/d7bfY0sUgjlRT/CvEeIP7XSjzah2vCEu65r7XyD
WZpbAg2o8aVV9/L6BBWehXwJnGyvtZdfzUS2O610JyAfI7mLgVQHEodA6hrEmJTBO9Z+sqZ1Kwqa
HjAqqcSNtqkQLCXGUauZe+UzUENHM2gY3b3XmHdoPIe8DqKSoWa1mNnypJJGQsXQo3TkbQFDeDsc
gOJb3l2fZu5o7/OBGC2kUo23Vve7wTaVgw3luOE++7Jn/yhNQRrns2wHvMjisw8pDB7OVx3EOWbJ
4jsGEadMxSVODV0S64rbBRrSpzEdLVQXrQGxJlt+NHgDkMxUAh9ICMVrQDSVe4/yjyA6Dv3kVinc
BGUtiNVj1uQlf/KbNTb7BgekeWWfSvXesO6BAggllIP7YSeefM7vWHd4ytZX/2WBzayGXQqJYZb0
bX48OOVGfwDFlzZ2/w2DboR40h3Ry93rhoMx93qenURe8yd7rM+0vUJle/wM0ke4kk3t19zAj7LG
lTZqOj7oWcinpQJH7aaQX+wcKLG6NCnEXAHGYuXeza2qr/IO0XSQYLa08wOMcI7a/OQ6kMYAK4ao
XpYz2GrB7hoMfGXY3w8YdOdB9UZxwL/ib7X6WWx+8PS/dqcixOo3D8rES0uZ5Jg9I6BpVJo31n3k
C4L68szU3UptgeXC/cXuQkuNI96tQBNce9HPxkR30up4AWZb50a3Q9om4J+HhnYlQdfKW9E/rXgQ
IxGE9vFmOeQvqxQY/J4xuHyF24wuOEJr+1oScxkqAZvC7Qr9StLO3stmbZ+z/Zg7dH/Vug+ujVZX
yzcz0MV9vh12UmVweqTTLmheSlaLUEiyCj2Y0ntUdonEtTDMV2Z+IExz8td57CQEbrHkvcCo62e4
KMdxPwE9wh8N4RhHMdAxpbx1NJnHqnrUYjCC5zLjOGNtgc2dfjAM0mWYXD8Z6pH+GSw2Mz6M+C5T
GGNMMCUWKXv29zn8m1ya+jiXFO2MkMuPlaRSLuxFl+d+1drBTj3x9mN0wywsCh+5jGaLdSSFGXPD
xGZCYbrOo+wDBVcOBSgKKORrcfZ+7P8lJi0g2jnvAhFuXvsk1vdRzKctrdz52hZNTUEkNx7GWKh6
8mYnfKcf/VtEn9f0BNGir3bhUjBaGM8rP1CHD0pRCmfX6sBNLdNUtPi95csZ/OmgBN4+VfVTZTjH
7l8VtYBrDRNDu2AyQdHLO49wEFCG3B1vu9Tg9iwMH1f8J9A+i0vcf4A0iuRZ9fPses2kG+Cxhctq
aX2oLcvUgSEWjJ/zdeZVbAQDo1LAMej6dOTEeWaZEkRz25jrf4URLY4hSu1lKW9b5kumXXRGCK8n
9aWS7Fop3FncsyMQ8LkRZP02oWX7AzRHxH7XwDh0hqQisbJo/B8lqSqme2BZePvCVfhnvVryUyYG
ll0vmS5IjIFRxHeZYRVGYvI3ejuJfYjtiKDAr72e1Xoqc9s0PFcAeltvfKsssi+NAUdq5icSaDxQ
uIV14c7MAxkgBfRNxgpH0gQEhUZK56qVd70rZarnRgPlHeRZlKH3Xv2RnRibOng95io7ivXefeyC
9tnvl1ZoQAYiyljyFIGeOVak9oxLLKPc9LcMNKJOOKm2NENToFz6vkttJ1jFMUj33tQKUCVTWXZN
O8CcBdGuHjl3BEslxYyBsnP8mpglS6So5LVbEON6TsD0/5Ss7aZVkbEovhaHXBM9RUhWtKW5SuBu
FJrtmy/AFr4taI5Ein+jgRBl63qRj1eN13CqdCwN1+yuku4oLpUzTNdNS2iCIZZSJWfvYpF9SqUd
HcOYMCEUC981crKKapE5enUnQA8W58oBgFqr1H0H2cJLiMTBHgPwcM7Kt6BPkoQ2sJWNYq6/soLE
BpLklkUsIjdC2aThg0M8Xnz9GsaVDPYHImjQrJ7giNcKVOKUNCaGbRYyiMCSGUCkipQ3xW6C3iin
n77a3QF4iSAaS4MM/E0rKUBECxbKX1U96ErWtFPd/9vu7Szh+VXOocPU0Z9/k7FtmjpsK0OKlfGk
6ukZaLJqDoTrs8amq8J0n/vmr6fcjAnG/nEItrqm2w4zSJDgRKy/2xWQTY/Dg3gPoq2rZRHU0c6z
j8/n+xtLYUZSjbDJiXlZGnrN26P9JAX6rCPPjmPktI0QFqH1ojTgO8V4EZE1tVaPn+kLSyBhFJU/
CbCq4zIpEYKymnI9mNd/bkbgkCo8dYRob+/71ZxxEHB+MXMrfiWRp9VvRierjCi+fT4AoGDhXn2m
o76FeJPVVOWKOOiaSEL+FgqT9+LzBNqqyLEaBB/tmxZpOa94WLMOJ4tANsIdUZU+aiFAoBd/i4uu
CG81YYbNR1gpEUa9Skl8DaNQTUjITyNYG6bGu+aGsUON2wt4C5lAA1RVWulOHgmNDJsVqIOkEVdQ
nmeS8LPAHglG1CU01h0Cr3CmZfU18lSgvNdVro3dvI8+jPIfZlWtpdw2AQgNgjiZS1anqc3CgPY/
Gfpcb/UDcywhEFCfsk6uSr+gl9w2UVWooleogloOZreRa7ol6HeOFBnO2enRkecLenoICoSaGTkG
HM0fBv7H3uA/e+ijRwXGeGpsNZGiAJkiBHfXRECsC3G51ibEoZGMkkWClkLK7Eu48v1ExmHWe2bW
gVTZ+DIZxbbCsXYnR86bZ1mYCdZMe/0EpPTqSJFDsA+QBVFYHznQ/LfrPI67DMU9yNPqEqAL4pGU
mG8YAh5OLl+TAPjtVbQKThaJoXzihrpWUl2qNZT1SsN+Va4DenELX65jU1bGOIe8O84Nf7B+ooYx
LsIuVfKHpQ//v+Vs26tuVtya1nBsYajLhLpCS13CRrAP1Y1538RMRHYsyNe7G17L3quyFcDkHy9G
oewp6XEpveY9yV/608Ur9nSxGIkq5bNhYYKbXDah+4b2qyLJGWtrGcNHYFHcP6eyhrbbJf2y3vJH
YfIstEW7e3S2/2DWTi8kt87TIxFhdoAH3q2bfnwYrFrxxMbc12Q6niL5beiUpqKU1TRObK/38qI/
caOXR89Kiz1mOPK5ciQTYbU9KcX5+bJgbNyU5gsZp97NitiaWHHPnFflsLM4cU52AsHwK6DNV/gk
vd9L7VfXBuoiaJ00eXD+5OZ+KLPBQiuNGTnCkaxwu758AaGiJVoaOb2mQY1HOebJnsK6mjS4vR/j
4z5f3tzvduAXf4zUmuJf4MBhI+DeL/dKWCA/ozEj9lNyy0glk2sfNNHO7bpm7huRpyRn+PTuBMQj
TuNbXYiuvmiHLVJcqp13aNfa8ojjN3n6v0EiIUk0i9na1g5Ybu6pDl1VT8/6IEa1hOnXdz3VGTAC
4wh4xK3X8EKUR5Lixb4ehM3NYSjlaOv9fuKFrumS5qnmt+3esilziDCnOfIQCleL9P8A2tcMhdmu
q7OxGOBltCLU99UOBtwbeXmAiKQTpcmkemORxHSUJK40AgdCXI6qgOo7MGcT+pHPiHahXwnMvV3F
GxK+tRxFq8DDS8EbnElGpdtK1nenSWBturNcqX6q7/ohDP19vd7Q7FOcNRy2R86ADZihWyNrSx8x
w/BHYmV2mK0CyjBLhmeJcXZ9Xzy5e1wxlN1ieLQokD4qI/NOlYmuy8gRk2Kj/nz6IEDz3N2LWwbI
r0IbaUkdx8cqEF8YhHGgJVbcX4aQy5CRYWnSuagk1NQlwPcOwLCrpouZx3hkriByCp7CB1uBxibg
7kSEIyaN5vBDuW9yJEGgMnMn7um3uSyG8RytYNTlHN53MlOf4/Rm62a/dDHdXBRHoy6jU4t3U9LW
OVV4Tw6kZJxzrupGoJWlcRiS8O8oxF/EImwB/3Moi+Ezi5uGjsqxU0t1bKtlSf9UKomNUmkBLOPT
Pi/8SFTu6tXrNM30jvARjifoyAPEw9sfa9Jx57m/SG1qyp2gwOBFRiDGCHDbzFC0rcp2IVrrGE/v
Zj+8orW4t+l2fdC4QI2MQdjed4BhuOCBUaM3kgrDuab1KzCWBtNhdxjoJVH/4mtOAYb+KK+gOrKs
Gs9+hAX9Eo/5BuBEPjwalqXasfmR0lc3Ym+UGBQXKMvs6h9aADgD1xbXvcal6nwhRHQ3kby23lzR
wBzUABcd5cu8j98xcIFk/hZtjwEOKsGPCGq+7emzVBmU0cH+ZTUPtjFoNqyczTa6Tt0ZktEaRxCO
U4S6dfgM7cwbNL80Uute/CnDORzYInV4Tczis9jIJHh4tMjs/qJxFNLvNMFzG5BLFSb1pK7kJXQj
V+AvdWIAv5QILERg44AYV8H0fb47Pl5f5NI/S3Q7uzPpv2Xoxa1JfIdMOMSKwOWwOlkKB5sGr1X+
nT+y6ckFVDN98n8uVCGWGPVQWhyfgZneZa1R+1UFkPLg/ecxb3atmPPEst9uBvvXIu6kFxDUMzbo
DSQJfgVS6/ZsGM7OyAh+boFZu8b/7L0MsI3lj3+E9RANo64rmOAVCEk00F3ZWVxIhbugpT02uIU3
Ypu/9sP8YZULLiRrqbIntmABySx11uIiCgOX4/FRioloZvcYbHLprDJDJfjrXdnLwAuLZ3cLv/mt
fjEo6kD5jNEAwX5hiwSfvMDUOQFGsGtf/mU7G+xfJGDcIetVy8z8oXY4EEEmZy8vkp1zw2uXDLPg
YGoD+yVXumDk3kvwyNWxxKmFQZ5EXGL1otedBNHziiLOjFXT6NJcZjvfpHq+0sCAk33TcA2wXuUb
oGbMdpaEzodiQzDgK4VcwBJZIkCt3dZiHOIpW//fFXH2Hm8i1/Pl1f2NNqkMZJIC+BP9skH3y17N
k2SoWhLdn5D3armIP1kb9VCjI3YZtEGSuh+RDFRl11GGzxw/39c4Q6Pjsj96HUDxb30kOKO5Gj3n
wi98uK9QprDHMh3vwUnYxiTfSoEBk5sbZM2Nlp+4c39EscKdiUYgcZdw+nsL/Pe8Bq31pzFc09sR
N8Uc7eUxgg83GeP0JL6zS6NgjB38+KjTD+fIt3fcmlkwJybT5U+I+F+cjQsLH/+d+JPVMiMb+MLG
6TNf0jDIFQ7B8e8l5Gir+bUXZDTOQsEwNCoqdBVQuGBv13GrjEThgn7KSV2GQdcWNDVNrEDQURx/
Nk4reDk+jA6owzQagWCUlIBw1jrFveF3AVuWnarYpLHE1NYbn0sMMQS1drB1slxPs0E01ktaWhMy
W8u4IRQbtazakJAN858Zd3QRG3+81pS6NerItAKqaoZfJUMz8VOZ+9KV9ZcJerPUERBVV+BANWGr
9SQi0QjPhUE8mg7+tk8ynBxEiTpjWsDhG9gGOvflPamzBkuESbuKp4WDeMgq3R7cHGszQ5KNvkRM
97J+RJf0oPup/kvFhEULREwNiuSDOUk9fu98NZLQi1xITtPr3VkBnJpKPa6zIAjpzUd6L+Wife8A
zPSZkRStXnaKghrwRS39hfq+IzZr8ruyE8blz8N2pTg6yjJ0mYo0BpHuZ6x9uVg9mQJFmoJrMNzw
OhdEmdFFx0bVpCE1EtB1DVAPlJXUQv9jzpH802NNAQb2h4s6dK3Lus2j4rVqYKya7Ik+H2D/v1iP
nBfZrxiFKbQXNO/opeTwxKrMxxEiLwzm5wrDyIj+2L5E/wK8nWH31vnM4rEAX08ImTSVlU6tazRr
WJlikNjfy4XRT2rg9kkiD8uUbDmTEcV6cPRT4BUuJA4u2mFSlDSieRONIgtBPqc4rBbRfNZL4Sdv
XFUL9CIfmuo/CBTyyuw5SD1DnMn/rgErD5mxlAmbLhjTnMsF0w0iEwUqykzt4VWZmlHtZ3RMCtaj
XxUNOk4M1tdxDVys6NSkHoKCm4qw9xFc86enXRocRaAI3deybEG3kgFXz3/wI9wMTtMBpQI81WYJ
fmzETENhwfZrg9gAgUiYwCHq+Yoyt5XGpYh8/txRhHtKOMGw+YUTrlhYYQy5BHjbzHNgz1ifxSX4
kAJ4bySVi/f0aEIbRT3Sx2A/qXTZGt7Unl3a+V77kAwjSRUZbee+QXi/f08DegrStZAFMNG5kkGi
gii16gFMiHyDhm8wnpteHfoi9U+7yp/zrp8Frxk9giUl4QTZk59EgA5k+ugwm7Wuo4ivL7HoRUG3
AvtivaUS/R74Jwy3xcHOHdNumyMSS1+mDCNPurNVQncuxBdg4HdEfrkniOnVkDWUhzNot6L7wo6n
qsZ2o7Qu+4Ln7aJHYorYgMQb1O3Z2YaZoGAqC/EcAf1p0xxetUANs5dfhOu2Xt8KuAVLuLqy6UEC
48FGml6J6DJ+RhJQF96wL9ZY7Js0rc9CHAV7YLMGM389VYAZjST4pfs8F2mPCach81asdC3WlfeF
fDIbYncd4CEcnTf9tY4dKkYc4NUZgML1mtZnyzjnfO4xYCZo0qaw5GaQwuPXQfi6Jj+WTh4uBgL8
b2UOGaG3chqTLhtI8S0UrX4E6e1Pat4Vp/fMVBsBdS9GzhD6qnCb44JDsB8uXwIgmJSnXg7hPX78
2QpgHAjhrezd5p8c7xLzk8avAAeJM58ANfuf9OFC9bpHPAyZD43ZiKZgkO2vvm4wITPXWYpCsVkr
qhz1HqrNqXnpsgwt8Pp9/171CfYfMTHacj32TSthmuxod2IOixs0NmTdm8zwGIm1rQZUF0orsSgK
QM88CLLcgs8J5Izp5nYF54whDgW3gJMvhJelnTxKKfuix8vh492EXjr7aS+0UDF3UdTGMTUjiklz
W7WqyyTrV1z7YzKCrszWXfhCI087q1COePbsozigT+2fjBW9tfOxCHFBoMbJm76ihv3De+Tt+l8L
a1MILXRLhQEESeCrX4DVf7Wtfm8SF9a937n2pyDWLPCGgHwVLC1FEGOfxyCeaX7xIhQ+Ruy1Mff/
bPzwhOipetcGznIT0lqu7q09mDF3Y+qVESNe3V8H6NAN6V0sNPUS1yoAoVu4oxC88lSfo54QQx2v
qVsfT2znnFpHWjRtHqI4QSUOeo/wnqzJ4iG+yi+YWX0+hVl11y7OV026k0LSVGxSPY2aHonsIpqQ
pBfQy/9hlS2H3SL75Xv/Xj86yzvUtsVSOMgVS3x7J1wIRJM++mDgAB8AjtRAcAuE+xIK446RY7fX
saot7OKoPt/lfzn7z5OEafo8tFQBWUe3DhlFpTyCz25XgteZNTN0BKlnlONbEBVqUZu0+ww8cQwU
sD26Nef12e1nllWRBAExif/ZXnGAQMYMrwtAAxeHnC07wrsjAF9z/NHFdBlmXzRpJwVF7JqXI2y8
XGMdocINAvrFawa76Ow2f4gm/4TPhnh1egC/Oo37cVyJSvBLIapi5xCi+2Yu7b2r4X4MCKM5CtkS
MOrXqKgyykZ9Zp9oBwzQYXv/j1oNYa8QDdcS1e7vrPQBk8l8zBC4+nU305fSR+SsdbjZi2DZSrOC
fRCoeFaKNuffO+sFPpghIocQTBg2SQTSXWl0GFLVeONErp/QEaWOw6t2+WhK5zb708V0Kjr5IsO/
8FLxxSVrLJSMfUcifAqpYqGYNautmA6VVn0MmsJDP6DxpKSIHAldzORz/I/4Ov6gf5N9RliIKkNp
P8GsYZ+jCOUo3FFrdaJYtofNyo4oWzkIpXNy8hX8UVbpZsQWRAHVolpPGn5GWtn+y+mdgG8YFlxn
OO0JiL8HnNhqs3tGw9+31Jwk5+MvMG3p/70mNQYzTmUbKGkz5K+Eyf6nes9TW9v4tq7cjazs+RIF
hqJuH/zGKlFCwUFo2xaZ08CSpFLZHsn2B4K0UNSjN/DhT+Y6STL7u2l77yrIPDfk1p1+u2E1yBNq
ZkAl2dxVr6ijmnGCSXnlrExoeMPCPlrgz86ZwSAbSWTd0O/Um5YvfRcwzhov6TnuM8RHVCP9pVWZ
NQvMZYikxFoYfXYJTNQId2+9L8Ur2LuVqBUtLcC6relMAR3NG0TOuymAkJsWhjz3hEuoXH3JPVl2
lEfvaZ9TmNPTZpaQXXzLlIxP5XwRldPFI75OuO3cF7zMXqLQzdJ2Wwk3gA4ngvYlDEEUIRokS3H5
8Y9Roavt0Ie/yzWLxM81MONFyGY+FyIt1EC0iFUVMk8uUMtMXRLogeilqLtB7/mppzMBVgj/YUGz
Mxox9KKtbv8OeXgTJNGycgx5XVEO0kpVRwyVIzx0mwTX9Qa6KwggztOGJITpWtC5nhED/q13SM2i
hNWzIs8/3WBUc1jEea7lTe78nljZmbHgtPN1FiHsMGzywViPldv0Y7f5xa2rz4rfpijLvgu28JWW
xKX60xxK/u8YgH4DsGQhz1jPfkZhuC+TlwoxwNZQLgNLGdEszD2pKYBgYTxXKa7YyLRBgde8Duuo
eRe2DZMjWxRTVxjEPXdCFenWYr4wgars3Y2R280mLaKkiDc2eZsSnjoA68mthKMWxgr2bKSlWpXD
8QBbArr8yqxsVkk+M7Wlsp3p9SRosFydwwqk/a2SfQD4uq7NsV7tgba115OlVTnl/2cre6MzikPJ
OBpvkszEoCLz1hmv4Iq2q2J39RskQVqK68VEIEJY+M7/zstNsMDdRmAJC8D6hW7/2udq5QfXQKQH
kPpk9XJqc+YSo48klqeh8GK8x2zwe4KIPPMBCLZSowLivjX3FtD/DLOEpejYBN639eLcVzARt0C/
0phIzO6QYaIcUkgzdZqjpZTH8fCRDaZ3uOjk+RXfujnV2GLjBdWpjPZfsgtq6PQj/tKZYG7WEBaT
752NfNJF7/iVpfDYGNnItjTeyI5W/xbFxH8VYqkcu7IP7IWY/zDyHlWQrjMr45babYMOL817cmpe
CQT4fYJf3IUOLsrqEy4SFBYrijq34Jfo++LAeNRVGhN12zjiJpLhSj40fMWVIoOI8UjMWpk/6WJ8
V/6yGkJNOIQ9TBcgMy7Mxxd0wf+A2A49Ge6TCbgmniRajRyy287AliYbF1jtKTq/WM0lDbsPjGFx
FFxOP+SGn58O83sfSSdq/JeIyc0/7uEE5YZ0F/meJVf/B0tiTmb3dr7lmGRZKFkNBp432xbTlAfe
5rmzSy9QsmICqG5VKoOH6Spre7a14fucFk7hpSdKtvIeuK67nE57PDNb8+8VI9lzsNb9+ELsj1Re
FVIWSvdXkqs6YV+GmWKms3kZwkEFtrBsO0Rhsy5qkqOJgypHlH8Am8D3WIxsIvRqF+y0QTeUs8Hc
L8OQm2aZhVnTgbK85fvW6DFchHF+5oI6gD7S3lDKAPSp1tyLKgd+oOV2ephYyBFcAJjev2Y8m+KZ
aJ5lcFVELVd0OxnAtCNLs1ZOVdPvSiRW2xhadCUhwk3pZC6YuqS8lfisXWdnILC26DTO018D2Hla
ho7vhfEu/S+f4wSPxUgkQ+3Ad4UOjI2ie7irAYlJygkAf4Nd8geCpSlTt0zpe1wNSc4qqkTOriXs
meKSNwAnm13rTPFwJ7tigS5GzFIuEQX5hiLwAKvlOQobWIHEIcV6Sgai/SG4qerEcRuptaBArIvP
6qgGs46xzxFGOnwH2d7zsau/e5l4q5z3bziy8s4zRlcX+dHIVcOoWwKoluPMQ8AjRnc+h9XU5ozn
OcHfcqINO/G7a2D19vvAFUmQU3YN0y/bqWljkDXJx4UaNpeaYzYym7yYLtvhxH91pVuV9NVvzM0D
n24+w8WIAUAacAKOHGkpsvBeCAwkWqd1NTlKtGlINZG1AM+h7hyPCws+gLppwW3LkL79yjH8/3pG
Oydro1LjL10/lp1ZAV/ZFcDisblK25glttUzK8WGdaETT5DBlURbtKPJO9WQGkejGqLeB6wPiTEs
h7afPH6CqoawDI4R3TRx5aNGhZh3eRwISe5n582na9SGy7oHPcpqBokbubStgm1fhh7XZ8NdVqrb
ZytDZO98Joo3XEjiZgjoNe47bOnSswmbmNpcNjvmOYwwmnLe8/lcLbpKEJLkxFcQjjqBT3PDHTrK
XyEgb/zXeBzLuAGrR3aIt7NWcbRQR1UTRWYfBq9VFu0ib4yjLLDKaeniHRBSEa5LD6t0FwWAsOY9
9Nk2jNtfl+lTNgVdxlwx0Y6OWpcFdQud+hTJDX/6X5STmpB0IETXE9IiMiJsx2Wdib61OShcAOq6
o8bW3Vyrc+7caDv0sIm0JzUkSMYtsjBDJ0pOoOR16n9e7pBWjHk4X525B91o1861aJgdo+AYo49s
3IxUH8Vo/SaTreFVaSkZdpokiOAhAin+6BW6++Rmz/3kVCmFxomuna8WX7X+/QjK7OvyYg7iyDiq
CIvTXoYVol3l9wEEVB0noPK7xLj8ka2DOx7TYINm8dLNhWQC+ltIMN87r/YEYbWewpBYIn6NQYTv
DQ4XZHfwFx4ikX4DjcM34Gme1dvRMkVfPxnZlF8yvFax6domM3DRwFw5tSH4em0uBrCPsCEhSWGD
VCelUy/CcqGZAilp5ckymWKdTwRPM77hrMk18Bt2jVGB5eGlPl9xn/W3O8ytIt/eXHHVi3YigbQL
KEOS8WAdgvqvIftsV2NpPRhZuhxUCNsDGWLIsCl8vuAPQGx1ryX/PQh15Zm4VE8gPh+DmjAmov93
hlMStvS6b67DIqXt7mRzEU3Sfn9O8AEiykA7IRHggeTriskZ1DQBEA2Vf//BTPLgEB10rGBOtN2U
qkJnDcVHMPtj0sBobg1r1IwDUMX7hY/5P9WH/30VCK6L3GvBbnYGRuzrrcXIED3JNGTEnvkmew+L
SBqWS3Z+qnpYS+2qSvSjkkGhSa5VTX1y6ehep6z33RLum2FD69tny4VNU7DOdihO+sZgtWG8ToZM
I2AZSv/q+Yp9Xj27DyRrZ3KAI0NgwI7DCRuEPhHiSzMXedJmocHGT5U3MAZt0EYVzU8rbUKF9oib
2DaL8EHtPhCsajEIy93CORf/l3VyeYgtrD8cZSqh0x3ivklSj/A/kAj9r2H6b/665pqb9UdiRT1p
QZn3VO5B3iXQoRe6osQvaT+IYk07ICylqM6wbx+njIm5xRPu8PQAyV3zkoOWWPe22H2zIJXfh2+Q
5LthIf968aqwUtq+k2gTMVNcRwBqVPxQ8zQIvrebNt46b3bsCngmQxy06L6B/7Udn/ygnf9Ygion
ZAExKLxjtsqJRQYHZnvP5yqK5v1PTBOKKo+90A4Whb0hQcBnpgtIzlBL4QyTeq0azIAnq28pi90a
m6bTCJ3tLn1d36fmxKz+wQU+iyXtISIQxBN5oYdEMszrXVupRQkrN+vUj+w1zHcSSAkahWqgNUjJ
Qg+j8zs2ljYYpmYRuzh8RL66crVwftM5ZwwQTzkbyYJyjJ8aJKjc+4Hi07f2es1yVAzqmIIG2nA+
2e7PzhA0qmq0u4gIsxYQeIv/gArUR1SqJnvn/gosbdBRmc2mml1rDfoed5ND5wpXwu1nPquQHoaL
/wxREDQ9R2YczZCRZqvZrjZxxfxjS23O1TXAlhxEjfzVKkJ9HG4ROmZgUM3woU9g307Rm6Hg+spg
2qazAdQWA8o515t+qJgGGN06xBbi8M+cD7xbQ9tHkcFSBvYANQB9dCTheC7HvUNDWtKKqKbCrTZq
NtULbmeFASysAx113Rp8gS5yu/TJrvK4PpIy7/2QR/jfbJbOe001ndQKkvAO/+9Rk2LuJ3TXGARr
8rUAle+GL8mUzfCyGGnWNnaKloBCl2TU4LE9nxlAPJm6hpqJsHRZt6pSvoFXND+cstSvGseXhNC0
qodcGy+r519GzvbQfvzUFljWf9hhtUYIqCWJH/gRmsD6zNeR7wMm2+Qzr1tC8HWo+0gYNiEsFsW2
BTyfjdeTKas1wUNYxQ/JI/iwwZek0BV/k9Hky2i0PJweARSrxYvZlJ2JxuUx1uy0NnKUUiH65aUn
3OGna157yaEHmaxkrr1qFNUPywilIGcXFALvsoTnX+6ys+ReFYDo/NsajdvdTBuJxPx6Z1O0yiQp
ETH/xlGRKMFhySTPmIuoTYB56nnqNEeJ6AJG6ulFkJEg7OpJPzfWo0jlLOMPxyGRJaHgldkkh8X/
sJavdOPqmNoiPIuRHg8x0XWQmQQcFX7mN++k0Ay+zJA4YWgU3Nu9qVAxMYlyCVWZyZFl5hBejzYb
gAtKp0izm4Nvw9B9kEg3+UhDYconz4sR1qTwmAxP3wpZqSz/ao4raIjy0L3hCr+qiwdCYtI8ORGx
sRuiq0zAp2hLgWspsfPobx4Bd0qLGlJjqI677kqs71zikUs0b9KOVAarQ9NCgXy6/+fLfpBDRzyP
G1TIQLZtb/mBXK5CKnwj9sXW3KxSX6O6Vhh39B87sGbOJbjiNwbxRm5m3V8GoLiICYDyZrs0lZdY
Vc/kE9/E2yBYMoacaQE5CKbLz82h60mBf6x1oUI17otecFDewL3E9ZUlXdR6ApRzHtA8V8HY4pLM
gMplI7Vy4DNt/ema2jz/O2ag955gc8mxM7qtPy5f2iR5Kynz/4aE/W6K7UlMufG8dN0OWpRv9Uqk
TyR/RNlLEFqfEt+FsqKNYOmSRmZT2yLy/2AtTY8nuEE9kK7caX6uGzLERQUywGnS2lljGiL4b69N
v+cAb9q1gQViJRibLqCLDKJln91oqDe2AcY3CkMxiS0di0VelUzlDC1E/y8ZKUurb++hn07ktFhm
iTGRfNjn6biGlebepsl+9+XW4zaZ9wWJK09klGZkzuOo8dNff+QiyCGl2IGekLZ55wauS7drcIzs
YaqivKgz9ofZAzrhdO6fHyUFfI1NQrkLokaY/5OpExFB9yrt79iCygNT30UANlH0AwObvFx+mZYt
PHWH9HdaDqrLUuATPLRI64iUKliQ9hpZHSMRBX6s+UXHAUGfCqse9O2RKfLkPtLzZfDAx4p5aibZ
5evPGBcUV8DQFHYwKSFJcaSCdpOkguvPPqTVJmR4uRkRI/Izzsck/JL/wBDAS0YfbkiiEMsfCUq+
7XwQ9ECT5LnYWkBIyYFM3XMNm3XP8PUFNV/5R7I8brrK5AHrglxTH2ZRHu07iPTZNdNsAceLuYl6
CS0rnkky8vQPDFelJCFanHMnkFerrL1UTYe7g/N6YyjE8b+/rQNVbRg/eY4gYB5otzfOtGzZVb5P
zHifm8MjW2mP7QKjwWKonQOrZ/UrmsHM+7cNEcskwuzthdUcHbpIbyncsbr0z1PrDIfUGa3scamo
GSdlIkV+w4SXHUxrtTXTgHEO66+qCo5255jXiQp3DuC7uu2Dl/fJlupsaadYiCniK/8+KTxBckBd
yqH+afvjqpRHGABiwl6IOaG7GgTIT5SBmOLU56fX9ZNo3EIP7u3M8E+0DPhiPVXnAbw01ZBXWv8R
TTzuttFaEjTNjPcHoOXJlFqfcNJNVKhoHqC196H5tn5UkAptR+BNwFkhoihT0gAQ7YJ3fOqGEtSo
RumOr75ZAUPJUcHARRyB3dpK5em4TGPzG/JqOu8I6WVFCgi6NBAOz1yQ/mEVDCOt3OdpaOQuEGxX
NVQSR3xi1iWU6SE/JD8ebRkLzrjI3+B8IPsjGZsB+Geai9MwC4eD+QDKH2U8C8qUBGGzcrgiIohk
8BroopEx268GaOquJwUW+16me5n9/82NsI0HWJ3skfMIwyBw7XJBGQ5rQlS0Zf9J+u+/MsCc5Mk9
bTOHI6XDKC+4vjfPHvPX7xJ5NrQzWs1y/KYxvyVyUXGQy0jQpQyQ6dewZVz0ulHa4TLtjYuxywsk
X+hLZ9mWgP5ESx0PwaVJgUTT7BxeG1jF/pU6KJwyzKHObpdQia8fMMQbLRK3XQVpp1/WtekBiJQ/
kzhsWr6OtGwcTKYI44EAhj/gZgRugJeGfZaItoUU1RUyYYkF614RpQ/cVRhy7XODKV55Cpsx5STo
n1nWLY4K6JbxlLir2PRbzfj5oIswEDPVql9uj9oAbI+qmpZyfhT6oeuBdO04DUiynVB4PCDHReOT
NB61r0xvJ9uiVRaIwiu1101NIQau2LBZkG+ZNSWFq4SJ1Lp1Ks90PWL5+15DlNZQtZ1InLhF8SuC
NW3KjTgjRf2n5FMrVDJeN9tQoSImfuvw0As0dhAcailOsTauM+8elSurGl5lzuKvH4vp2MbflkIP
echITr4ItWf3bRqHFvuvHLZx08lpQHDA9s4B1IB6oRh5m0Zvi2Izm3W8PjIGO6lx3/dU6qvIOdqb
3nX62qZxEcQtT0M6AAyNiCcLmtxr1kl0PAfQgJwX0RA3q5gyx78UMMU/EkIU9NW1xgf3zD6ctAjC
5w/K9Hy2qm0WiY/CpFpPimD6AWlcTu6wlP7V8J95rO3MxA6lf4ueRH0WU2ckLhR1Xlg9dMVjwOY8
/8aR9I+7HQTNym30nAigAgFcB0jcTT1YO1d2NbFTjX28zzxowQk9jSzb0AG/M+P2qiRkR+6oYPSf
OLosuMg0f38z0sfKNChuxU+8oNSRJg2MhTOJAYeqvnJMLvrOG5ihrVicKw6Jitb9bzrkSxJkxlVM
05CUOG7plDSyU8MTlOOVCFIUBQ9PuaZuz5fWkL82DRS/7uyI9ZkdxOlEQ9/FmvhGJS4p6MGgqZAW
buzK8oy0jRSgQXwy2Bp2V7+luK4oBt5SFq+9qQPjIW926Eqy8r/n9cgynVu4XE/j2wz2GclBqVWU
erQcz/wQuKkh3WSIkmpdo13jVxMAd4q3w+UFp+5hQ3hCV2AiGwOKTkG6JVfQIAhS+6daVVHZHET6
elJU6fr/Kc7I/awbJuUZQ8qe8lPWCUAaIKxrf1CPku6u3hb2koVBimQPPFzupuXOXqQAe+AU6iZZ
83txJdtaM/EKUFviQpUfRI92IkM8W9GzNxXsXNQcN2/snRovXT6wnIyKxmlXQNZF1WxK8mPwrVf4
psboYLMnKz+WS7rMvlogxHNzkDLReHeTGqjhCN0hl4IFsCD73oaDSSAQmCEyvJ8Xu2zr+Pq29N5S
5L+q7w+UqoMI+NEK9sdrEFkd2c3Hu4XeQwsP62jkobFWp/2hwwhffHRNdvK+UAqa99/JQoPDfoxG
3CoLU+mLHP9Cw7SlaAXjyjz09C5nY1ajdNEiSn52DSmrg+W1prUsHC2DyGr2CwIDpizBRyCB3W6I
Lg3WLBwpnM8IBs5CKP4q+X3YxDUDHRQpvlptIPMDo+kUwCY+e8R6Uio0CXqHQ9LSzfT2fUp5ied9
ZLNNn5luAzQlb3zdf5EGucZlmIA5hqVOEdIaDU2vNw3H4fm9ala520Y/QtfL1dOYVGhVou9vhVIK
ww7YS7kW08cR+ZMUX3J9skjm1huKDw2d4d1KaS/Ei7yohUgZTNjjVcPRVgx8E4+g8S9H/5nB2Je2
CEzzumlNp/tJIdOrdrzv85xZZwIldweBnVbuCf2GfNqVQ4xiz/LWBINFeiPx2mLhzohYOdlKDvSB
pv/XN2OBiNg7Xodu3rjeLK+qKvhB74fBTWQivKmf8mh02WP95gI3qWitKH7GQpqxCajBIZ27X9Fq
mDFSjC3Zp+dpafGnFL76ukjH2YcVmRORERtoN59f1j1r+32LKn6fy9aBEf0eG7WyXxb0WZ6qaZDe
KsC/9kgl+jQKABkoUGbSvwyU0mkU/wmJbTQ09PzE09rpaO6UpHY/6wv3lLR4TZnee33TEWSKAw1c
KM62vBHnFlWm0WbDHEV2SnL8WHJjteCZBG5LwkhfT9x1sTFlzXD2DEe4/F6o5o5xGQDcXSPXxi9d
b1nRFQP1LCLFyDXKlz1wYaMFKDf7W94bC83hOqaffm3V3eydgPZaCHL79hvtMWIg0H+dCn8Dfq9F
95LHqiCZZneiJk7abxMbKLj+ICDeV7AAYZxdER0rjaeFdQLS87tBqn4ydyHAo5PAbk9iQaNqAs0X
t0DtKox8fv0wgBQ5nMjrsiMLg7mRJp5zopqyZvJx9nro1EfQ9PT9GWeB/niHc56Y1J51t2uBRlfz
4VHfXedbDz+ghbivhPMxTqu8v4DG9Juuaqzvrz6REZ0cNDSE4mPxAkluRqKhK96Gy4uy9Q1j+QMe
Tcg2iUy+s8WhOi+T0FEeM52fGqttq0Ut8ywINBJMgkav2fnxeTne1Yy0qu/P4/AuUWUAq0GTEvJD
HjgSZQzhVeoxSNF3pwKxAtNhZROy6K7rqSTeucQQ9t+NH3+cFd0Nct9ya/WmrydtcY9jKTuFAdx9
RZP1or1VQ5G0tX5zblX/XI7/jqwck/zHqAGa5YIuT7Fbl1lj+u5fwnHZBYGlOkVZDtxRWehdyoi2
wRNfMzHbRijQLqHUtKmXU6nXZeLVDdP2oaj8z9NAQjPIIdaHKNeLVnaUUwGyiaoGCon8YKvqg7V7
Ow+kS/mL9WfhWOrTK1VN0U81XypywAhdtNk/mjcKg5fJQWutoBMVoijQ/laLwqO35sMPDvTakyNy
Y69L2m2xRU1qKab+sps8JHYyqT7+OtQFduOqw7M0zTO2cIu0jUeCtiI0Wq9ehR5/90Y0QDzwxti4
SMdu87CXwWmAycJn2vrcNyFtCiRC35RqPRuo6N/sdn7KIFE40kdnCdSWBrFb+IU5ZVSsnRW88wSK
mDmUIiNX9VNwrccg5IslHy+tN9c/GtsnOum7YziG+vR8SjaWzO6WO+oOhF72LxguUkBqUYH3dibT
iI+HAUfewr97Fz5cd6qHr8b7TwFNHQFo1J6njsAvRodqTWVm2NpacxWzUA/688x06GyWx7pM3Opm
Ct+0YlmorvBtBYxgYnl/64KeXuw+LJYHjd7HUjZFc5bqXULgh6QlqhrSF8EEZ5I/pTtSXY9R7jKO
JVHT+ETboN0CPsEdnMDhd1zkGw53jQLdmqb93LiMONAYq7op6bXN23Vm88D9CeahB+VA1B5IaxFJ
awNUbvnWeY8UZp46xOb645zkG+ogHx8rtw2QSIW2f859I1pY5S9QGOka3ipXkUF02AuC6btLvssT
3l9dfaQIjWpznpCu+5iTY2Qomdi39HF8MDvWssigtchE+gvgGStOrCk94ckE4QG2vBY7myBU+CVJ
NqefaUVrYoUlesT07sXPXCrOYw7IrjM3wdfcwB9jFx6RKY4+mVTGUP7iSqIJjhtUadBT7qsPIijT
vaVMNtougWZAcntizoLUUlfxLqN65LHA8ggumZDY/JTGHn9Lpz25oB8W+k41MZ0RwIo0G85yazO/
fKa9ntYdZ6s/iDyWKdiMZSGY/clX5fyGTw4fFS/CEXmc/vP75YyAmPlMUobW/4oQyHxBhsGhW1ZB
hCpupvcyxvyUgmOLuKLQXhHAn6Z5eDNNfwjNexvK3jR9BXlkMCIgp+yKF3TE5PkCRm79ex7m7jiE
DpZBNieh8z0DFndpKtIRW7sv4hESup6F7Lhu3dTO+h3Utm1updOD22shidGhIkfuVTEXiKHNnxsu
GSItdg8OQBTUoPXV1e+aP/uMTQOleYrknUgxXHXfx0Nhcf3CDZS/A1HbqItD+4yaf26zQG7ZUZrs
7QpO1PPp5t2i78h8VbLJbCNI6Mgr/9JwmZaVKLenAYu6JInsfU9g1bCZvllHO18pDX7/+gq9KttX
SPWIkqqNQuzPxJobAhGC9JWmQVuFzLUQmGaP1wGT3vg85Wd3OSRkDEmxR3KNLfxQT6sknH9wmza2
aYg2YjtGDilUOvkTZRLHMD2jRelNWonkfcLa6SLE38yeCuGdysi2g9T3buCAHmK5V5O2uv+h0kUf
73VTXQCi9LCBEkw+1/OrvB6G3iK2ZpIL+1I26w5Fcym+ksVNza9hE/daCVUSbIdXbklO2+LbM+2r
EA2gUgeN8EEV5bqaH3BlIvwtODZWDygArBjLhj2vPPRcW60KHQZQ5Ocw6NeOeHN1M4NgjH/g555a
JfRNY8COrnYmrsNOD+3ny7jwfXzuBGX3EBD1n5SPs/fGchqPW8kn6Z3jcsngA04sdEpVqYpeIHBR
I86Ss3bYKEr8rhm+75nHQ5YUbNjnGvguFpRxxqvGD4MCmU1xG/+WaJ/iwqc+fciQ+NQB9uHPbhFO
M1N808sCVqz15nd9viqA92KI+Brga5Q9dNgCx0WrMnzdCYxXMC85L1O73BXRWkOUm+cEFNV4h7D/
On+FMSXCiCrccxDpGmhqpUMQ633lWJuZlr+H6s7W0i2pOc+e3Hh9hUISSindQ7/i1OdmqxmcHn/0
ynjxQMZnQzz/G/s4bGMlRwXrYJNuOQf8aesVptXEyuJTUMDutd2vq849b9oiLaAdfVga8FfkZpb9
00XzFkR4YnIo7jqJR2c48TA+TBAKgpFEPxGeYMFj7Iq4mZGVb1glYNsVUUYLM68swJh9INi0tscv
vk+TtSw80c1dUxbYxxdfR7T5yahfBwmahCLHK6non72+KBM9ouqpHJ3tFRtl6WHVnCfmSFzwgcVY
t/yVqNYyk+R9poWYfYSotbG4u2l9OYjR/bX7XuYBw+aejDbZVThkvKLILdrhHPd4hewwtu8RS3xy
1Leoz8kNt99OI1WYQteF6OXuCak3fVrg5LBlYN4AmvoJCnZh1exiTfaOvbz6fABl0wt4AbuPD8W3
v4sPxmJcvswFfhg0dPp5AHiJcX7gzyK4+0tWDwviSVa+uUPrmqDoTm4R4mkNuiZFthbanrQpofFf
hAw5F28YqIL3grfJZlTJB3/Ji5T6v1xE8ES2JJACFqTY6Uwi1r87lVl3TQ5+jTyj53C51m+jeQmJ
HkK1grisVuxkoJZrpY7su4nQFeE1Fx+y5Y0KosZElHJuJsR7ZkG8aYncusOxR+J2q7X1hN86hLGh
MossB0rhGwXf8TRVLvkEpVlfCg0qEeZqJJop3cA/ai+4TRA/Q7DGE/bVAmhF02u+qLoF8aI90Inm
CkbzRwmfObS2ID6XoG9ycX8zag5F4IwFzPEvsuQ2jOEqsBqYI4L+r7fzFoGS0WxsiiCmZcQuy8BQ
jP71eBe9Exzu9zrqMRdGUhO5IHpLPGq3yOODIpCHoh86btrCaQTZoOiF5QGg0QkgC09adY0n4rku
t8r2tvyeA5SQczNHmGXCx5fSTCQKBzvKl6tzkamXPVpyF9dpV5IM1BVI7kITqDi9uiokldZbTxtI
V/QyhNeIK0iBYTwFBBoQ4LYOGAoJMCC3hucFjJl5ryKYUFCzuRgJeFWA5uGNuXovr3A+rXztONqw
KvJaUq7UMeTkUEJuVWVAaf14HLmTzrqN6Udm8nn2D+kyCHfYHOTh7aZ2+xL/uKJa9zWNKCs6/App
/hAGGsR1WA/krxYXkPBdzNHMWAfY5RFL+3+2GbAEVSQ08iLqAyLAezmah10IhMz0gicm49fhg0z0
PVFHzl63MrxdJKWCukXYgEWWy7PqELFGvvvS0UNYJ84TAEQ1J8yxiKdshvy2gq5Zu0ryjUV/npaY
1KdCr/2zRkdHZ26hoirnF5ubdEdTM2pnk0pT2b+cTkEeAHad5vYQAZIroxiB9ZYqE3jlDnbphTyk
Cz6pHzWiCcHC+dXwxvX3o1eP1kXFHJC+RntxfVo/V+nyB4eaABJtIhe8lqdxC61jDre89yCJzbY9
/hqGCe2zNvVHB+nMdHVLeRkgEQdkvhGYz9svHA5VJ4YR/misoqL7LRpYdlS+BkTDdM7AO1MUZTwj
FxymdNxo65efitbkdDeqqGchhwtAph5GLAZNXOi1yYkxPvXLiBbEWwOceNERN4Zq0KnC54Hq9xnb
xndtScAvXdrZiPJd6+LJHjq8R+glc3eirFiC0Tnt/OIlKsRPC0Esv6F8Cv3pyMXp0bAUARcwWAng
sAMh98CBj9E44BQa9NiDnLL8gJ1ouFELKV5VitBwkNifMQzqIkRU/A4/ZkUcp+YaBThxwXgWzuon
gbPdQaEyKOhomQoZl0GheO8uRbbEnjG1tCjSvcenaOgOEOfGMrshVQz3A13mB8XQ3WHL81AVA+5f
QMZNPv+14OToCV+9zDwu/AFrjukWkVd2O71jm62rEnHEdks0GQbcjIwL3mqdocM1xo/DSSdpct/5
0Tx6Vu8dE43IISHNs094JDIy90fZEMNUYNz0j4z/8+WXcyK5d9M1ToDR6iYTaa1i+ERsyM90Modu
P4zg+7tKM4aVeNdwH5v+LhL/upZtbdg7/WrWLzF8IsDcJJoQpS8MowcIT8mFEF6HFzKJgxmc8VS4
vkxKLeKgiQ9NqLMO5nM3Rrcrz5m8UmDSJQop6/BPPc51Q4SYTlxq5ZUG7AO1A7c7pjK6/gAb7cgM
S1UQN8yhx1jEhs8DjlxgNHt9ADzNqI44oDGTmCBraAn5Udf8zyG8Fmn1IlVyWM+Bc7eeExkP4bQ3
wEuZI/WxqUm8Cn4P8JvY3O/rh+RAyamo0q3qYiflmipez2Qka89ic/qYQAXRzzrwZnx0BJHND2kQ
ZaxjkKW+2knzsdjQfrAsyY+MnUE1TAcFpb8RoeBpvPvcQfNTg+gHpIpoQmDzrjZsibq+gtyQ1sme
eEROMyllf/pqfcw7f1uRc2TLSOvwpQDHf8XhjLNrtzOWNij7PdYVh7QaGle4rdwhHbFnxKD/ZyCC
KGCxumNcAybBAYauQEFUN/nqPvvc6WJJyLVKdyUIrUkJ9VxJrPmXhZJ2oQmcYy3T+45HOmfz0f09
4yKet46FIyCoa2TbwVC2DUwSinGFxIh9xHlSgCzWFoWzLl9W91I06sWNSnYAOIJgEBweVBzn+oUX
D5j8H2tU8ABHxTdkbKU9uh6JPuVzS33yLgOMwV8wqv1FMpZifRyv4s2dB9TvXskKy6EcwD/Xrd0B
DJfQZhoFCwtZ8KpYAS6/4o+yWgw3FfRbhij/0U8vNxIQeDiTVUwObzzAkCUbOe2XjTXkk/eiIL76
cyBzu0KlHLTWmyvCLjpj67Y5cW6aMzdf6dt46qOq7mVJhXkju6BoI1sjoehTdj/cATAvYfPmtgfJ
iBscxk89L01sCqDJx6reXd2s7NXdkcFy3ggdfoLTDt9c4QsUHx3OCCKI7CXdXK+3Ib9OdFfKWdKR
fRB+bk5rvyHc+h4nztipgY4EFgjGdDDWw2GvvhJ+0QaKz8Y4iP4bz+eLwM9xRPZwQoLZiSvU2y6p
yde+eXvLR905RZLAN88GkCN5okIjO0Yk1ybY5O5P8rg/G/xFmcxoy4bFHFdCL7NXprBphfQIv+a8
Y43PT0ifwoZXVYMnb52JhKyG7zG9nz7h7IxmbyhVv18miYayOU5TaKDt6wsDbH5OAqtPSqLQtMGN
Jzcw/qpHwdBqy6KWdLzd3fBr3w9m835RY+ot3EaKLkou6ylSRg6JpLiPkumrskAiEy/mN9s/k1H4
VpFbsar/H+imIDf5o3DcwAhriPDLhaYlISkh6L091NYiq0UJgmwFpbH7KyNOUwASOQ09B92ZLWHU
rU9PvQIa4x6kUcUPEAYVIcgssdbE1+f+H5ObYIeRsSnWeQDdFwGEYRNhqoeqwXRSavC0CsFJknFw
JOiq/Q88UROjcQWoKWO8SSckI8w+Rgyota0IZiUTAyv+VtU5meHj+GS5/2U5erEy27xAY/PjgGwx
TRF9OF8WedEdqkXARk/rC5PK6bm8GCsED+HVZlm5P9cx+AcerFlWATmHLBRuKR70dDIulo6aWwY8
9YnplG9OHvPCtC8xF5Ocrvv7oZxWGKBlShs5AMPtCeqRxGrZEcZbhHm3l+pfqHdEnRTrpKpYPCPa
/ZL3p/3js1jdDdPuabOrz3a/eRlxwU3Vuxoe+J6jUbn9UF61rzEyHyot2GdksPQxIszAeOs6IxWA
UjMXgRX2jiWfhe8VuF02HrrbJBYL436eo+GJdKbDH5qXugs8cbVq9WCzlL8MWpXXpQ/loORGyjQJ
MXDYSr/+3/tbQrh01MwRrkecHrtoon7J1ercHloxokqXxC46ikuZtEOD+308s5us/F1ksB3Vuado
tUmpGAuyaGx75Iw27jSILl6Hyg/4xmPzWb/5G+kO8gfIHqJtS4L2D+fdKLrbncadqda7hEnKY7gL
5D2j5TPLJUG8P+lHAhfNbU1Upen8pxMWc1/lKJLlKxbxqxn87vZ8TGgulB51N/bxusCL6+4XGrmx
UeS+dCJdAGTYGwHIEvzCuYL/lEno27S291C9ewy+0+x7OOVAqMqX/dpwgmR5dLo1WKZPf++XjHr2
fZRHWJjGlJMks9zk1NJvkhR2WYJpdKrmv3NQ03cLEJjZA+QFg1np/KPL6cPhZJ+/S30AkWWQ4T6l
zzW0uy9wHaJf6QL6XHAV/lFyBwZScN+rVgQCR3TlAPe1xXswY8CqPS1n+EhI+4Pb0xlhR8TF1Pxl
N4vVVprlsmPr4nAVHHK/4+OJ7BsuCaOC5WlIDOueevdhl18pmNIqI1/XGW9X5EWnMdHQVWKEu9VU
aIhaeOgKI24EC6G6Zh4V1q3ZrEm3aBtSbgZ+hbMfSvYh3QHZaSmDwY0yRnuTpvwmrIWSEaYJIMtk
WNMTRazCJf3pnp+fwxeOEYGMf+V3VUq+U/zbEDVGtOoLuXmxrHFiDWlDzCBHnFcAwHINtTOyulgf
Nbvqd8YJPC+PeznOUMIf8pQa5dHlMxewemWEc/8cdnxc+UYBEHxCA7N2Mc93HZiCw+LLjPZfo4fc
bERrJyK5kN6FfYQ6OhoZBszbcGFf0+3dfCtdFzoK68OzqIMEN9zVSGvc3iDGG2FTxTP7AxCXhYt7
2Lh54765cVMr77nkZInoywOqQzxKyfeTTuYWrf7ceFJpU8fmJCTDGDpeEjEWXDLNtx8cWF5YXzEf
MEN0b41FE5HAkZPTcZOk+OQvXf5nXd+21VSiTbYMZNBTd21mtFqaVE7YmjTpmQSEaiUTvghq4H/E
Cqy68Rmt7JNVNFALatG8C6gIUdxuAt780bd07c1zXz6SJGQYZDFLKhbRZvomLll6OgGAN21cUlyM
2dS2iUxFim1jHsBVTTySTPkaHYeMX1VMJqJGLpxeTsh6qJxYEMrvlVYWoAnQtq0rHG/Vn/scsC4L
rPDddeNT+uq+s+sHwsPvUq7goYqeilktKj4N7ZoWFrugJpuQEDlGFcELLODuDxD80nCFSMUYCUlN
vALO3T0VqZzp0HlhItTZbzW+m+WQhYtlb5UQ10M0r2N+FYBwPgXTqNwJ+zsolLvRx+8wW/wCmEW6
Fijc1LNTFV+LSM5wFHV3lX41brgCAp5Vsd5bIlhvKi0Q+iadiJFgGyNwC006v6SPxdIKLjnmdWGe
kDNfCSELxIGRFq5Y9HsSGyX/D/WyR+jAidd5jrlmn/BGNIFeb40ZUZtTY9cEsdznXO4yWjIIUcFl
yy8vCOlMIEgatZdOzOFaabxiP0Svt9GIxB38Wt25PQvJtNrIAYKHnpo/v58UD/NZcmqrYOuImdx3
N43tbyVbLdJhsYVrt7bhuUbn1JHHYW6LrlxworWxw0PwI7kS4qYsFm2pvcnou85vU3sHh+kkaaPW
P+Zm6RdMyAcjH6L0zraaOWkWT44laA33FEO92ynT3wQBGHkD1gZxiYuLnidVhAzxCkQh/WyLeONM
PtQ+e7DrkUlljnhXZZkSBOnWt6Fto3jBLYl8Vc0wNED/ycKaN1dQJ93AbvWWeM7Sskg464C5mjC/
rlcVki9URiBHsyxMFB8AI3LxJ8ZIPmey2K+Fwh+Uw+EaaDQ3CW0gB9PF7KMk9SlhBCM70drCsTea
5I9K9et8qsrU4eDFDAJtF5ylIzspWo0nBgBGQtfDDAI5aiHQQLeeYiEx8ATBqhfDCB60x3lf7+bc
+eAFhQMFQOMzTYYGQ7JVjJyWS2uzdPILzrSidQLeLDop7FZ6mmJu8vt5sxjnk2lDW2uLTdC7efc7
OtFkyzCySa44f55M8lPUeIIdBRkYklF9sYgNaGXa+gTX4fiH+9JJqX5ZVaZjVbd3lp1qJOnsZ+v1
NljF2Z6X7S32MUzR+8lMDv6n3KaiFkCuQnkaQ64WRVAfkwN4NepwxdpognbmREKyT89+Qk7Yt0VR
/BonQ4scR2+g4aWgHK30Ebkg9mSX8XRPmV25/pVsG4ttS0hBa4MFh4atZYsoo7EUv/Bys/mACpGT
sOf+YVbtpdhEOq6+XtTQt/VMZsZozuLvN/AxqbV/Z/wq+j4M4ItDorbzbqRe/9KrFpxFTzWSJUbP
dLZxifbCf4tFEnk8XZXGLBVy7g1zxNcXXvz0VJUn55T/5IPoXNyZgeuzy3hQZTjUNi5l72F8bnNt
yZ21W4NiCR4gn3zXS2l3zKP83PjoHI9HgOcWbZsguqvub02bwDK9mKyyYDxM54rArXdRiDGIbVje
YjcVqtFBGAsAyeS6Ho1vO4eU3zn4J2LrdkyPzewEJ58wfVoBd4ZNsDrCHkdcbW74V3Av/BHSgLGJ
IXGR9qbf0WG0Fq1gz+JoWsogIueK9AGA2AUrxMDnKJIMHc73mDCVA9nG18LAdAswgnU8KpXXeFav
lPoaXIo2tHuVCAkPzIZ1Z3RT55j+KsQ9YokoVf/hejrZ6BZkimvRzKLUepMOzT4Zlk8jYXoVps7H
dzkA8ZvwF2uF4bUT3YboDHiZaMUHH7UBx38yhFiyF0cMpMt2kgT+U8DrZGQrGn7QRHZpCVenp73c
jrmvw/DQzL3O3nLKtNnA+amB/zhUjGHD7RWC09YzvUQRivewn8VnZPPMXYxHLSk3x3WuA0roOY/Y
2IZu4llgYir1j2vBUtBz27xDPj2Y3/QbpfYHAuL4HhMHZCIXHhVBpK978rQa1jNQhRjHyGIHHWNM
BATWgYgakToEGwTS9VCN2lvqyawGunO9IZx9OYqdVLokO8T72F1iGeB65RVOE5kVDmepbnyHPAld
m/bGf0w0Pu/7hdiM7L9NU6t43HqUv//Rhn+mRegx0IFR5eJ6x/ce+zrqAzyUqUqXgVG+xxMgFpij
/ImHzpiKfRjK2g0AoHAlsd3HO8Hp4Xawjv9cb9OTDiDtl3QxMBBLqZ27TmJCym8Vscy1hL5fcU9q
3FNfQfrwW9sZ+HwJAHEnwinMguFkAKf92u6QL6nHCzvUslcQfZX8CxZPqjIQ2g/VXRMk33KAz5iC
JCAo9OXsr/0iKUNYNi/PQbSqqLFVoCB6TOTYDTTYG4bN3rjeJTqTDhJE+DCXohEf2GSHNINhd91W
dTz1Zb6THdKgr9kKAYfrURhw60oABs6NpSUSwlyybBE3yyCJ+KqowEltr3ado0RCc+UdBalQcvid
51wkY5RPwuZPmC54vuasjYUBhDz07HdicAdHawDyaluiRGQ/XDALFsuQEyaxrT8hex/PS2xlm1tC
NWqwCpyv0T5pc62TRH9i66rR0TiYDwTZynhTK720cO42UmuxaUvZHlwF8MYo0mM4lJBInYC2+Jp5
7fJPAkbR4KU8ZaAVJx7kT6Jq3+k93uZnoXKe4f1eu07m9yQQ6YyOw/PqxATTQ5GGTe0O1WCLtwN0
My5YCa88HuufT/Hg+PlowS9GTgtt32zxAa6fC2Q1/INcCk1YNHbr7GrhOECJNkWElCR2O9AgIctX
ecx9s+v7dV77v4KeOxfMJansxIL3p2sqM6Gv55sgrfTLLMZKIC4XYvBy8KroEjtbNVfCS4JXcLEM
sTm0/mu4VH8pTyrUBXxTCy56HFaUTH6eC3jNM1kRzBYeivahaU5mCEG7WPGfWJGoJHwTj1/P6lOl
dZxe3qtOQciP8quZG7ba5SUOC9mkhoq9bLNiloz0/XX9t5VdmRka0aXKmDLX1F/2iXvCCr+h4EUP
e7erHnMeXboefrJKwcUnKBWCPh8m0a9MvJFitzYcT18ckFw5ILLMw1bvm5lOB7dsD4Pn4WTj1ubV
xUbmfOTJrkNN2/wbSoenncyNAX6nfUpiBjIEbg/WHYz4h5GyiHcA7bW3RwNAcSzBwCGaL8MVbCjY
6LrtoIrw2u1qbCWrwEBEVcuvGLFbbAyCI8EjUktY73ezcTt46Fs+gHuEc78Ji+FJ+j9QwqfVzD7C
gr+L2OohUB2PW8LaeJOtU5FCPvw+tEU4qFTvTQf0eYPoMQNGHTU1bTHq2653sZa5MFzrq93Md8K2
r/8gVI+MqlsetVeMgooxGk93X/kuQhLD61kbLf9HHYie9kQyA2n63SzsAWo/EhQgEYBgdbwICtOD
BaYVHq+XQtfV+YQF4Mm5SMADMa/zDkSsFNtCXMTY5XJyIFpymp7CX9ofYetQrGtaRfZtm2TkFX9y
yyXxsAs6stfs2lNmabMRKPr3oBTv+bf3C7FEJ9KaJO85uRSynlyjyklcdKFmDy6eoGEtLO18Jjs3
uzE6ihZSD5ib/yEEPudgOted04DKyXU7E0PUP3wWQjSFxpjGqkAOYQQPwzTZDW/SZrIYKKby8HzV
xcdlM8YhfWIlj3TnW3BNVxdpgPlISZs4Wd80YykS4iAIBCFQdaFN2WVmWuuQ00Smt/P3L1RzPMEM
LVdYcvCxcKcRtQ7Ycea5PRYFxLM2sf7zEKm7JjEXkLjONAH0owoZ7axo0JPwa5kmJicwZ3l8ttXr
Pkdvt19yg46BYVOwJfHMQMOVblRUuwanaISJf4TYl8GTcEwK4Nj7JFEuVeHuXAgLMqPzxoUBlEWe
FcZuGeuGrvsNhIvVndXIPQcuhYtH6Qu5OhUwqKBqbjnY9XYCe28/EJ3s4gguY6ceHpmCbXiOk1FT
OQ+NL3KoFUE+uHihYGm6bwzL/MfN22ZNf1na7HtMtV++cuh5QKbwVKirKue7mA4M23f10OS7RZNK
kKHOfdUOePALokcIy0NPdy3IsvpQfzUHOCBEIIQsKoZmaC7ARutj8JqZJx9xniBwn+dAyCTp/I30
AkpKenP55QXXX3vigNxauAUi85uR5ZoZF7p5H9OrY5YIxhtQarcNfUAkYCv4CkwnJ8QbcxyVZGQ9
bQtgylkM1+lm1e2lujNPI2tPPfgdGBu/5W0anC85bv6vEgILPvTeNLBR/9Kx2id9hboBJdBvvIj1
LyGG1933klZ5CrCDzqNdhNswmnA4NJ5wOivhHpZSbsAz+L+at5V1xgpMiYL0tQRPhvwTglEZPTOO
fFb0vdY+SJ4CsPmqQXL8jYy6UUUTOxfPGSXupP9kPtaD6EMdTveCVEMNs77lELnRwnxA6xwXLdPm
9EoebQsO3t9rqchNng7gDCXuZdpgFfTMgGTaXZ78paCgbSzcBoW+aUP5eKTLKCYZ4rsE4yw9Vx+k
5Vj2lMOenCmYYFijNEPy/cnj6tmUgWiWDSusUhvITx4DOsAYdsYNXPy3kk3fHHYO/FgcbMVdD59z
JcfYTI9ZGIpCRmt4laPlEqAE43iQfwjRo3pK35sGiSIxU/23s1wfAOStsCIz9Mh6i9WaLe9fyHP5
PbMsbEXflC7lRwnCEShtZzW0vKrUx1GdALiZeMp5+LLGfcHFAl/64kQ7ePQ96xq6Zxhk+AOb3O45
oBp8woM02f6pCU+rZkwgoDx5FSZLir8Wd3OV55XyPwsHXrt8oRe1ew7dL4wKoZFGPpO5HbKPEtw6
toMoAXeNSrOvnPxtJCIzwlF+xUz1fVNMG66+lpgS5ouyPK8CRApS66lYEueBTABaEiLUFTotPzK0
YIr4L6GPQezOYBI6Uin4ZENSjpgtSJC9B+NIyxj1WFDuz73VTRHhrQn0qvS27mKcOjC570YNMqBU
s798h3gEVI40UfqWE85x2ovEE0P0A5flZYllWqHr4TOlzNNK1Qu/blxpzRW0x77zoincgAiECiZV
I/DSwLp8OR8TQzftmE2J8XreXVjAhGjiZ4tvvrJfLQOs9cGiVib6ueljnhk3oRJga8DPSOJLflCM
/ts9Y4ndYhA52TZ/TI+welDTHkJHea/oPJ4y+iznuvPzIJHhhSAR2ldw2Uq9WTrW10hKy5CY09fa
GDXNSw7u68QYIGTMrKX2F7Rbv7XnWYDcmFnM2WapGAf5LDH8B6GxQBg3sNs6CM74zJWnLRpUgTBf
Y9YKUl4vC+C19lZd7rF6Ho62YQNzRjq71LaT4AejhbZCnglblYFmWp48EUd/KJbZ7OeRJTX2l6gG
gH8szl8zX3mPiQnqW5n5Km6uIbq/DfJ6QsymJA+VX9pW/yONm33EmdpXxMQE1O7YwlsSfGfTGVLS
3sQYkbpxxhYhUX809EOfmmLEyk44Q3Tn1fNReCUGyi1Ul/Qs1MyRkdkeDtAIiRqUIv3XeFHiUjbS
pHQpoaeWXPQsxduNuaojl3H1orUBoThlra/M3/T+TZuDDNO/GVkwT9ajdQExn8uxU7KgHSluIPam
C+JJb2K7IYkZvxaaveqj1mktZXHDUxRoW55p8/hriOEh0go4H8uMjumVUkWOnsk0d/7L84X3LkUq
98pqFnCakIg9ghfh+R6zGTQwrfkEoSyWASqJkHxyAHD0M5JUiRDka4AIvNmhJbTyjideONQqjOVC
eo1MIovGp60HXLsvNLi6rI3IL9MVy1ZVetK9dEnDROeANbB/mrS568BzjaD8HuG6l2IcAmz2g+bu
5/iUCoafzVMtgmuRkl7APQQl3WXs1xN4XqIp4JmgywIPSvs7cCPE4tGkjTThKPJQ+Fk2nkM9nEJf
eKNzltwjNFulN7SAWvoKtwh4j9iunU2UDrnps+4g5J9czT0m1MtPPS9GSOsh8ZcPmCLF15AvBqwB
TXPWWWYSpi4YMldioENYwvtL0fxUuvs4q0di3rTRi2T0VbFwFQORkoMpym8ddGsIPpWLaxPKo5WM
JxofEhaSXOaINAPn/tqhXTKtJwolaHX2iiymSjpivydzWIsMBAJMv8suGXJYP1PK69nEF7bIkKG5
5viPlpWbYRha3YsDojByRoVLvru+nq+CNSAa1w4fOP7RDYHsNV/fMdI6C2op7SHPdXcXiVrkt6AO
YYuJLNhdK4lH5u39MmxHuy4HaNDLin4iflN9IrK3PogaDb8PiwGGz+zEJGMWA1VoR3BHxHORsd87
ygIRWmCPtLomwX3Rw8nwZwhLgafkTte/Xf0Gpuxj3o+tS/pbVPqvghwLw3Q8t/Mh7cJUU0gantKK
hsAlB7Mthy0YfYDLR9serPMve0fkgqC/AjfINRC+XnVfJgAfN07E30JfRo4PRiCMBYcT2PPj1bd9
sj07b6HJ4AY+7tygjXO5HYU3dHir5gtgsX2gFT1ik5rO/EVnqOi4E1Oo7pETK/ZxcR7S+zyZnkRT
msm5CMqZxnhY2jEbwHiY0Iv1VtRun2GqM1FiBQYzB0GrKl70KERDsRGxseh+6RQzZcIRE0mo4T0L
hFItN66OW3Iw5KziJWR1fzcB3M3R4HedZrk9av6r3lKCGNffBa71xRr9MQqKaWrSvrTdPYnF+FPp
dou4leOB3DOmkaSroW267UkvqVJNn1Z/iLlMWzun2VX2JVZnly/jvlpwcQEmo6b/Zcj6MD72k+N9
kVhWTTw4M/cxe5LtKppJ/t2hOX+z7LAki6p4LLLGtCNaYi8mbj00muXDg5T/lbDn26NCiSn01xd3
ejNxhm9uWzxPVYZdOV7LEoIy2f5BchcDuu8/IRZ2NzdgxoV2zr/WiAAPwmaEWNclAyYGdetD5B8F
nBlrzFWaq7f1Bx0Rx5NFz8x9F9Y9eQf61Cpa8Q39NgC/oDuJuWHihrl5jfm0bZKvZvVUzTnZnmXs
WIvBmVDKHcNlVBp4M989QhC1OkytarG2dctjA+U/k3uA3p9RxV5TKeK6aTeWW6hG6okRKM1SARkH
tTvOe1HagJJonUOZJLHeFJrCsdRzJmX5u9vPJmk3Qm5MRhlUb5plc60N+ES45nQgO3zAb6LjVHKx
TRHgy1noKTKr96jCvkPsZ3pMu0n2uFZu71FIkkImKLfCm5eDV6bQhiMBBXguJPCwX4QHLtQwTgcp
7tYG3+jwVS9qzlCqdjyuOGcd9/ByaTf8FwD4DlMMyVRHaOjwrl8OJDfbvN583XE8xivzDbqKsV75
7aGO7iDkZS7UQc7J7vi1N53B5IEzV7uEWf1gZJ/VAorE659d29xzn7jJfjiYWUzXvWFarRnpXqlk
1NRBBoEpl/ytrTcv3AnkeZM8hduNHYW0c0M0ixPgEIZURhMiBU+wPIvQ2cfKFQ3KPZvkH+Pkf9yn
3iRsIm2vCrMvvy+ZkmGG50cYhUCLB8ylh4NvYA0gO+i8XvDZW5yh3WtNlbPGJXuAlmXxzTwFHJe9
O11pve//KUFOfUxIzzeq8Gb0OezxNPMWusQHZj8nhbUz0Ew+Iqy+Vr0xw0+JQY9cxhoZhCsxx5EG
9TUT25mbBn0fLz4d/yimAz+w288y3EV3c6bDcwge4qTEFnR2CaMpsEnyo7debgY9MmNIi6231j0Z
KvNk/hkuiib/fJMTq5kr2/hvkUeSh0AQ7bWODZ4noMljUr2scQgFPcJ6EK+JPXFz/sR+R7ipiYOi
3lvTeTJj12z7CrKOHQ+NrJj9L1swj95yL/GJzAS5OqTx1C+lWYkEMYfsr5AbeU+pBJU9vTRE7+sW
bvyXnqcmGiDz063xbBJmbb0fcVMALA1K9HCzJ8VvjNBm4A9rY5UlVxQM8SC8lmlhh+7OgY2Eul7J
3i++bS4Uy4PpHcYAS9RWp1UPkI8uwHdPExlMwvoa6g7UlvDlDud7C4wxCLgAj9lKJJ8aUKCuIfHM
jBRin1CLg2uLRUkRqdNiq4hsSj6eJDfn0mqIBj4ixi50njH4rdnMiLmDjdUwxbu9yB1cL47POIKJ
8S/zo8fDZY3Y3jcamKBx5btlypdxA2tcZeOfB7XgCz/2yKFQCNC970qE63s4i2382NINzKgiJSg4
2imGdbVh96AqW09iPpJS8rpA8bjNXaVrkU5eNCYDdevE6CRCjh6UiKhdcsFRpocmcAds1KRjRYb6
cdkzqJKJRJMe8VaKq73QCgbFDKFAcoPhfXSovPTD3gWHKL4QySnIXzxArQV9rw+yyb/3bmRzxldO
hfXzgbDOw4D+2rP0y42iuvtBjScLd7ueBtKEL+m8lGoHieuk2uH8jcImyJbtwGs4SdBsjzbauS15
zsahm/0gApjaEMvqzE/h3UH/3DyDg/zkQHQnXm8hq9eHYcHyRo1aEpc8ANEMsUOWsNSpJSDG04ng
b4VdWABwQX8KF8pKxCWNBb3F4u6LtGGxU9pP3MNJV1Nf6MRXKda4zCTT9D8Ex+Z4NVKMKFAGdFaF
e1CbDmZzTgpY+zAKVmNQa+/5bgh4MmATkqwq+QfSIKcCKveve5uf3qTRgQnlmK/uT8IuFl8rJioe
uj93SEZbpR1POvKRtIfN0DhIev2hLyLWtTC7Z/P3U6NSe28O2jIFasmN+eU11y2gBb8JkUMtXi3W
l85x9231NPU1FBVFxfk33Yhc9NfOeM2MCLkf3AvH4CqzyJvC3LYGGwZK/w6hcG1qx0YLaOtpdQZY
PyPoy9MqERdmfvy1Q904qW4ZO35Xbv0s75jwwmeCQGXjm7XY5AeNxGJKwvDZ/KTaQG5kRQK8p0js
EE5MyU2lpEfRNC/S/+8y3C321D1GsrL1tiiGFhlXBHLoH64I90vecyXyUwhQd3dJs18+0+hi2E+S
ObPr31G3YS975ViJbc8jw++s3odOxqdFYxmRBA/R6Mi8QxZzwWtxFpETycr1HZcwDugdbQiv2x16
zTEscMUzE1VCb1yYUAQMrDqpTIJT52DUS/OvQOz7E9wrGusit6Seo/EUsTi+UzhEotQO0E8bpdCG
b/qu+tTJ64Mkwga8rPTNEWQEVOoYXCBUCJdk7zvwAF89HozV4S/vOsiFuxmmrzAkny/WDD4mcgFj
DrS947l2QmMN13mm+B+Q9Lguex6B859yeXRDlhVoHKhZfDAcfPlvqOzG5O0Di18iRkPlE7vX8Pq3
WNb4xXpoy9aZ54Nbjqrzbi00UzalfsA5XZyA6anR+ac7vJgGZHxYK1jWedepdHBwRQBAMk7XUh5Y
uwcb6efc29jssckbgBivzrznDCj1XnAdGRv8c41QHOErvkMTHZuNpSJ6r48re/fuZwAMuipPFzee
gs9k4JeHFssAcw4HwVlW4wOetpFCfekIMOMdIDy6k2zv8q0Emd/KQhbXEa1he5czjuCYQ8NJSQuJ
fxWLv1F7+g6JEB9NgVfAGSAQRbGpYl+SejN54qNpAdOGpeUNmmta89iO0MKhoAAlFT0Kcry52mzO
jd+KRK2/uX9r7vXlqRcXQpxiMITFlz+UZFC4LEJIZyyGXTKNXJPyUDCJoq48WOTP2zynvYkmp9gl
uHk9BhBFumr/oSTOo7xY5I0rvell1N4+EaD5iyQFZrt39JK+yAF9SWEyi6QPpLHf1P+PFciGBJX9
X3K04ZiuGk3Uk7PSxAQ4hoCpNWDk2xesTJIahKVL3S7hIlY1MnOZ+VLyjOPFJyielB3vhVF6pymK
md9hp5YZKAd6gL97zh8BtzCl+4tdN3DPXjRgDRG7SF8agAHP0wobzCr/HRgKv8OkFakkGnTLy024
Ms8Z8nlUhw4CQQFrPlmxAFEtfJ2MJFLGoR2cRZ3owllHaGBLU/rgC6jY7KU6mG0qHC9ieAO0Q1or
0EsahWi7MCPpgcW4vXE3oZfyUwTMAgXBdGjxroI8PRjvkwKvYi6QgTvUujONP7D6DYyPgDbsL63q
O/8aSy6INqt7o+omlSiaj6GYI70alhBw0TYjps7mNdlAMt0PfNx5GPcYfVmjKADFYIrbHUbvyJsV
5gFWhFA6UgNS8/A4P2nQTpDOY8O/pdvwEuzyBvRhec9lrOSiLMySIDaG+vZY4cjuijDgtexxCU2z
uwxSPTIr+SxtKweoAoAXPuGr6/55/ia5blzDSCuibPbXuuhZ87RQAXygBw17AC71lFkqqBAzT5Xr
Ysd+ldpocdW9/+ZHyv79lPAg6WNgcPAxgudwsE0okuoBjvspEYn4N7KyPI45p8mdy/1UMBbbIZsS
oPay64IqCFxzCpGBw7+fsvLm3vg/CfarV4bZ6XsZY2mK9b1WNZKxDl3dhm7kN2gUD5pu4RQvqiIM
f4TFnGMJ7qKjfm+72eINQEPmhMjrO50BogYUSyRO9Mj2Z9Xg+WUimZyA9Z9+2MFZjohmHzu5chjt
cOP0s0UyDcm4MkilJH23LyxwVQfeheAjJZ/ooTC/Rf01uyuD/RH8AfM0kNEJEHfIQBKg9At0wAyU
GgtUus2xjToB9bWGEk10Fzt3k9NSlcnNWpb9TieMGMDCJ10ZUPTsMRCiN10Veut9Dv6ypd4LPvLd
pdTNVOJGJUdg4GQ1HUEMiO3l6Ox+n87IxFlNhXVhU2zWbTpEGgDkuLClcGEbGhHtjrv5M902U+Ce
OEKL59jsoj9r2lU92apnfB5C55ExUlehw8CT4efqO5lEkV0iV+l07lrLnFNoJAPbxCzbJa6nx6Nv
FIusB7xjcymlBGKDjA3HMn5KdCXUaFN0+rrir0w0jcEktzwg1hFXD0tUh/OjjVOA6naHwUIhzBHp
10b6T58Ebs41yUWl0BCA3ZZH5P+v9XNT+6xWEi1+uqOBn+9TNSLcMPExltgrfz+BbV+fil8pYZBe
hkuBVaVd1B0M2iqjl4PnBtsFUQXjAloyaoav/sNVV6ovBW5NOICVhPGZJBkiCIqNhmoVlIzmnzCu
f3USO2kcJhDmwV4zVw97g4tIj4iE1zVKfd4tZr0JWQcHjNINsRUFuKzU3CqK6X+ke9BRWYbFoZDI
zCmkagpATf0kbnzyml+QeAHVIiaMQ4jHTHyiJ4VmuC79dSUOjU6/q/A9orszpkhvyH+pZMNTZSMp
rK4Px1i/IENo+Fmv1lcRaJ4vIk/MLqIdfQbGZfKvYRwOZL+Nksv6lPnlFNbXv6M6k6ml3FqWoq1j
hkfietVTOCBI2ABV2c2vYiOTpJCb9Du+p0yqlAydFMLDGbqkO9j79dKU+8xDKGXRH77hpt3Y6b0S
4ug+gz1kE6EzaJ1nX/kwKnoScGvMYB+LnXJRiAxVvO21h4K3bywWd2/wwIWgop8EFEckVrUEuex5
loQuO8ujJe092RoOHIg0xznx089GJ26kutmUdVEMzy+EKb6SN67AkiWxCmurqh4UE+N6S6fwq5do
cz+XTefke1A/GG8mQ17x8VOLAJdFNBUAuizjiQTo0FBPfdlrg9C47yoQRSFP6cvOECFl9MEzK5Dw
zEoCccGVJdQlcTp5FWf4/BlbE8rHQLNugA9aF1M3ptQ00sKUzJebYGxiVbIy+Tbn9ybfUQlXJRBr
Z7qgXP9jLJliPCcUuGQ+IQ04h0RQqA3FLioV+rQAejhUzr0EJNRz7jvuh5WH+ah18c2slPmZ2Uza
4jKRuaV3E7sQzQHr7epcHO7Tp5I61cbfFmMuJ9W+hXU/JSnOS5USxEfVjlvBpNprcvIETxV+3Bjx
aULOJaU15Rg7Lk0A6H2tdK9bZzSLpfTaNzVNa2yxGuRPCFThG8cKD+r8yLyl73br7ltR5LeDvoRJ
etmUTpxBt1JKxOBmg3jOq5mhVMkLmOOjGRidDSN6j/3Gzq0D/KYPE/Xr1c4Bz6QinDfV+uLjLySQ
fRJD6ayPk5bFd9khaFYyHocWySGhNDobXy/27a1VmHMHOWd6TXwfuUBo6Wt3+UPrS9au7NgFeZ1X
zl1fehhxXJrhKSCCoaOenKJ0mb/xw4fcp/lCbxj7Trpk5woUgC3Z/Dbs8PAGFtse82IUL6lFHI7x
HJolev+oKFCzIY8O+/4xx6tjjhhU8kyRjSHllZoPsEQ/s/nVITKNm1ScNqvWhvJHWUUJiBYaF0IJ
lyLlW8S45URiFDOeSBveN0yyOBV2xqxPqhNIOhy8btk8TA414PdaXzgoRZyPpUqUcTnjd5XeN+Ck
OEia6ESpsrAGdk2n3p4jwMilM//oX0xsOHdblMP2NQv5remTE2+nrYLnFRrsgVSXlaHfbAv6gzu7
j2TaPbsmx3Q5aU1fcZs9P0PXjxqwaepc4oUCTiiva+FKCxYlsDOuWivqMLyxEr+6bb2KbfjOWoah
/faC+PJ5YcTWCNmMAgjR/1t2tTuqsbM8P+4hmlS65IKAxEgMR+mTJ0uDziqkfk0qOUrsTHXUMi8J
a1tVIolwHsv++Q2k44+31LzYFss3hHe3gErxXSkUslZa5zPB+KAadnWowvhN3Jk4hvFZPdYv5axK
5vKAn5yXDFChzIl1Y00hciiwmRrWA1rpKmFVjQtvoAm7dw90Tdqj5js265Cozo2Re+RaaVAXnt2t
x8kWCqNBPKNRVuuLf4jyJ7XSk6sQBAyeoBM1MyisPsMB0Gm6bLR3uCfwY53FZhiSZeG212MwJ4jk
VybyRK9B+O5a+l2XfSK6grhA7HNSi2juHDZvnvQsrM4X+MFtnuAzFN99+yjxiECHm+CNZeDWyj4=
`pragma protect end_protected
