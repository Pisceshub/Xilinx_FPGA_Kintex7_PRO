`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7440)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEJHsVDFxnvZhMRBzEZudoRsXMKxpBbwEb7RyQmU0woPH5UmM6grfa9UO
DIv7sl55VCEbVesDazf0epftWTNxJoXYO57S406rxAFPttEBkRJLq9ZdabsR7DDC8al2T5q6TxTO
DHR7gsPax93Ia6nR79yia/AvVFU+NF4B1CfLBsRUTiJl1hbJGElzxb3HQljQjPUXCcKxpoMz0fuw
PtPzPArBE3bB4PHjTjo6zHaTPVJpLWs9OMgeQb0t2s8htgHMZLckrFZ3EX/ssR/JlxuiFoqfYgRk
X5QJJqsrmwPwBThBVRSScNvSMVXSn4YdEXwyKHdySA9c+CQ3FjqvHMf9AXcV5JXlZpMJDa4rUX8U
YKrWlLZmXTyMvtKlw/qYDwpW++az9WX2sN8sr/B0edvCU/0wNsTxK+z7wgaT2W9rH7tGT3aW8mYZ
AAuSUi+o0ccjBFnpsgkXmuea6/6Lp8dc4oWgJjwDyxWTix1uRRjD7fZZ9Q+C56gx96kP+StNBQq1
o4uZ83gxUgaig1kv3FfL82ofJcoYZ0ORox1kENUz+t3a15DSuEALWgmmykO8xAHrgaKLPsKFIUzx
I2ccuL0rln8tTNxBX52czD3NartBXvIn4ALeV6ZgCfQCOp2q3j5OGz80tsZqf15vS4Kka0QUMq9Y
QXDsom7lJ7sLpM04GxaxeXi9gGSk/iSIrGAy8EGXS/N2q765EWV5VoQ4ohLjC8yJrSc71WJOH8mO
YRVUveDtUxTnMPKEz3XwD45OAa2sXUr43SBHD8GHuPxdCL9x/kHkAOX96Uq2lrwxPDnetK+TuvJe
46QhlGt1+5gidcmHfAKX4YIxeCgIpXkflykeVuYd2ZsoOpFm2bxdHzdx4n7q2wMpF1L9HnOp1CyO
nK4QNCTsm8RLKgZMb/G1MZJktLKPDcdRGPKwkyHRBjAZ25S36lbAPiPCGS9JicGFZVMPVLzR/F/j
kLc/gzfGxrvbYz7qpcUvV2tomVqI+C4NrAnoRjZGvpq6k16lKL57JcgC1eQhzDtBm4evQG6mtUGV
cS2zRMPdac/SoI5thuO+uQnCooXMyKiTJqarJ8gnf5TX5rk7P7LiPiq9PR6jUDgHv508lYC/VyeD
nrCLBLJjmUqj0h2lEjid+xM3jteMUU+yLlfOF81BucO+x450qcOxTvqrv/LhX43J2SF1FaWvdN/A
GpxF5qxintsiyGBm/D6jUA4DaquKCZkW7G7jfVa6yLK8NasM5EAe4We6pY8uS2LKwSDs/ut/WEFM
Y5131F8Su8LiAHJWyLLvfXprFR8/p4eRGheqH7pzmLBSr7YYSN7QT8U7tsmaSNiDa5DKSG6PLKPG
O68yACz/EvhnSgCzmTAoTvSwhm/SsryHUrFP4cVen6vnuPtl6VqPsU9yW3CF3hBo6JfEhy5j3Tq7
xVBYxpdvDC1+lxwQ/Z5nD4ocLKoAtxGt2mnvnHjk8QMDX9kVq9Aht8sxe/QJOGk4e7ZQERYorRel
mPvN/H+8fDquKKTKxmfniiekDJu/IG/+40sOgvogNyWjoLoDHEtcw2+Z6Z/foZ+nWm8bA90CSdvj
p75pMwRrqcBb3K1IW5iaO5mHRh1r+7NlI6TOR+ZG2IAFUSHZeWbwYjit6Mdpo21O2xwvTDxUXqFJ
xJT9Eyj0eDrE7fRvfdwfIiZqarJ/hDcA2mldTsdlf/huCfu8tgblO2OjsJD5MK3F6SGV5zk8pu4t
xzFF0w7Mp3/DveoLoNesvrkYIcl4YCFdNBhqPBT1G6WyqaG8Dv3QjcjIM+P2crwdQFxze3VnimcP
SVnnGonvEgPLEEDSJBEb0JHHCnP8VQ6J6tKc+87J1d8FAXSWHyDjM0Q41qPjPEPeHxrSERnPBqDy
urGHkEUDBFVoxYkv26aUvYy82xaCMMDJrpdszdB/WraDgcRhNQoE4Xjk1F/jX/mQqEKUUiaak8Xd
ckhkA9GO+RYNYcAb6/8pQXsamRB4VQ5BCPzeoLrRhzxjIVTpDCt333nO4sMQvHV/QsjdjbfusAy8
f6wgv/UZMqq8ZPkRV2ytFcrM4AHXfvhv5LGT1WRduPK41u4O+cLcYtjLS8C0GFW56QY10AEYSMBm
OM+6bGJH/lcKIzyUBJWIoMrgIrIRH9MTMHkp4WtXy5JFNeFKf5g2rtZqLaOerBDBIFETqVXMBqdr
VYiIrs/jeV9N40jamhIri/yrrXNEm1VcJjtuszfIB+dMYHYXKBpFqQvORmosLIvNP70VCzTKXN0W
nEmFpj5LV9oeR1BVwVzs7t7LZOXfav2Gmfb2LRH1l3L2MLZILUASgdFqDL/tuSSgHp84OwfFir0L
73axL+rxT2UC1WMqd+XYdrkFK6dND+X4N56FKlbDoCoTt+zrtWRZrz634BYpqN1/RIpC+1PWGvgJ
jpLR9BHe2WzjA0TM3QWAwV28Kq0LET6mO+ZVn1w+ZJXXcyi6yai79df+H9ItYbGa+55c9A8lyBHM
ojxo6V/E19GcbXF6yWetUVyvzOVQydxfBT6+UsOzR85Vpojn47Houa2V39eSis4cXMu88BH1LSol
fP8TB+Xgju7NM7lSuq99wfYoDaG9I4IRoxDHJM7UAToGoIu4hap7K7So2PbH2mxPsWSykUKONMwS
79If86w4niUTnLBTAWpytS8zRuIlQHCtNqfrSpfSIbAwk+2svkWEL7S7t+2re6KFZDHHkMkCLOMG
05uDMl5zo4ow7D/sakmCAc0T5qn9QLnjTYlA4Ve3UmIOojRww7FxBUQs8Gobw9IwkNNpDlf3fy+i
Wvnnuask8gxRnDMAQhChJw5+XS/N644k5WKUUH5Cp+wjO9S3LnyY73KVGfZ8Pu3p0WSHQ3lzE5C3
MXjOyfeQDI5DimIrKzOO17uo2JIHoMI9qxpIKZ7PFHkrtH1fdnfux0KxGaeh+LLqFguCBul4APJN
uin0Ik/imWIQ5Z1Upz/ouKr9pZ90Kt0qG6+vXkdTVrlPQCLMDD/WWGpmnZsOPStUoqekokaBmlu0
fIM470fQA7FqExPwrX/o9myOPrMwJP1qbrpCyji0zLZO00Ve950rZDAuMdlKrAbnK8Ka0Ust6T1G
LNYhkNajM6O1l3o02DvLuFpV5atyggaEOON4ESKGkHhlEa/fDhbPRc1uWYyTjgNdjZfs95I7i8Tb
gf4q1OTGgn06wn3i7BLG+IUBEbVtyX8PIAh7XEcFvVPMdhj+cvbMaaGmv4v5PQc9h21o71pal70N
nj4w46sLeiZgBZl/Z4ZkL0K55n9s4WTFiqIPZPzuqlv/SmPddsacV+MGyLj8RhFJcas/G/wb4sDZ
WX5dRkyfNMdSVRfWrABDPA3RmkaFuRN0xC/o8Y2K7GaMW6hjHCvuMMPJ39zFUPwUcRLdIgcZIfx7
CuxqG1YgJ6NuyYcMcoo3W8y5RCzKzmgeOzn2LdMDDKe1mfuAaluptq0krv1gdOxBdphUbmiUhOTD
B4pRIxItR7rb8AkGl+gd2KWgJ4dx4k9Id5283Ww4HWXKA5g3QOXlUT1eEtLkHYGAXQzOwj+ULv1+
2Q6ewIG6R2Z77tHly8Iv8ncVJzqtgN+eTr9yyRNDqqZsOZu3+bBNLTmugljM/qpNaDBI8UzaVuyt
v8CXzSNx9r6vS9j5k2qy/UT36uGnJvl7KvXh3d91SVOjO1QQn2eov4Tu+YriWGexFdR+4d+rqgB5
fQ6SKzs1cBk5RiIS45uGqruqiPkvrMBmgwFXPit6TH2zP8vriGoVK3fuIT4O5eUvCrBKwwziFdyq
LxhZCe0mYgdkGcR9h4ZVAU6etl+0Y6VeEE+xjarG6eyJpgnRZZTD3DOl0Ha4ozMFowysEOzs9Pqq
aGxTu8+L82fOA/U2FZWyQYLaT9u4EMo/Uzi1BfiXSure7UGyXqGydSRYD2mvUIQ7z/LnY4R/MJFn
yugT+5bWv7U0KGlhz5SqMow2xEZ16pCmlVMaFEk5rPWQQmBeCj3k2YCDK2+SR6ffdHONX3NFFGgh
Kc3LW6BLj63Wq+NATb5bPhypUYI5JMfknDJAhO9AffsGsMXbEmExusypgTk+wcW9Rv3JHgAcxXkh
cbhYzZ8UzWiiGW5dPT2dhy7MKGs4mS57YaI/wOq+/YQLJEHNFkOXVl5S5nPfQgDO08QIIJiNZAI0
JekFFZxWmUxRXLU85oBb7sMMyfs1dZAqvtmOwnO5m5B2MXcd72/wtvrI9Or12/DmvhYuiT5qjLUi
PvALLEIITibc9GCzm3HVFv+MdEH1juf0jU7XegXUVMrRs9D0lx2hcmWFm1kO8evRX5+ccy4yxtCx
lInkvYBnblUlm8IWLU9cA4KDNLXbTv7KnN94m2k9cGLvA6zv4aOt1qnSW8OvcCzBHfNTSzpcvDnb
96O96krU5tM1jQQp68Iq+HSov4quKS6DdUWdIM5Q0V6BPFwokBApX39nPN4s5rT19oxQhSiu+f6E
D7d/yXmjWs6TCU/5VF3TAW1tVxWtEF6GTyJWWS4KxTkGuQv21TF80GAUSJcVQ2XeS1GdDtQkfOYA
dmXjtRNg7h5m6WyVwLvp+Pu3DuL4md1OC4dl8ZWJ4DyaolyRs00BFkyrWysGcTs/m6Sp/an0wdGM
nyy5YSEn7cw1VgLvBDohZM/+nxypyCC2avv6VSHzeEXuI5PZnzKDhcc7FtXOCUOkKa9NEdlmlEVc
sQUsyrKc1vW2VMJMvG9c9aWV3jnpQmk4uxjJSXLN69FKTucufy85bFTeeYVUA3U8egCX1Vm34HtB
jpxExGGVuhw7VTP0aEHWPwRGl+QcXjeIyQlo2XAqarKLN51p3dKzMCHabeWaVg4rqk3B7h+ekB+h
6fsxm4JGhly98sEpNpK318XIKP8jvizFZJNR0f1TgMGfAaj9mcQqCEs72ySc9StI7eo3fn/X0Go3
CTBtCRYC2OCwbxxyREfjT1VX/3kAVqGvPbr0sBjsfHTHDaSBlrdCWxF5zuHYxQfoCkMrsjD8vUf5
cd/K/SZj2sofN6N+TrI9DWiwdqe/RzyDAXQ4RqIjlV0eay1LDG+316m/luIzv1d0YqAxgJyYV8Jf
D8Pj2H3IlfUIBJjMswwM+hXpzAvIsWcKKclwRDwy3Sns+vuK4iRIdiYBhd3gcte+XL/p3/w9+a9+
MuXiuXwk2K4QBFpFB/pGM9kXfyf9NvAS1RpmX4FcQ3TVAh5ZbeVVyyd3hdTGqdkHR2NKSHYfPJuF
QGx0GszMXMaSsrf0yttp/iUuXVur5hJ1LTEj6fbyoFV26A++AvNlZOryh7TVHMoiRyqW1dHolS97
mwa+cIZ1Wc2Wi6Jurp6uEj5rTgMnYAVOMsQrSDWSFpcxpsGOeAtVSCvC1fP1wQ3CgdQT1SHUMedU
bJjSqM32j2tkecsyU1uIV34OtZpgFwtdi7O/iZU9zIf3EFGv/1bxCzIt39gevygMhkE0ZmBkj3Nd
Iayv2bJRveMM3BTG359uKOu0BUUTlicoD1ew/UV9tg2wR90YbapmRcI1Li7jVfw0IkObE9f7EwNJ
FwkOytcXkJj+toS9NgHovP8EjfUlefTWgA+Lfyk5mEazT158vJj7jgTQO3V19IoolkGzazDbZ10n
VnSm4MKY3oDt1IrqZVQy3gtSwOlqg+Oi61+EED6+Wycf/jXgNw3634NaKHWtV64lJ7mlj3ydo0/H
2SC1LP3JvflYN2aIt6HUzFd3nwTlU1m5kXkWy1Q+5KaJiFdztNVntLRqaA+PnXYCx8bVJkNgifmH
znPEtko6rF9i1EO9/3iq/fudwvehCB55Ew5+LSe9356SIYLySL7M5nT0r6CVTz1k8Nfkdi45t33y
oh5/i9X8TwxenySDEKBwiaPzQLwONCCl1Fit0Pegmk21vdRpse+v5ETJBy8s6y0xcyYmrzdZ8kKg
FuZiO1DyuVzrSCKSshZQSbgdRoS46gTd2HIBaol2gV7YpOfxoKskZUN0Pv8W3rW7CNS0yop+VkWC
fsRJDZYsQ9B+Fz2wCwyrWquiwbCxpc2A4pWnAdUZ/zPUSQ5xzpGSuiu01nUjQ9AmHoPgut/+6Zaq
6dIXUkeyNCmShA7CymNuuYgYPenGTGnDz1y0khIbjPqG+XRneFV2Q+T4KXWVytxTJMQJR4kp0rQh
qSdEc9L+mVx7CMy9HFMYmAZ5ZR0gekaZpmrFGvQ3W6DG6U1CnFDrsAPjscidWGquHW/PJPF7ANxS
XqY/tnMti5d7j5G/NVDgNfLV9VkMIxC0uG1Bccpptn+XSY86TghiyW4IsKua+ZS5XiXTWkrsXAGC
fARZIFytiXnLZaH+0Fb/idSEdB2ESFQg6/PwU3kOcb3cCWsa7I8McL8g//va6h1aEK0r/VdKO/Rj
trTPyYztuns5Puc6QyahgAhgUJIrmvk4ioe0U/5+OYhPtwnakmJidkS+8RGj6g9W1Q9GNeQTa1dP
9M+CBlzCFuhS8nyFDCOAXEqvwRhDEh3YVaKvRxapaS79hPmaOHtma/4WFtTqs+2nT7CmGjE8PVe1
01Ly9O/B6llE+DkKZBKR7n6hS6faN8epJAkA+k549JGhMGVezMcCM0SMYk1uLaaI71iuElkvd+4n
qZPWO9pAvrBSdiSYTLhrZEcxLbs1yVHtPadpO1ZIKFaW5ywb3bEc5tKF5882TaMH+7JhkqYgboIk
JMUg8bVoLPf4w49BN8E0UZlsek4W2crQLuCKlj9mjFlhWjfmpqV16q/yRA4wtP+t3PQ/T01wyAHC
EAm6EU+EKEFcAkS6+aAAa6YqH0DTHJ2C29VDXXKX59Ac8OTBxrcoIqq48gcbukV1YHMxTqj4BOKV
8rfs5FjVC/mGlqpv4S0zpzFVxq+lIYaw0JBIBJOJ3r9OaO3RT+WolwotlwYyHCIRlYKgu+uzox6B
4XINN6GfegyNvzvxWyVkagRh7zWL+uvHnThwSvPCRm+qMH8NwJ9X8mIvioPD7x5l6tdE8cQp7Zzr
/gr4UZRCY17mfWbFTERW9L7PjF6lefzaba6/qdOj4UlPWKIyYakTfx9eXtUT14HDT0CuhvTnpUfh
s7V184p2HZDMNmGBD6x24GoTNTk6XO/JF6a8sUTCMYK6Rz0nDza90DQgaLItTHIiAhISoDpC0ji0
lyF0rKJmO6pejoQ5JH77NWFGot+FiI/7uTEFiLrUXm49UAi+P/oWT4P/5NwtAhuXjTIHT+P4fqXl
Tq9lyIMOIE6w9yDFVILn4hAXXrn77brpuJEjtdV8Pp/BdikXOfF39myT75MZGDoQDnPTOubinmvg
mjPd98LAMbB4Acgpziq2RG5QVCu/2yXzkf8qZZznVB3LDO8Pe10JJ/XExXeCY2al0gWVfJ683mga
R3PWbIrMsMHvNMT1ZRYec2TbjKiCTtWJLk28x/sweTYunYVibX2tTpO3gJ5lV/8hMLeI4ldgif3v
O4hi4aFMjrCrUsSbzyFCnVCLrlvF4bsr/YSIxSzujbHuzQrx94NC76bNqDxA4icIeD6cDpNoKG/a
VOS6A3XQJhuFLMba01p+ict+BRfaNH3OCeEup+P+00qxaYf5XMAwhMeiNGhQPGa8ZMtJG8BttkO3
blcrxd3D7IZkXaCU1ToMaYbjUDwpQUyTsvTqbLhz4pae+qZGqhvKXbrP4J7/m+AQU2VE7xIcHUb6
6v2hVSJvbBZJx0MOaF0GdaBUcsU0rsDz6uyRSw72PbnPkccw/Z1Oa6UwzMDuyGJpO/shTlRsWwHr
iDXRbTgMMnJKufoTWMeje7TD83EqQsQDELrw77/33rOufV80+kFmTRUUAHeHtvferbSuhfhXYv7T
13NnW+L71iobjnKo/VIR2f0zUbXnlf2d+MkprwjV+w1Wys6YStp5isqSo5LlKN3QURr3eOUHROJF
U+s5puYKWTFDWdfLVjODpRkQYdcnLxf4xqsgR+y6ZJJVNaGmrgEn4jiGe9ht4zutSN3LgpVXLhz6
mu3lYRvoi+TMKZW9+LZeUkfBuWLA1sMLc6JjNsusw6Esj843N9IXrbJmlMA3uNYzhaN2LFOU19jQ
xKBeGdxB6fXsxSLW/6a2ayQb0fOK/VqGKxk5Fc0MF5N5TWO1fnRE+qHD+FqssQZROQLNgakz3KA5
vTwq/lUol2Izj3vEpMLQ2thCp0tVPPRkSPDYzg2wIzNwTMGfIPH73Z9BNU6mDXiZ70QDXfKPFVym
CkqnbZnwpi6+U3uldDcYAvZxpqF1BcG6hIGN83SVVfm0oqbc1WLpWSdJW32/Heg9fZ73OItKFFhB
Mj+edwJ2glLOjhexu09T0RXDQaY/qabroILcGyCe39XI80106QstWZVX32wQR/9qaXf0RMZH1/+J
S1buzj2zFfciBCs7lURopajhxAcT/W4MFv8192eYaqA0yLbBX9A1LxE+1vsTF64L+/+8p77d8RAO
BE7izdzX/8dmYNBd7J/HMFhJLni7M6uamoo0lJgei7Uxc7/NTUjhlSguP/e21HWGX2LJ820vErCw
iGTbBITx6RXy+TdlK18qg9c6FFMKUg6VqTg5+4jMZA/3b9HwzPnDqmktJZylzy94pxFwE+O0dfoV
mbkGGq9YpedHVKiputMjM6+iVP7AsNb6wwz9Ne4ILeL2HUprzkaT8K5K1cNSmeopO6ZFdqjIe4H+
9+7KKlyJcFM7QBRvo0RcfEoyw0ahawW3x42G5CeN6UAcOn1p8mLdPTnzsJ8Sy7Ixk43uFYymtbQH
mc/2nnMX7eBdiR/tEjhzkSkTXPNskSViWpTRcpXs2r0cj1QQesW2SMZf7YfNkoVRleWlmkfczBF5
2a+8x5VBPzG3ZqGKfm0DDS4yZ38lh8wl3ENQODA0fBZ0aTLMwgk3n4r9QCii7bZvSKNsldCWsTx2
CG+y4J5Ta7a/1FFHg9NPjrY1lHCrS9nukF4O4kyoa2fW8pqTUiE3atDqfK2XJB5VZof0B4PjlotK
5J39/lqznQo//9+DCWBln5QoeajGYZggo8097hISsanAAZXLvH7xtqy2Z/k4Fa9S63Tu5YAGM72U
OCiSlqsI4zki6HtY9ylkysf6+0b11rjCigJ+daezyYgHMwiOHSp3wYDgFQQPVoIlet1RgPDvw33Z
SjJbrQKE48DH4BI8i/Lj1jx2fkk40kUSdXh+5Qs8hBbMNUh/1Muz9CQuMSq67pdaZbtLpObDgECz
HjrdfLhQl5GrO0EQjGsmUUR/2e/fy8eI73GFZj7X/DqbZR+uFYZ0zCOJ+fMXDh63he62tzTwtYeO
5C50FxQKCoS/16AbcKJZi1NuVp8snwITpolw+5Zj75g0Exxf/4UoyXIp2wXgSSY+VemV/2nmQQTE
/0uIic4EanNrW53vRH9pXwFHTo+ED4zWyl1JKll4sVtZjFgUWxmu9GLL6rmhwfVSiZWjGTpoFRib
oCWN9UhKgRJ9z3tJK5f8B6DasJdrjx32Kd9AXtoFWNmWjpvEATIeslCd1IhiNp2eo6b21EHJ5JUQ
VU/apUKjxi90Yr00XEmYY/KhXoz6XLhmNFrorF6LrvkWpSmtSQ5Fjk0yBKcTnMAs+rqkUJUKvMbb
BCAgvL2l3ZVD48CFve49kMZwZ1tZX1Mmdz+8brUUzETBmxG16Wptsi6d4EpUgMn1QoPBijVePrmf
PXGXglsrXWKD0F8g5eg+tTF2HByPKjjKb/RuKkveVu1k5ndEopC5qP5pMQynJFz7M01ZKWQKQhcW
iWrfO5R59sEcItFciC5fl6a5bgwE5dMv/L6w74CnLj3Xf94ppOKbjUOUGhamKSeJb8dcZExgYteD
r3+I31ZmYVPp/O7N1I38IGJgsvmZui0pusroTKeLWNJdI2n9RVBe4l0Es/nNYTxr0G7nbO3O+E5f
kWE/o9HQ6BV7RlzA2Q7+ryqxIJoWPsJBRbBdYEjT
`pragma protect end_protected
