`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
UVUeVClc20yTY4qDHWGpRdAGVs7hKwUNlvcKeV0hdPxORbQrQerFBArkgGE80cpuN0AvSOknvhu6
YkjHdIiO4g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oeTmEiQbM1ka7XzqgfHZgHkgAnj/QT82N8+aOVJRv2obDgfzYLphDpGsbZYrWZUjp57XPMd542/D
4HcWuMKjZ+NreUvtMCPBluoQ1tc4bO2STu1iNx8zY1wvQHzX1gX7044+mjAAs2w+sEd+Yi5bBhQ+
9zIJxVyU+T6sN5a8Omw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
vkLRS2RdQLKC8qx7iuv5W5AtAWoYm31sdgZOluKLHkLush/7fmf5ryaxgAV6hmJVUCnefRt7c3hr
Rx97eThNoLzSBq5R3bhmbnItoRbBG8FVF1XrG1qNfW7u2hEmzlkZlq4iElwLHOnZpuCkTu/hGvWC
T2smQs8oI/x8MWf8qXt6MEp2Kd1n3R0E/dvg/OFGTrFjBiLs64l+46SjGDqUPD4nDbFrO0XQVtnp
+5m68nox4e48I1B6knXudXCfQnpaHxtaxIifvzH5PIjB62j70EEIX9b+iOoKNAJuB++5zYU997tv
VSxbdJRv+l4S7bj6Q9vDGxF9lrCHdUvOztnyHw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
U5ba5VGWHfHdMv2tAQ7kikAnjXRhKGS/4bNO/Y2PJw3c5N9ujojv5im7jgcCXq0TonXPPWPJLJn/
7xu/PPpRz2O5SEIaPVETqhVUjc8F9HajgmbqurKULpWA15vskdmQYGt6owCpaJu6MPSxTMZYjwnx
uxGKTLbF86Eyd56tVyrkGpP/saGlwCceac426Lb+ugDxm5z90CChi1nzy4etFw9KZLcceFwvPQz9
58W8RZ30qqEoSMq6adyrvyT4+IvzXAUzQDv10KXKGqxinWdyBEegZ+J1SdpSnjX+Z4l8qZ5YFxxc
Fqy/LV94YZgmMgOoBjwquDxzkWyjoYAtJPKGtg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Rqv8Mn/4chYzqTTb8T2j3/MxI70dOtwbEHtKj5xS5glfAgFdhIi8ENexdFk8V2n50qdAi1jHh29n
+vlxhkqQ61GSO/56wavmByzZJE20BgS+TdFANFeYye4yrcXYSjp3abtZ5cz1LWVY9ytrbCqa2BzB
NBTDm2YwqkFm1CeWMVBRmRTeCFo4Kh5JOUgnHHziyxXpjJu8F7Q+dnW4aztMDBuKsiqEvpyvjjAz
AWrL559msVcP3ygsM8tlg95Tok0rJT2lsksN/+5TdEdZ+D2n7qZKnvxdpikOa9hF+o5eWaX7xeoR
+C5eID/gsNKWPEFGVCVPpqA96P6iWRlOYK6JTw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aTBPcOUzbRJfTcc26CKEu9GzKlGTHCrqUvnfH+MRnzp1xRnMuIfu6Ce8amP19T70eplvDyZ62Fsh
nlHvW/VePfNo2iYAHmIsExEpFqLqhM0bw9g6P3ucDISkLzHQ8a4MzqRGicVftoCciRgrBTiGG3Qa
18AyCnhVWUBWh5yxlxA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
LVk1pdVEPPmz/4wAV6yS6f6zgN36XphdMnOYLX1C99B7oBTeT4+BkY9hyZbxEdsHAtTu2pdmvUsQ
mWSNq98UogMWnGLqSCzU51tR1CFIr/hjlkJBaKYbbAzz6JBLBHZ7Jv7FsvrHqekqDPSoyihsR/vt
IPkjKTTQFEy/kHB2vM1xfp2nLFpgUn0XfUcXBOxKDfY7OTdB+sm0n5PFkt1uv4hmzNXi2kVmkyRT
C6mbrmORpRWip8ljD26vKsxjUMDLebbYzp/kfkIdz0TLqeNlF0LL5CkiXgtbl0TGe1zPLUbeyGa8
rRY+yPdr3rtb/mA5dJhprvl5zoPbn/Tq4MM3sw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 123984)
`pragma protect data_block
Z9GzGQTp8hLj9+qKGo5z9MVAJWDJHNzPOTKFbvhWRW1Wt7RepD1hSZa6PJsneFHAFx/n6opAiTNI
UHTBXvKJCnQC+LyqG4zd+FkRxd3GmJswYUYAMhGTQ32xlVP13NjDz25kIbzhfj86OAD3dN5UGJr8
4oF9XXu3hv5YNcz9YxWv1aLm0l3rAHiwRrmB3r8EU0NWpuFkBjesQVXtfJ0krkFMC4SRojiQDwkE
ot/yCublmSaX0QNU6h437d4nIDnBrki2DZys8dQGaf++L15nvE0KlI5PXx0TMKzo2DMlOAMGqCVF
ALeKIPlci1MvZqdXIdVN+SorWey3YIGAmBU41mcHlQMV6XSov1XT4g1Pos2uMVihqmFFaOI3c9VJ
mYWosWAldvzHshGyl1ruT31mbBIsDJVfu0CZxHVZBU3+I7deSX7UWPkwCopyqntUOVlS71EK+FEc
y0CY1nuaY3hG8JaJyJWkHgiqc+xUNBU9DeB5xuUgr0lbkWLD2YdnXwnrliVlStagAL7WMHnhKdc/
6wQVGwYnSxBZ9Ko8A7dCAEXGAvGPUVrMlwPRZz/mvnxXc+/G9hhNez8TPhd96BaZHWYNbbf0BvZi
wzZ0+DdhNaOoeNIsEeTn/aiaKhbHfIm6CfVVZEV8tUrMuTjNE4z+p/TkUYPL8llFalDRPGRfW7Vc
+jTvhwASSwlEHikSUICV539DfHNl9Zk5XDKEEFBgvo9+lZRgdfNl8WMYmrC2/IyU3PWHrKwDucDp
efG/UAq2IpAawVWi/vOm22BCRIs/JaUubZRxFRivKX2QadViyo7XQPOUMoD1KRaV2HZbpUcyIlmb
gbdV6G7XFrRuuuFZWIsHANVUFbGvJlnjlCYa3abGaDt63vsvjTSUgCS6+uzeS0+9faMPLJVqTkoE
YHJ7ndNTFK62tOv5Quv+QeoRj2uueg/k5p454f+qPEkH2qV0BE7hXkXz/3GDjRdun9q6pOOmmlfM
5m5RXWsaclVSxbFMUBJSJeOlVcBk4JVf+2chuL9dC7+qJH5QGemxIDVAQGBeXY8pC2x4MG5mw/BD
pp9W2YFfjVdI90FgPtVFsPWL2ZxC2/lpudAWcNciO1ovVRY47enL2uHyy6gYcfguitvcOBJAWoVo
C4fF2uejMlwjYqaeDKfaAveiBj0+5Vmb/6rJVuFuP0vCF8iYTZzFwIjllERvI5faL2TYRAZkz6vw
lmeIyvLpLdv++Cxj6LjQ5aN3a1QH2+ef6U1zO8Y/q0BvdcR2xsPSSFJ+gTPX65rifzDRlWzP1hs8
L9acnQ3GN25pdtsgnpI6bSU7fgyCmisSbl+Pk3joRqp9vvHbbBrqG+iSgZWpzgKMgMHx5e0c0b8Y
aaPQ7dnfy70ZyeC5OYTe/mQ0UC3WhGuiKx9Fvg3apUx4fbykODRImqsydYXdlk3/0EX5WGhPJdpl
/qwsSAcyxI95LB6RcvzPdt0SqngKsrqmTt3jvu4TI0C3qeZ3nD8nzs4+D/55P/oV2/QRInVe1HPz
ScyZaM5Ul9NpTD4zN/lmh0Ses9Octb0ahFqFUv6IkeMHhIsROnaj1KkTslBXEpHuAikghYkdBeoG
Ze2wAxJboHUf1Kj9Jpf5z3D+5vt8LrHrAZU8qZXRgzcZqqHQsYk9yEnKkD3ZK90nPIe4f6qPWFsi
YHBgEDEBYsnjqlyEKaBLDAjr5rROe2odzEazbhMsEUzso+0BeoZNd+XYuwWgCv95DwN/n8MEEsYI
mJUUag+akwySNOyRH1wNUCo8JuRRXB6iIU1m8hHVnk1BLCjKEul1TE7ViXpsj76zfnp5EWSXZ2nu
JawwNy+tq54HWIalrvMhiVeA6rajc8QmpNUeLq3nP1LSgPTelGQ4j87H8l5QrbEdIHpUCGpsaKO/
rwEDGSjJc/lVzK7x+Yw8WH/7LbTRjUHrKI3vA497TOgYoYmibfwYv6FiFaA5KOGfNI2TiATgU/dW
h4/XvxVvOwI2u4h6xHGAGi/fJA5JKIPToo2PdRYeyNDJaV3PXP5WUpr2WngHI517NkGq5mX6lR8t
CD5iJ8qq7FDM7iXJ4nU8K3XKfGYND8t/rdCj3EDykSQsiD0/L/IQHr/FBZA274xxadmSnGi80AC9
M0JRZ/griH025Y4G46wE18HWXRCdni6RJYrriiymvGFDSwF8D5ZAcJgPtSfJyfSfT5WLPa7pXc9G
NGwf+CE6dcsBfus5qebouGifODoUI5Q74IVOQZgg+WTQD76P+QZxu1mINwRNQS3GO9X4V2E237qL
z9X2wCDEfjS2OpslHL37DClzxU7HoWH8mnQPrS2AGAug5tGmVek1Sv2ZPkiy1fs85sLUmCblQFFQ
wYocys57LgAc6CdXIUcKmaBt/QrMOaKDktgk+p0eQg1haMKdDI232icbQ0zqgw3PcRNBhHg2xeeb
udZLIHcieg2CPgxMwuWVmKQhpIwmu+sZWTKDtas1wflBq8k5/4mrNTrnggOI6DQY0S7uycNpnNKX
UvMelaOW4g4dIakXE/FXKO2VccZxWSXplnlQGRqHF2dyH5GpoOOqbrOJCHD5L0uehh5uNRSx1GlC
+UJLLcMTX14ytmx0xechtGjFbvu0yVg+D8wR6GFPw587sYBQpv0FcIewEOvMmHxrGBwbRefurzqS
GNicjLtLZeB/VPL6w8sTkfkK25hGj/uxwRddGksC1lP+3Vz/7vLl1CEqgiWSTUInIOkt+FBZVGYH
jWJ+HGYcmhKsiD6PO/HYEvx/d7djGBcWhLEL38BSjSNwGatsdlRWXIrKsbg09F86L6NZdFJiZl91
himk+xm9wjUj+aFBniol4dmXghioC4i9ymFUtXmiA51iS4+lewke7B8RwWPPHaQj63luq6DvpDlp
VSu719bIy7rJXGLPTeWJuxVhh9Sg3NRnjHdoqoyYoFESarh12NBmHdeqr2uwbDltjGiDXuerF4Ix
9l+wqJlQTt+cbTjBeEbizn6ercMJSzVaO13mTOccInW4G1D7ApYvwe/Iefn+PvsMF0/+mjWjPS2H
pXYaZDtjwITZuCkx0Rp8A6jbU2Wwj0aHxEgAhPf0+bJ8ym7oQWoS634qyKLyrnucZsS8+iz1BjE5
xEr3v/9b5YK8alwZSv/7Alkrt2acIXK5T5khTIoWtF4fJFKyw8mMgM93mjg9vgqPhnekctEPMOAi
aS2ZkGEWyyUzLnsZUJSCxXPTpgqdPWmjtGr1a73sZlHLM804rDmGoNCwe2eUbYrI4NAbi20xaGN0
ch+fwjF5Cl5nze6DpWWn4j4SgC+uEOpeuGpYfKoTe52GayGjM5rBG9DC2wBGQHYqK8oOXEBTTxu4
lw1NB1h2PTlla1i0kAfij0yhzIPUviTHxLyPmwjfWjwLYSMn3v4FaERxU0z2EFdVTT1P+HqYh1uc
pMu7pmDKqqdgkygPo/s+LZtwlgITsmjTnkN57Fa6qevdHqbTovWqo4oUGN8tz8KimdwzXGzjjD+3
iYGSY8zlBAGxQ/oX5OznMN5xoxgTdQ2dK9IoKCQ4/c9osFRIc7Ll+Y9RExW0n1ATxvrdjok1N76r
mED5985F8+0Ik9Q0Sg2jQ/wN+My7fXPhk5lusdXegYZYCNRQ4L5swc4dYxpF701GFk/NDbgvMx0I
XrkGQ9sreWQplAoskAvblqUBxgVj6KuCnqgUwwYwExIV7Ip3df4fuVWzvhuFuKZhKq1GvHM9BvSx
YruXnb3hWK2jrkaaTxJ8JjdJXQZtckN6MV2yg6C6G87vA0AX0hiMOLgUMu2no3bvstMFf+UcIUXk
++1qrFYQOVZNEpCaFtrXyW80C3zzqsNWJO1olf27VRqhNOPqO01tSwk2hFxu6+tmJodmH0Q+f4Og
BqPB5H7+CyIrg/uqCD7fOvVyJkNT+j+/o2S7xbPRiDLG4jITYReUPpdKH2Bfn5mcN/n0qXxghHn0
P7HUUhXZFx0AJGEb21mOJi+l3IBsbPq7VyouVVAwjbW2Wxq1r3CzIn/84HRenRnAEb/bD5gw/sCJ
96x1qxVDHP0D75sHLJiW1cdZHhGgfv7vnZtC65i2to+j6qooDLnQ7mqXVZTltYS/wDfvaoQ+hHfK
YkgEZfUm8VmJ4Rj1DFyF0UcBspbTy8L6FiRgG9JqCMn2ATTWzCTt6Aa531cXFqft/a0v5wGrvtvP
Gv80OhO1foJKh3dMyNrnlkyvFfv9m7qnmJkQkjOprsYTpghTiQFzXtPWu8Tm0zUdGOD5l+m/hhxT
KhLUM/ZJJs7aGJpHzaYzRd4nWZRG8scfsEkWfneb9RWf7LGTmGG730RWS+d4fPOP7WfY0zfTiODG
xeWYL5BezkVgDj1w/4qdLr4ASy05z66xGuS0pJcnNWyiXN1nFeXtNcCJ3zjN2pVT71tOdmadv9Nt
v1t3482rqu3hyo6+68aBtuFD7NqAFTGj/lgJ80qRDHkb+nZCvCX7GZVyXtkpH+RzERWxESOdtLWT
dy1v0XYJWtOu6c2YXZEZJbMTtpqvfgYGuFuIWuFG6GYuP38LkrdbDFk+NXx1cvvkNxd0mgSsqEbr
5qLU4SdqnGDxPUqgfrv5VH9kkAj4UPJqBhXbK8JpvIfoe2dvEZ7rrVCsMoZtr4Ht+UZQOBi3Tr4j
ENOAkZwyyH39tjwz6ojHkP+gvRozIrrZ/JOiQ7Sx/GQqy9yhskgk6AKXnAJdUKfRGhKPQJeOt6OL
cAOpBVfiCcjaTdvdL3MJi9oF9npHKgN/1Ei1nb2N/s0LIlkYnluVJfaN2ijHKHeG/ovYj6cIhd3v
yWyUmdvYh0V0u7e00qL7ZG5NGJ8oZw7eIOMMA63rtfJ5vp29faaGXvuGnFGDZv9tEDQtvEfNrXx+
YzHqaKGVaYc8tK6HZ+64UWouCCtmGQJSBrlaHLAaHwVbIIVnnb26fgQtqlSakwHYFedLvDpxl0lE
bPaEoD2GczvBfMUfICLhBDgLCfP2oRBMgWs03S178/BW8xwXHS+0KEf6lK1KpqixDn0SE+PwHgPS
qMmL0JpKI5Bw8WFLAg3P93bUlnjELdK2K8nPq7ZIHysS9L10PkmVfCgm1BDxIY6LB8xgqGlFhSg1
L/gOPudshBYskeScQmaQGYSZhU6LKnh5KhdazzRYfaHsgigUyW2ogg3/uh0NJzpb/pqRCjNMlJZG
LwEey6u76alGgOzT7B+/g+w3ujuk04ZM8cN7Wq4mg1fnl1uRCKAZ7v9P5oeAiNcp/15dPjeC+kTU
H7wC0W83dfDByOHx01dFSGsKNmgXj0tFgjoM0Y1Gs8JV/KU3XveD0VNOYRU/y3jK+Mu2x0VoYIOr
QShpVp8tAtSJV5ueNKSFK47q8FeKQSxuQCGoxJ4BAqYx0c1zA9TaVkYuRYDCGn7cnqnTSlQ29Ja0
dsaledA+41N9QDAuJcK6d+8v0fOxK+Flq+aSvHA1VZF/rBOP/ZW6oCnxicPsfRFct3toDyL9dgOU
swwOmJILRla4tXDedoGiYAZPZIlduDMi8uSfZ+WKqR7WzVLguiC2K4l0aT6oy9zCeoL6ciczDO9w
D6rXNUng+1QgdrSLm3Pbm2pbQAkYdg2TrHPt9S6qRuC5N8sLdqgZKJOEwTCdL/8M0Vt0IuXe1WyQ
2QR8t0PxlAIZvsphEuFdJKLZRuqws9eDWdekoTlmtnZ8igcddqGULBJdGXfnokaakNdejY2y+zjx
vqEjH+2I0oCQqlXnuXV2ZBPIddOYUgBXGHQ+ljn2Qo4+dRZ116qHlpCyzY8a2yzpVyOE8/ALSDSE
fFIsJ7JLTC+3c4/DZ4I23SrArnM3TGWlNfCGcxVz7ti5mKj1jGV1bmHYfxZu8+hfVqbFw2k4rDpn
9nh6VjouckFLYC2MtXo8XMZb4ox53zE1e8+za+nT9619zGBTzNWR+edIoZiSA2eZNn811tABtxss
MnnpeECBUtnUoreDtJe8G6fukYzdk6GyM9QBlgIvsRclpgqqlbPA5bAth1Aih2TipvF3lHB6Eiq5
b6QySg8sxn0WXgPMVL6IBpBpb5+zJljLmL8LJ1lJmE7qiSLzZoaAT3sHGKMeclknGLSupOQa77dU
u8Vg7UTmMfxWgrhtbF1nuXzYp03QE2LaZnNBh2LOHHPjscdbSNUpE+RLnqxR7XffL2hMOMMri/oN
MSblIsP3fQNi/rNWo8c6E+YWG+1yH5is0nnCPgYY7nBp/YOBiRE2xNWNmYm/jOWO0K2ut8aNqty8
ml2CzBi3J5X0DKMur3t6uaqoY1foowpBt9XbQKxHdVf+wMccTUw4fqcJ8wCiPQ9nZLSHaQhfvpT6
m95daMxLM6tppQD4ILNUHy0DB6QsVhT/OnyuiAuFLRDqbzNj+xIVhTkaC3kABHJBryO7ZMBgQ1ag
lpCrLjc85JqAQ8lY8wxefDd0dQ7LdBAk+oH0QTXiQFb9vZnUE2+r5KqErDE77SVpFxtQjehYeMvQ
FC2+PmVqFZnspwXk/ZEwaMoVf/7ddKS2lZluKtMwFUZ//+Un+r0paegWUVufts7dDL9yoFXktvXV
QmJYqTIImhmKYEXnzoM9D86ZsJhxMN2d9OzZVucTF0ymV5F4M0Tpo1S2NJZYTfw0Ks2hEQTSeRIC
tVOBF40l7d/ZTPJmfO3tahqia3kB1GJ70iS48KinwOwWHGlqv2t4rMQOcAkLq37F9tKpkmU2bH9Q
Lr6KejIKeQc9c6mgqXPKTgZTHxjjihndAq04E3in0rg6zgo/dUn5ZPGY01fNR3uPSxHEYThzDkJR
FqFPCRwyjxcR27doj2cdDt5vc57YmDsDYRMYFZMY9OtvykXFiEcdMa4QsRZ/QlOnUkRvuBnGTvY5
OqpletYWr058TeKHQXMSHTyqiR3ANtWCMlGtptG8eM+svW6UehopTtLgFIWjB2oBurt16tV57b4D
jyzVn9LSuu2QBjhaEMAGBQyi7/CiLiVW/Eai+M5uMpESyIGwHtAV15qOWyQFjufWunH0jBBaIZXQ
r3+9GMqZBZLch7pv9Tog0Mm2H3v4D2YO+VSbSbh72U68qdk7P3n1rlzMxtchn7AZEYTUYScjQgex
prvDXjQznzKqfz8yOdbhIe5lZcmllyEBzDIhfLc4gyGOXJLFMPnOZDMOdg8oTl+Kqi99QXi9XvWs
4XeblftBPH+gjrhIGKvTo3CpFr5/9SOYOhRwx6kpzh8rojXi/IRH6dqYu/kcJjd/L/whMGxp67g6
BbIzyEgQz4h4qKPNXJCVe1YueY3fK4pqQJl83+UKe8KA9shrfD5x5ENk5OFhHvPgQIyrnw8+dVIK
9OIAewKnbj/4yBkpUe25rbVuchORbnP+r0ZDEfanxv2uWJP1bSJPQKZxV5PqY2lUmLRrAjQsOxmO
r71MXcLAlBTvodO/qYlKKx5QAdunHm7bmdgIU2M+3YI7jjbIV2/ddYjpPWUspriQQp9srdPLEhbw
5noLo0+iga/ACsXC4UNWlLVDitoWjYR/UKv9iGOLdKWwCOAWtJDDnv9OZwEtzm/gQF1qwUyMrT5D
zETRdzfe2voyjg4Nm0r1/8vZTkEDH3agQ1+xk9JE8RihthypeI/bkKSmeLL3vVMJPKlmPwVflZqq
kAc9fT0o6HxZTLPWINGOTDkLDd+OzWcOBnOHK7ddZfeg301T59E7QXK1wyAjSE6I2kIZU2IOYrxe
0J+SJFAUfPDh2jXGjxN2LrofwBIyMvLXgxk/toouRuo8n5ccsTaTs9ETZFW8ifYWnKI0UxGW0KHm
mw7JIqlSsKXdZxNS9iyT5HvClSyLkm5R649JHxAmlqi9MBXxhvxkLisNZn2EkL4It1Kp/4xgw3Om
rDvTVMuvDVUV5L82XE2hD6GzitWxityqp/CNZQ62GGOU9W0t3TMZIRlVwPESpwMgUFMOGcJlY2SI
whjfJcsRQBcoAOVwTbNFLj4SS+KbFb2KL1qvlI3c5QZGQoKDDurSNuqX9PQ7MAjEOIH+8BA32n5X
35WzmO3tFSmKWDzC1N4DaLqVNdwO6U2wXoFbfVQOrDPHOhyR/B1a6N5WYJixULcLZbFi8Bx4Qy9R
e/EZaPUf+7Ko1m1pTqa3bId6nMrEIQhzTYgnLf2/WtSPlViKn+H3ZzjXpA2czJGSB6hF5JzzVlY0
kcjVqW42y9Sjgg3qCd27yzWdzYJrqz0WUfh4AuTpFrX7pjdJMCI4fd+6jSY4aICWKjhF1PtyTF2T
gCEPkepXsdLiq6QycfdQQKpOr7Ssk2sEKU2z+AOTofxNLmF3wTLQM7JJ1TR2dv7DqnHyTwYdM28g
RfZcdNpte3jgmHGfYBz6ikr2DySqOhUI94DEV2+ON4aE9WZlur7vo9zX7jZ66fFeW0euajXjV/hT
RRSqMZQfDGMdDcBl2yXf3sBL3T5meB9S0dXXa6peHYBXQu7rnT2Hgy3z4lY+Gjmg+tQisG3EschL
zUUnsbTcd8SKKwMh7F7YTO6O1w4h8YphqimYQW3lZaNcOIW1kmDEk6688A8XeL2c/8LFAWacjIfE
qmlLWTw879xTzGOYfUPyy1tfIwa0uiCPKNscX1jZvzIF7QBRWEMsYKijmPEYWTnsLvSLEzEBa5nL
apEEjMrkqfMm59V3MhNdEe6u6YNfOHgHt43aZKgGgUIlIr3+81jkEVobo5YwGJOBToVsbTN23uvK
nK5yw6HkyofS0O/7YHEhCT05oyDs3bs3RpmWQvfcont7RuyF6UWregbQVVe9gsj3TtGtrzOYcLOP
+j700lQX94d45OYn2Kl2iLRr5+d6TTVDBCGzq8MYkzqgD/ViMoBALuNOI2p4vpSjXaPI7qy9bvl7
01RZazoKX3+Iw+j5qmkH5SlwvnrVfj5Y5VzX7XTve/w5fcBrUa0bgikmZJVpaDe/Q0aY3ldacvBq
D00n2PUyEJg1Hq91rEHerlL627gGeQhbW2piwXxANmbz28aGt2XDB4SVFV8sPT4EH3aASzJkTOE8
w4ru62MUuJhZM08cQKUJSYD+CLttSClfRekSfB5N8tgzY5J1THOXY5WuRD6JtuXupOLDfl1oXrOY
T5bGT7c1hI0Cy3DE0vd320wqmq5xGNqs9ZVPIelbFtcJI3XKoEeB2m7a/6T2vXkFiNSEKFy73/Zb
+aFwvOUPLkpFLjDUqYW9K1iW55Fr0xHc7GhwDsyz/QWS5/w+uqEReRsO+MgHwH1EoZwG3Yo0yUq2
85WVr8hGr5v3G+llV2iAc/7q2csX022B1GJTeaLqTMxPjyCLlhNwDiXMAeeUjDZxO7ucxFVyegyO
LMMZtkjzJ7VE52UTPJ9eLO9ImY/tcikAMT5UL2cD8jzXH5dtB9R54tmumvG2r8tvAppOkpLfOgc8
40Y7bgX51oOr8KSDMHK7cwiBacv5Tj3HUuKysCgsCeyixGEMyFavZjKE8gjVZdQ0JZdUrmW2sD4J
FtF1NE8LIF0SZ3uQtrMChYbLYZ+LEMmSY4QQrAR7C6Y/c+NF8G1A2leAM2gKzZCUgJZbY/0rCruE
sAE/nTnEU4tduGO75cquMuo0I8V1gALQW6TlBh5LFgM1HNUBcgRv85C28OUEKOBfIdqBNoMN40uR
B3v8fcc+h8XJBZnHvIIy7NYPFS/rMToPT+40g+oIm4NdD88CIaI78FcQLQvmXZDZrk/qpYLXjpcj
7NwiPtnQ8YrU4pqWc+aCex2rIVvuXmERUfJHveZskRIbM11j4/56AvDji3em34RJVBjsVRwLDWqY
mRysJLbzsFtmGGfdEU+JSrlAcJo+DnKRvXRb4VuqHkJR1Thtp3VItZ0XB58ya4xozCbMbzMRHWkA
ZxF3J8sC6pP+bfvsv5eoeJcrHql9rjoLN3wwGSgei1tjZqgdMMpyxd1w0tnxlCNGRjFmkjrDGKB8
UtGZU6MeTPC2fz1FoxvVCHexViO2Ky6Hf7RtV9nAEOtb0puAttcuAkCVURByCMeIALilMpiCM+mM
OKCfyT1ZROTKSrGhlRHh5ifv3NuKW11mk/9KbU2/zM5M5+lzscLpYRxu4b9/qOHkk0S+uFgON9eb
HYbZrAJw6qoMGrrhOG+Tjv3nZMOf1mVrRBztninpFoaOrXKcP3mGngqPJ92Q6J1TV73DwFtuVbwC
md+8KEBWj7nB1xx6EmEwuC0zh3gd1GSAmgsn7qMXw8xwfLvkDGTUm899TrhDQVhsVKeMqeSi1WNw
mjPoxprPaFYpji1lgpQvWuy2rVKylToUz4UZI76cTP0YJnPxQ2l2urxr7hofvSz8qCtTpBtyHzpM
n7GNSMocM3PEHiWnBZGWeMUmTQKp1SkriQFK46W0ac8qwTcFlb3bKC8fkkV7k4zvm05TNgmDRtJB
/IIIAEUkmP+gEhrDUSKj7T4j3I4Lm8YX6Ol3H8IoXMmoq2Qs+mF2ohHCAdb7TucJVFF9PKJ044U/
5QLeDA0HT77DcxTGQOsX9BxylagEoOGbW5tl1O18Z2Rt4UkkizmfgKN37mkeaskDSd5gp78yKp7F
85hPXwVgyzcnyyMlfPHLt2V+Y8IR9WNSYIAe+o7o3DguH0RhWj/URjoz3rjJ2FS38f/Siqrh0OeI
ARLtwuroRLucjPrwy/TdHg2xHmnv6aBZISNmvqET7VHKMFIRtBS9/1wdmf+8hMdOvKQ4d11eCQBH
mikwvBUbBSLuYD1q5B8EI0I0JHHOSUew7uoQ8xQ6GaxM3SluGCqnk0gqi4YcqFdfXvtS8TIg50Ni
Z01evrsABOr5i/Ae30p45erJJkrvJAAF8jALwqKUzxcrD+Ef7cE8LWpe+GbMcflGXbAPPIjwRHvx
7f7Aq9UrktPO+H8OETpJANz/oY5jhDAjpZbX9t84GetzeeTzIsE+mxPIgYhiw0yPF8ZRLsL8cVIF
uaOTstU9+BQEAMtwzkvcXbp5kavTl5wL0vU0H0GYZ4JQuvk83WqtjIdfZzCQPLVsyYEr5E0k2ONR
1jK+HJFQ6th5Da2+401wF+Xdgnr+WD5/PnmvDYc/Ec1lgpyA74r+bvYH2iOMupug+Noz6k87SAns
sGlYXGhSySF35jRg9z3smRyAHM8frHKlJPKTO0I0Jmb5pcplr52t7O3QHGTYbzgmjYWlffW5VW3q
8WCVQAxEsOfCH3+vSOcDM5dguV8NNH8nIz4wgiUg7QJ5gm55fGV7XPjUOxdBh54CZwoBXudOcG00
MwYNSERWqfcM80rA2v8culHANVckjJ0hlStQxzrR98JyfsOrfP5K5jCL932LFuYkuyd1pUvFUgFs
Ium2aY7c+1T2Sffo5Ll+gxDrIFlbNRJMDFruoni98G796uNCvn3hTYNFQf29d4R2RNQaLJwYuk2q
fDxxAZJsDQELrnUmyBsxFYLtinNaSKrh/2893bl4r+uGAWx9VCDn1HYkNMI7Dk6c14om3qgY6doM
cnneqQGZHHvAFV+KnvoWjZeXoubq7qwKpebjj4t4XSP2eOWDSfSeBotl5SEtzFaGcRjnma5NpY6a
XBJh2EzUlSFVWWeYyvLuiTOoHE0VLWIjT2hXeY8R4Y9kFr/wbWO2aGsuGnnyWl/11cHWKFNcW143
1VGYPU1fZU2h8tm3uTTprfCnFmOOFO78W42K1mMtGpL5Ka1NIldnOWO51rDrM17bKKFijs5k5DpL
2Qxq79Zp29UFU94yP84Pv+l6NNmeHGfPmOOqgiKegcluOFHAhQCdRiAJlr1BptghopeK4VxMpWnM
0CxzIZMEiSKOp+9M0/GxruNL1p/TaR4BcWsOillEhFWwM4nJGroqdbGijdeBSe0gGlgljaxGIIKs
ULfu7zMso8BA9gPbz3AiCNo4uDWv64Ixw+1/Lt2JBcdTb5rQfmREhYN5oKfD+8CvO3EPwvEOKvrM
ODGe36znIbwNa+hLFgvnINHtHMlKhbeqBR+/q9wZYZypK/wMrsr2C3AeHtI5vDQ1JDOYdgtyqLzt
4RzJUpJHcZDoHqx8RCyPKphDAguUpaAyv8r4BFYwasIBCWAdXDV5EpH7eSbpRAO8DXBA2sMsWINp
zT65aWfzQ7qL7pZeITbUHlKtie2MwlgYFrsjKCzQrradEJgtoBfYT7/tQhvtOutCsH+Iomb8tJ/i
oMc6OMNQ3x129JMx/VbkM3tVmVOLsKehzyB9kHguYXuNswZRsMcOTg5vkHT+VyJci1BLXnlRy7JF
3pAsMac55Dhm6i1NGU51zFM0NQnI1iysBzeYrexoR750Xd7nctDtv30bNvYdPMqihUIVQfRmHi1x
jAZ0H+zE+VZT2onDev3os+UnYPPvQOJXAUkGKSj5QHMQAjDemPXKkfgBeOqC4jd3t5bwkeYCrjPi
KJOvtroYB+8Erm1bM+rliJZy/Z2kwlICBlrlr+KTdg2qLgN4dLSmXmeM85kOa44wenmQRkoY3IAs
1/yMHn0PXAeMWDpndO2hgQRS7bjNnNGnv3FCslvfq+atBYmKuyownLKWlINgQ5MEkYz/8fvhgWJl
ebs6Cpcv3Lg4PohCFR4nKGYNe0i3sUCsZuLIk97UIGZucqMNrKZFhaPFewCIK1mt7SvQYDKaqDJn
bjwJmyNLBUYbMRf8U29Qspo/Y0JlEEwVRaQreWZlG/wZhqTsVK5klUiY2LpEbOZtcKBJZMjdqGb4
gBUccb4o4+wOZj9x+vzlT3JKAD7jin9ZDo7ZjCxAio3CYtse50SCaPgCEmCLI5H5lvBHEXU6mV5y
fU5GFCEqiaa8+xzZcIew9ooNUSJJDNWUBQeVnkIZTmTWg3ApmODaeYpRVmM3VqsAo4spSi77AEv3
Vht7oT05bzzLkRxtKtLM3ky9/KcT8QEXMLWFFD43QUCNTuu/b2b/d4IEE1aS4QneELdhWziakuAI
ddm/MqvSra0/5tJNxYA+yRiJMab0OlpkoRr1cLWT5puQ/DkJCHg4P259/NxkEbXqeUg5M0qCeV3n
BskJE/VGWdN6kekbpjfRZpXpxayQ7uT2EyV7r92YJ2bctolRa0KNK1sWeXwKGgbPc9Rurh95hqmI
P9QFNZqISf7dS2/d7v7zHEbHe0yaE2xZ/l5hHtfaGsQV1xt3pypCkG+h7AAgZOwD2cs0I0AGn68+
lfVTzpf0TZfyM5r0+A7JPPjw01rVBZz82FeSC2kuygVeCFxuspZG7v4LYTKYvoYE/cR1FFFgmSJI
RgFVMCd3rIzL+RcXtb0RJHZFzImAkIJQ0XLzJdTq/ZjfpS0cJkCS5CNfLOzu/sw22L9BBlQlZcID
B82+uUaTF11ti32ykxiMS6PdqSGeIKcU1dBaYr+zAKm/6Py/bmdOMe/n8HrRvB+zVu4SrNKLiwUr
6cv54ZlzHOJ8ZTfNmuGhoavYgMtzGbAsQOQlwrxLW0tqSoFZqxj80CXsYzobt005kJ1W+uRO3M+R
5zeoj2BJcc3pxyOIuegcNKZrziNBpbANjy5P9Ma+WixZ2kMPLp480b2YWfYocmdalDwbG7wJTh+i
IiF9O+NvKaNCnQmc4DAPaL9IA6hTMfk51/fztzuO0fy7OVEabba0BbLwsw7096S1NggWudaivnm7
1q58M7tlANONvteLgja7UEtrAwuXXHSOfWqBdd3vSbzMneOswN0OHON+d7N0IXXVyGRpyhms+vKi
k7ENOWbOLFF5wzoc5druHEVHMj3C6mB/4cURqmze1G26g/Or6LQ/j3UoMGPtg52qLZ3QHuaPRLFm
YlsArlNOyH8cRI3s1ICudXIQtimzsvTA2nBajO5Ru1kZkBYNKmPZLcPjkTEzGeID+LjWw57wGQaS
T19vt+04mPWmabxBDYag1NGQJ8YReYy+BwKYn/vkxs/ALOTwTmwFxb+AjhPbdBTBovW73HejtCkC
utgAddUcknKR9EmzG+7C9v8JeRT7pE155QgyPPqLxOwE7lEZNm9pD/WlrK9KslKHwb2ph85cnrGB
+y0z5KsodsspaCsaFztqnb1tdF56YUIvAdIVXEiIIh377Ov5V20o6As8bKvtebp/sX3jyn5bT7WR
NcCNV64J06n3TCUxntBNkxZkyZyi41G6xkTMTx+NbX1NpdEXDj3/qnANdlT22QNErCcol/lbeWRI
FHiqJ9WAePGvzl2cU8AaN3CYbs2/LnS0ryxSW0D7gcv9LepxbGRLG6aFrL70L7gcL26Tr/1DMpOl
5nv+WwQ/NoMHzC9ZJNNCkXoCitmH77GaF94t89og+CvjdNSkMCFcg3faAMA9/VfdSNROfTHm0FRc
QhbR7ruG64ubuzsPlqZvrOadyoQYXCOZNGBVAk/9/CmyvFGd5MeLjR3Ybv+pc6T47ydmVhoeNNSJ
ykL/7hTw2dWZIlomf7Srd2XNyi/74ZKAeXsN79HMlECQTkSpRafzuNEz3F1HO/Sc0ECu8WlULLys
UbPcRyD0QFUAHI/lJP8eC0R6OzFEdl0X1/hk32XJ/ThwZ/alIUZCodO3PYLOL5DfOT65nvfokE4C
2df5SoJE8KHT68KQsOFwyXPk7qCc3733yBAjSYs7IquOhYAi04vRA0fNPyMwvZ48X1L51TwLhuLP
wUA20CNRu/vTaS/VhPhC0i/mWuU6UB3wwmG3sB/OTkbFLNTJlezf6uaN9kQLuDymj60chg5+hwXG
F1HEJovoK5x1y0KBKj87osiU4+LpRQeyp9I6hG9zbKr7mBmGP23PioYiE3uJhOviMd2Yfoce9QZX
DBPMhgRpi/aaO0kiNBLzGrJIMXr3nncnATlwcB3dlqK+RPuTP/fQXNEi6wYFfq2eLA5ntsy4WL98
8czqG0tyT5UTdOwq2OqpCYyKSAZk9qfltlBv22DDFH/F/fvab4c17TUi5xc6ykab6sb3Gv6iSe9K
hYCFT5f0IDqkyD0fpokXvaswOb9KO8mCPxkaj8Diqxflf3V5FAT1IzyjLq/5h2tpKCfLBy5qLztJ
sXmn7DOuL14ZX1yPD77N2jCQzJjF/qh1A6epLZNyZLVw1v6qSmVQpu9ZbW+BQdTN5OYCDfUUeUt2
TtiDkCXYG2V0s+E7ipX8QpMZfsHG2/OAF3Kgfmn0hgQ8Tssv6DPN3YYaCdlCh520Mu3+VyCRyvTW
KnzNU9s9p6mnD7n15g3zHR7z2PKhJ709VKFZEypnazQnL2Z3Sc2C34TClBj1hZk4iShGOk9e4rwR
5J0f4m6YuNrY2tYBo2qc3g8XphzdWkGd1nx4Xr5Tt2iZloMqCnAtRTomxl99FNen6Zm33HmqrAgl
kDh9+Ik6SWKKXuapmJjozQbL4Nc0LfMPt873NqobGL8+sB5Q4AAbP0PrONzP2aD57yfPXtDif3I9
eSIVKdjG0MwzOUCYEX1CDeUFinaF0oB8+3E6T2ei+Xrw/y3jq1udx3CvCjKBhPN3+XRRdWJl4HCt
DLiv8DPhaN0Y3QAqFM8JBl4IloJSawpVzvXZ9SCjDqpjV4Y4JvUafs7QwNfkrxMhuz0/tim2Scc9
JQsjkM1w2TfTEnJ91WpRUSYGRQUkVRoRP1To+qZUhMIs2qjXE156mEbc4svA70iACTGRbnJAVJ3J
/xlwQyU+uJ36+eqwjkezhygmYbbb/mZAPZWiFXGyV4P5xjzFeKZiCHfbyBw9vkEGU7+V4ovLvqfd
UtA5KyUwEFhGDvrTyUOEnxbz5uwmdA/Ex9ZOMnZ6YxKxMcXH/2lSDk6NkNMlGH/LF3af6StTz9FI
1KNCQL7Tn0UeljfRuEGbDItV7280ykHImh5I/CkDAU72s3/+lQtxuGCbbNK4mdF9FFiy5bWL3S4q
lSl6ue5mgWbGAvm+UszRHtQfqZOrJi5J5L63mPkNKiDpWQjc+Oc9zco1uSlcZIIwCVuDnVGLPTOu
yWl7zCDm6GkGAmOlZG/mnI+hM0z3WInLRte+03GdPpcLybzS95Zes34ngywODbhCCggZHdX5WeVV
9tKbOs81zfhcOEEYsoNJO/lYM07u0izFUcGyrZbTAnUixvE8u/7Kui/f9PEjdl7xBXHuYU0NxjBs
3zo945glqwTtQDxF6cMDNrW8RVlJfDECm3h3s/i3L0xNucYzIttTqvBJrbXqGv4gR8spddhOBprR
o4jxA7iBZyqAtOpyT/9Q1H9on1jFIEuzGd3aXZYWJZ8YRvd3tjCyrBReLFm+9fK+0sEg1QS4tkuC
ZGiXH73/EbP+/hmn2v1zVn6i6KQsYuu6bZibkfA+fggc7ND14Wbixl5FOhaNGkoB/Jq5aQbhYeXq
76ik7ak7f0MAYddW7Sli1CUqWnlgxLH8CxuEPQ/rbOAkx9lPkZq7f05IgE86LozyvQBNYFjhE1nO
OgJyBuHyMFK7M7DedzFUMwpMXmOr/0es7r504rheAgk3F58mM5md5wy9yqmm54GKHw7zZVClZv3Y
0skSrEL52PIg8tRCnT6tqNe3BzrOuwaigh7Z42XNFKGYbWPMMEB6gAayQE2JX4HjxhDbXJqanNLe
5RlEEUBy+ZBQ7gU1yyP81GMIO7QR2yhbx1TYnhPzPIR3Wr6IwgsLch9Fgc6N65gkdMigQij4gsF1
NLH8mEoAbj2a8eM3dYp7phZP1ILO2/SNoTX8nIDwMJnNfzy2buVdCbXCp7lkXRsqLd5rr/DBOKiw
YZ6qDnAZcNeHChI7k0MxPa1l4yHIrlIIINdGoOzddr0Qu2ZO3dLIPaKRP4MQGTVZCQMyNd0obHEB
442Vx0ItjKfGd8lj44a7S74Of8Jc2h0vkVHlUCJM/ptJ9TDjiaCa3vda2n8ZECAskY2z8AvyNt+x
SvvBPxOoEKHXhAyYUok0zkBRbkI3rmg3VHwWD31XMU/yR+4RN2PjBNRTHLdOlwEtsSPvw/zwTye+
vvAYe3F3HbI56IXUTof+7IFnR6QKWdHTLiLTUXdIRGv6sJmVdqRNNGUBi+tnvfBO5RvAl6Hza1pV
lwgcw5pI8E6NdeDHiQUWpoQZH0GySQkakahgB3a6OMYTRcEzYDe0HAr4WWxzvUhYP6WIGOZfLCSI
ujhRmntKrSfl/NekVDzOVdRyfEP3UgpW1jDar3sEplq9X1SmpC7UjEQYCdCx3ODITc0hzmBmhNGv
mi53osPuO1SFPE6d3BhM+TA24bRyCR3k+2qAV31HuQnZtVNA8naMHZZRJKS1YEW1YeaY9Vqur0IB
QupySAIqKuOU2IG6oNZpmNSZP9lUOboELYn+NVAQZzmpLk7Vaqw8OTHHoxNfZ7zhDqLnScVK7VpM
7zYx9m1lJ9QblE/s6F84s9LNuJ3mMEb4WREO8ZCxIiPAuRmW8zFXtlRczwNWVbTN9UEwdlGCKVfB
cCRIpLxsy5z3Njaz6yQzc4tbNY1k8NLK5rrd9BuUc+78aIFESBerbR8IjZVpBWjNpWZR95vMzhID
SbRMIaJJpVVCswP6ZgglzfCnNvaTpMmyo8VTKB5W52EbUIpfJNHE0ZrMS2aYymGYSdy8Hrr3dtik
bSFaIyX+dSY2Lyb/YqDh7ZJ8WlE8+n4O4a1yMzl0zTRoC9uM/2IZQZLjyjzzExk5ZyUtih9IwcyN
Vgt7w39f8dItUDo49ytQC1Q7PIP+Q7iQUdlMqjWaF//qc9YzT68GaKxfM8iWpn0l2+UnR07UuXiI
ZqrqaQVtXLUM8cexuVWndwRo+5YCFd61ZmBjbDHA9WyA5+3IxGL+pzjmsAa5RylcA5UkhtNqU4e1
qz98/NX9qzwuEsilTUpLtOAcL0R2eAoHBkSOPDPdUNNddIZnuJoZSyn/V7jYRAZNxS2V6DEsutmM
2eNSG0O3vpv5hdCXsEi1ZZ6ex5ewTr4ftFHk6unn4YLebNLKcylFt8XkxZDteY87fo0vfgPPepcS
8f4vI5IMQIynYYOmi4iAedR1CwphzWgYAw9R6cxalpsM0TkqUHyPCcKbNgu7Pl3eJn09vIEHnD6j
uK97iI6NTRe3Q9PWhWdoQhei/uymNgNAkyWh0Fo/VVx6e3rryG5ytHjInz82hJQMIm8SMEBA2bcp
TMGoYVeRL/SmUW7ClfDq8Smhj8uftaSau4Mr1E0Z08kOwaFclZFz/+15uOhYjLN/MeV0mkiQOKNv
+f+wCkMVNLuAfOa4Q1DWcQDiZ6SnxtiiZOGXXJzDEHIMBH2ijk7arUCK8DDUiXvOfPrGlL37XHEQ
4Yffqf+wIdes6/AzDviPfy6gBdcw76nI3YF5WeziTku/x6ESdR9Jfwyd7B4dMOrmDb0//+wJGCX8
+lI9iKbAXhijJBMSRkqIYrHXsxlbJOfO2r7g2F2XGbfg3cEBpz5ZcLrHtYrmcKDzE1KHtyvhhGzD
2YiNqGnCvhIr+G8wL209Vbwlsaov/AF3d27JjI+Rodgb4E3Y3cI00f3AoGtqXyoFcphX02UBdvVq
TbC13W3vei/pPemthoL0z/sY8y28dalZuPK0fBwlaD++qjxRF+NER03lPgM0jzmPJEfghj3mo05g
g6MkmR9P6ID6I1kMTBUEvw+sMHNJ4loDtJb+cgjmBuS8RIlYFNNFS+P7gIQVxpy9l0MVpvOfLVyD
PJOb0udqxoGaFK2eYWHmezlnRu9nGR36j2nEg0vpLvBCuu8zq8fYJixZuSBnFGEVKLx4TK3t5Pf7
xDZRnuyi3PQcBo3192JUMlarmsVw8GCF1auzHoBb8zxRpAvh1BqIBnEtLzWZUSkzHyeywG+w/Sx6
MJZ5VgZE0//zBQNocRcMTEuUbJz3fLEwrOA+RR336yuzNmsqwOcVySU8I60KGjaMC3mgvH4ZZRQf
y2RIOOqG1v3aQJOm/u59wkWLr+gv+jRbY8PhLFmMoaLsCWoMxZBg7OP2qdn7KkE/gRZqRVFZLovp
QET8sRoKD+1rjBChtZEI5KJiwjpD4SI2FM/zmFmqytqZyaj6Kc6C+VnsBkAR4hUDjxynLrwPomoW
Bd4OFRdTzq7wo5tcJA19TRVuDv1gNbDR1FfHUU4cOMvGnS8EtP/PcrnN+Kr3XvSx9ZZQFO991W5j
eE0lsKRuBW0Q5H2kB9SDmrC5LrG15BkudcWo90CJCbaOUPe3C/dQHV3YhJgZbMqRMlnX5dUsFAni
Es9ouMOhGAptyuJNn7wWrGzhnySo8L68X9LYiUzyyqxzPc0JRIRJpuECVpsS6IT5q66ra+fjCsXi
usUE2NcJR0y48Lts/J+eyDJc8XWDxg3nBwGMuV117FYk07ur7ZCUF3zFcRfb8u0FfbiAWZkLX2Yi
rF6fOn3VJojqGJEh4B9oY+TmDmaoI+uxvBRF1LDxEZCB4pn86eQNoLkOBQzwifjTGCfn91v3HF/K
hb4L9DBXXLfNgcnrNPa5w7hlz3k35Xo5tyD3Npomj62pKkLnhk9JqVRKD3xky+IgGOLF0Ns+uI5K
MmwvimF3GpJnbyDH+lOc/feyZksMi5H2VVlJVZ8F4SfDqA7eAetxj6HQwXSe35SoJs1YtE1UUdTJ
Rbi5Af+5HSx/zyCumUbw1hX9jg4J8/FM3HvUw7YzAsYhUj3UyT0wVzY3dgpzeQR/r54AbfcOQ7W2
D2WjSXRI9EFtSGRgUJVqDdUwllpbG4JxjwpFaVrx3ynvuQqNRtK2pPLIvJy7a48bXv3Rr+NumKEe
yfCVtrfNzbcfmp5fe1HxNhcyzQgZLja9mJTIyIMWEHkdH//HgfttXX5Z47t44IdvOLP/a4aPJE+x
zF1bRwqNvh8TBAH96mX1Xs6IiYBm+UmEFTpLiLhRKt20xjwSBNsIy5BNq/sAbOF6zowEXI00q3GZ
wSWjIDKCT93UKgCaBQEBdiJLikCOE9zgsDOW6RtyKQw00yKmdvgOuX9jvNh8aw+Ele8NLVyxX81v
VXaGjwaBrr01giVi2dL/laaedeKa0+FxmJYrB4YN23668qHzOw4b33CiLIm7+1NYo9kvwW5FsTM5
RfA4gvOrxQm4qYHVoPLFmpo8ARB7wAE762od8sXAc73WOYj72rlUIOswnPSPfigrrTPipdK2RNP0
MW2/WkWVq8Kld6j9h3I5j8fKL2r3YbxmwPAm9q53IdnkoREXEY4VnV52fbbljenOgmSTcLHx77j9
cmGdsmoXKDsVswfYo9blZtMOkYm2LN1hzbhmkvEwfGGXztTjlaOdAJZ+QHuiXhE+Qp3x4H2UKTIO
24GsO2lQwUczQSYQ1rd3Kt2m42tLYDn9tE+5whc/fKsdBzvvG+ALK777E4qHrwEFm924mFDVmVnE
kqgr5L/uiP/Wudte7rtE6vJoxMFbJBDsJWjLJpxC+jFIBtdSUjzJH6gj0AEy4j4fXer2AYPqntUp
yVF1mH87F7aA56aZla8DHJMXH2bcO1h+iHVE+oSe9XMn09B0hn7VmGoueSnD/FM3HMXn3reh69lY
cmnV3xj/JB39hkXv8EqvUeZB4ucFTNVqH0V1F7BQzxviHBWvffWQCUVaN944wxJqs+Hp53FminNs
MQE4lfj4LbW2DQUDOSHsKhHvOkQZFOEmhRi5hmxPpeh359Su4Do8zoBsB8NipBoOOCIGDHF1ecD0
+b3QAE0OOU0k3dIfdSOADLiMs5iDBH+eVH4mcjDBhO4H6aTiW97UQEQMjCr5n2/qeFRmHK+JRQst
XEugCOFWAccqj4+6GEOR9EYOrwFtL90fYX3IJ3rWUfN51p+EnFEuFV3682cTMmDCki66VmTCOcSL
LeAtj5qCxVqlUam6+5OMP2O7rspPGfyVo2X2cPZKIwb+SE61Z6aH+AYc1+atSMpY4/EWo6pqEAYg
9g/sjaNIFLIAMjnUSv0a33dH9oqytijTNwgzflRR2arsGuXPtT0m+ReN1SwChwdOBtvbBRq8J1Tx
7MQkF0Q+OCzSX9Cg/QKeXCQptZ2VFmxnUu17geORoHjoPHxhHKzJ5Q418d8Y4KzKBZTmErk1hHC8
C7iXuLawZT/mtl9xE9W57WvVjXGcBx/Mj6d4IxdgG5Etrqyi44lpAhM8jiS/iSku1ZrPRfj8SmDI
if6Q+lbWtOl0Hw4KoOTMRcE80QV8mWxC5xTtG3GYiZi8NWGdaBdNzRK+Xqc3uWXDMlTO5iQ86kzG
HSMtg5PnfQ+5LiceFmBwWNaZBY+z7SyAgzwoGmf2qg6yFHuDA7Sss2+2xjGfM5URS8GNSSD8Jq5C
/M6m0A8MEd8EVry+OYkdojbOOON7FxfbgIA0MxEYiWLxK9cEPomZS9ystU8Fcca7axJwYfYX8Doh
ksYk4Kbn6JG96ixhMGX8dbd5gFOYe42ZcTt0rVIEbOyyLtGQXTgbucs2jWCPE3ymkug6inqwVMG3
zaqjBj4RUEpwNJoHTg+1bmyXcwjAWPhhEFcllqilohanPUrPdarv094eKfTzWPZoTNPNCqZd0Qv5
kZQOZxrL7B7s4QR0tFzL4DodAy4VU1KbdVLPA3LPumwg4tTwtO3zJBWw0bvbft6ZD+ORrOYolb9a
IKWOPu4yB5EEFfRXcOhJ2jQd0EH4BBnYCazxzOL/pJ6tcipy4Q2kFgW5zTBP/Li/C8nySwexFvTV
MFSwHPuFUmevQqi/6BuJAhsV2eiyE69BDOQ1++rk7dHrpRJ4j6C3KzDZuGlGQiO8SvvmPs3lRGlx
u7IIb1XHQV8+zmySn/EBhTkEpo4+Pl+Tysg3Qy/v7x7rohVkXSRo2RMSEZ/SpUlm91fyDPgUxgKE
xLuqpjl9sa6wBP1VznPn0x0vdQcS+zFeO5MD7bVaQSCysq9BuMQN37rR9LvWwLFInr2oxKvvCf5b
KSVI/Hz7kolnYrbT63w/JjaTpQmyEGyGXVZM0DxyAhOEyZvLKBVyE+J1fEXtNqtGbhLqohMTGhWN
ujzYKkQOfIjA9cAe1lFjuhtdxRzgWQpedMg1mPegmv2RxHrT6RWUkiohhZQrqKajr1FbhUfwi+Jj
6XCcYl8fivYI7fdbwX+HHhiuzYtKbw+ENnIwmSXbR82nHlKd6jAQeY0liFEbP/k9Lwk9gZAq6BcR
6Br7F5fqY4tFr+wqQdKCfXCBPsVF3/YRDonb4hKwY2JJSogpVU3cPf1+bFxVmeEvoSQG7dqY1tpP
LLCL/NLourGbMj/IF6GDCwLKB/ZQqAPkawohHljjDPEARblikbFkRxJ6PF6ZVSHe8USTTh6Ssr3T
23gzNPsYnQSXOeZD9gYQQjXV3+bnb5Blkm96DV6uuWwLxJKrF0WpUwofZVB9JZz0D7UpLHx7Oced
Ft0XOFI36u2Ucncli2WciRdopqck4jZeeMacmLfu+VlDBVOudF33L8nXUKL0OLGFkpws2QpRV0Cc
V9I0gFcbeEg7wSkFMxlB2hsUmFow6wwu8ebwTVbXLxBgu0y+iaunZAwGcSmI6755v7pX8aX69l0a
eVN1eubNDcAVyNUfhWvoCJSqzPxYujc0x8olnRtBT9kV+3VKxu+99/reuc4HypVL36oaapsISs6T
fKvjbG1Lpui2lSRbbzFtfkSGRmg2ISDf/brb/0KgCoKgQP9dIfdXUbtWZR9j+GrVUewP4N8BLycA
bv/llNS88XvFp21MUSdjmXRnkEUHb+Iz+UkfsNh3El/lCZVPJcmKfC5A1bDhMw0bsVQUAzWUgm69
1SJTlHVjFOCjAXyC6qL/5aGYm+pPoS/zT6W2OZFO82gOdeszeigfQ0eaq/7y7TG/X02l8h8KXk9D
AxsTVHHLku7BHsNX+W2XyfQzd4Xt+4CbLufhUGxuOIq+cH8Soo+YIHXQVKBd+bXxdYb8fAx7Wt9C
/jK5ygBjxWJou2WQIJarXhU8ZMCFSEPBpyZWi9WJz45h1Ndi6WiDJxfb1qpga7I2bjcYLZzT774B
np4lLMMzf0xR13uwnEfxBMkBFtDn2PgSBouYkBAI1n4qQ+6iTMpACuq1HKvNj4icrp4kWe1T9ZyY
JZwldl7MUCPYl18d+zENYisS96MSV5Xn2cHBLXw3kKx1mSxN2qLMLqQHP/XAeDrQn327PZ/B4IIw
j7mKTVLAEwPLM4yKvV4s8doDQsStaPC2u1yRqkboJ49kplGUS2w15cGDgRtU9TIoaarE/lSvAbeM
ZxbmAAjpXDhlYMyngP2RFSASERuYFT0XoPL3Lg61prsrEzJGqgEH2BdlBBXJr1ZnBLaVH+mZwoGU
UbfG8xLCveZw9znUjonADG2aSRQtwYglxhyudAMH8/ARW3bmA/9PHiizPyzEb41KB9oM0uT3bldv
MxBgLu+ilEMVvnPCLvOSNHVR3DJTAp4D8ep+YjZjxFvv7rLHyQfCkOtWELsyrJVICEmxsjZUyKVx
DJYTZnp1GweR/mqqHWzWS+Vpq0PcT8rnOYkY0zk58iB5j99F0hOsqWkUh7RfAutUPeSNDqMf81St
NtJrYU8Vs8tLYW4yn0r48g4zDZACINTmSB16IeF8eTLY0bjPNFp3rRLmW2zkPFCctfTZMWu+tx+e
mEHr+5ZNyrkgwOqmeNlq3H1ZkZGxzOC0lhK9TPuAwRPyP/h57b5aGelmoXk+flsHZrG50gJEYPCQ
D1e2j/uVSTDMwoaA1BjyZ+3jbovMU74ItFtBDuGRdymKH88vrcrCkgA2LzKE3mEXnhSBOuerzQgJ
1jJ3WkZmu1huO352NHL2HLZ9rSOZyM/jE9xOEyhprQ1JXgpvgy1FXjHtlRVmEieBJyXcIblwL/0n
F+A8cIDc5a6woK9leDPRngjkKgwgLony/NcSnIUj4YuwmSZk6lZf0e3M9t9LZNwQJo78/3BPNDov
DAaaPkx5n81q9EkXzBegSvwHks07piNQe74mxTxne8LA6FZsaQxrYZOcZGw21l0vQ9WUz0Hje10V
pQo6lB819QxW0DX3GGYIBGbUvSDOShDgNr0moOFDf2Orrzr9RqVb/MjxXBEhFg8au0THnBHnrkZ1
j8UhspiDQGLMbKUBC+nxdwJozge5bFh38DS1yFJgpGABVaBLq8vTyMBatwa+GOy6c1OmVzudZI//
w7iQrYTEqTND6GqaF3Ica9YGsAsYjdIFY+nnr7TAETRYpVuEEdIe+fyLB4kYStsUhScf1qy0zAiC
8kQLeLAzeyJehZwuD7Sw8eKg46aaqkgCq5rj+E0Qizv9lKEqZgOEGFtT6I9lAine9ivjeAhvJ9XA
k1JiOxMfYiBaXSpikKg+dYAgs56q3pxp8/4IXMB5G9SiEyQUwcOKwBcnb8XeSMxVYO+NWkFPu/PC
mF3+Pu4ALyOA/8FuwhJXjkCsSDNZBihPFpZ7KebuGL2O1jzT5ywZvc0G9WL/DTo93JAxQnY/SAWr
q5GFRSqYIBgQB3HoSRweAcd9/UaPMVghr1qnqQyI2u5iR5dlmNzlhUJqo2iSKpxIUpashboEBqso
p7cXehD6LMgHClqPqmgftN9roHAyoV+NKXxH3KqIGBMW8Vj0pYwucOBlBJhm/YwpmThSBdUWYNc0
62ngIm6BMRLqi1vnsic+J7jmGjTzM5/pGEvkxzlPSj6E6h64iYEtJVYwQeuceh3ArrNZHswqUjE9
rx8CR//cL6jEI22AyVDRfde63yXpTuHdjAmKnSjTdfSKVD60QEYmhOl0NSYfgjlKPlugCZS6wsek
h16VQ37VmrJFpXxv9gAtCIbZxwdI1hEt7uFfBnVEHXCr2ziQpIxgt8Sd35wNgRh0ndmB7hvWQibV
9LoH1shtfKwc2XfcvQWjNzfVB8CvrAd6JGTjfGjiUs+kY2tGlJ/6s1wyrfj2ML0g3INE0+84DqHw
4pHJkO7t/Wzv7+gN+Zmq9kXOLn/CD4mbv88qDURYKTiymS076m1QLeWG/UfoyBUneYa0TLKYBTNy
G+BTE01befS1dpNaYianoeMiNt3FHkEucfuW+K5YNjNC7wlvwXhKSi5lkIl/jSOYyWNgVltxm/NM
Cc6haUSMdXAyItT6ONihH705vmv1nRSn5k20J9weRoet59Cj96ZnTbeHWG8J0ZpGvN0ozvLgNLCn
Pak+S2GgcLJfx5lu2WbNFwvrjpOSCcL8wAhbXJEK/bxd080w4JZRZeDHEvI47ufy79X6QJATm4aU
c+IjzWzPgPn53kKdePmEvCWU8AWQNzurQpjLfMgZ0PzEUPDb6guaOrOQC4ETVbh13qN4T5Mew1rT
68cPPj503JZafFoCzrBtWHiI0zr5WA2YlMb5fCITN/ijSqD3xL7U0xaxJDCzfm9uUUktAjhsVqgC
xq1mAuADwcmz77J3cAWayFJPdF9AkTfUuEY1fmvkLLy5TpwvSnIw3j8l4iDjbAK88J/kc/bIyOwH
/4MzovvMVSEInDpO0HeRNMNu3s3IEguemlLqZJHJAG8yAfDyzhYOoRLi+fYvp+KcMUJBXzKd0Sx8
0OHjo8jMdnG8XGtO/zGPtpyZTBbjzDPTQbrCYdrd7jcGbho+Ip18zT9ukJqQqI2FhxlNBWvix95Z
gzsDjZ/3NffsWAhwlDOFv181T2IOy1gN9nlkXOr3Pic5u11MDKDNM4VyzDkp45X/6XjzbYr/QVtH
Swbcd3LNSji+kQH/YzVkDI7mKQF0OAiozmkwgH4lST4lkLNie7YUK8PVefatUBQzuJ0Pkyi52UgD
R/IPi+h87DR8txFP3Lhyb9N6Mo8AT347pv1wZrlLATTwMUKdR64SMBX/lopMs1vqz41LmZBeRaAs
8VnV8w5FxZRu66S2m4ZKiuz+grLYgDPFu9jJhvt72RmF/ydK3MIsm8tub0Ww9GCnCLx8Y3bWm42g
PcWn+RG+PX7mHZdA3dzc0iHc2zSuhCtIMTeu6HOZKFWbINjvfiWSSDJxrjbeG5BxMMrcOj+GWAuu
ul19ZEaoFPPxxzomAGNd0hrIz0qxkwBaPR+mrRdsXWNXiT59rYtwsZcMe+YlB79oG4pU5dDHYyzS
2M/j0emnN9R0I2mhV2lOgTH0Bud7qkhU4HPR+nCi4n7MUBMIT3Ro3TSMArxtYryugtGcvu0XcbzI
GopYheSzpL+F2WRwtd15NvrxJmE5vQwCr4dSP2zDmyoHXAQ31eTc3lf9Bm8fRcSd6O9JM98qleO1
KhVnrORwGzA+Hc8CUEALHYO9Jsydi6rXW5jyd3NgBNTvpyIi+b33dpFQ/YB+bxRafPsuESIVq7cI
KaG38/C+5YXhFM3isBoBL+OhZ8/W0fTBxcK8G3bNDTX1xpKlGtVVfKI9ocQe27+dT1g1EfvafuW5
yTxsgjvEzPKmbxAXX6vCUsLqzdLuGTVN9eDVinb+oCwUQEgfkFPaOgaiDkBIEIw4W+B5hHWpaEwh
WpbWzAwekhYZUqVsEzKy7cBQrjEliWHfkSY22v/r950yts7Yy/7IZ/HxGv2ZllOELth99m1cciRy
WAJ8u3xQEc1JSFYbWckTO4QJRdZIzoXxPk5PiYwUhurPCjXNipwXuHkv4tEEucqPqlyjSmUVHZKE
zfZecif1x71nuddQdoNWccUopKluicgeC748tEOL/mTelkrBFKWa6/IlY4PZc3rMb+Jc+ANnIsU+
AthBsIKEMQ6qk7xLWppYRFLUzYJAHk4fxlq05PbVCwuYHN/4M39euPQURArmTReUEmqAd1j/t9Lc
rUGvsDHuapQxLUJMH9yJXvdTCsZB4gQmE9J+cx3Nux7JRLa6DpOWq0LGPkQv+1B4viQAlrKdMjew
u7evlq1+T+SHPZRLXm7q2WUOnzkDJMsGYiEa+SoJFRqbkmj78T/UHyiCncCytD4TBVMvO9WU+0Zw
ghzSUs5lf3lno4k3KBYDPfc7Hm1QHRN3ykEVXbAYAth6+A4NjQg1fa9NXDDxxjQ9VDg9+MiWM9Vl
/btGLRMYoCCmL0zkK+/AcMVjAttfMSqng8sOWEJ3Xn98Ospkrrxc4QWzRLOVAH/iKTP0uxVTf3SI
6LwKnDV1LFzGRlnQDiHdfCgZFjk51mGkCuTwDbpRVzZCVMSW34hLpwnd2wFhRVpvFNJhDzd3OxMA
M83VylzAHO6jFUADe3C5P12B9+e0Sae6O+ORZfX6JRptNrd1gDcAdowA5URIgH1FeMgylv0zID4d
l4drmiEa9FkS6AwUtOWUm7xQaEggo/34JH5uU914NIqxRLAxFztABvFN9b28m/zw5nxJiHYr67wA
Im9PiU74B3yjHpbWarCiDoQjNElfvGIRrSafyJJqy67xnHe3YkESdCP7sVA2cn+flM6ZgiA+AuPi
567I/1mn/9OPkNXPPj42g87Uqmeo8Z9BuyWDkGL6XF5MALdfsI9MW47zZ9Wbrosrg+NiQAIkcQdR
71GcCeltgW7i59u1Pp708Xq51q5XdTTaUxehQoAGRKdyUZak/ZcYk/uwBxEUmwe3EbA35USk01Iv
8bCq/clksv08DiYztHi/nNE85GW+TeRStPIwr0AOXYIvg9o+3kNp974WUyUtHKkxlfefsKH8WaoM
Z4QW3K7Hcnwiuj8kCo4FeM7F+G8KrHic02NLUcKaldebKR3DbLOwquxl8+swoSsXqk8vRoFmR8co
kgwyz/om4TmfgOzV4g/Tg/BjVYe7SQW71yFx1fCB/vvmOeIXCs4btRocupR3mxFK6dDeWmrxHgDz
zp6Cxa85spu5OeuvOzSQguEH0Yr3R60AwvfB9sPnJlVq2sbtbXJck8e+UhcYrx36A9GDWDxYNFHr
Y7DU9eveHgVupp76toBSEVuVDtxDNlFMrO01xeoa5YnGQ7HARbNKQZHVo4oqFbtK7vWW/Tsv93Ix
nCHIEhLDhwjw5ybUlY4oD47eB+Ya4Y0dXYSbi7Oi7V8aMvX5IV8X/NAkM8qkFw8GTp3ULDAcH3SG
OLXesVJuYcETvn1vpatC8VRaR57ZUz5YTBeWxBHELFR+CA4gYmDrtcAJcDSEfzWONb668shQujsm
Gfi2Z+4Dp1Gns47iDFyAJTlkUd0xfAB8fyky8KVXalO3B2Kuy3zFPa8GUrt05YTwQcc+S9Xzssft
oLH8EEyokiPzQs4INgqszVPo1VNZqI5QIiUm2CymwaIFmk++kP1PAynQtq+9iiIDcvPhKWZ5nGEZ
257ZWs/6w4AoIg1c2vLzSLH8QemcaV1ucX9HcnN4V8Idj9qQq5WBxS0vTiJeYulh3FD45cHqybwm
bd+Ma3brsg60Bxm5rvNr7rA+aVYnuqUYCUMUelwJCytgderru9b2JycSgsoLtZSqHMMP5mfoRT8q
JnyTAzJGAguiLjNuCt0ATR2+G4YkFVoutIfEREgpKnRksddyXf5CORylbsr4qk3w+SZsrwUEuaRP
c3TyEQOPhss9LjbYJOIcT+EjWESgzrz2/34sR4Vn6qjbpPIQoJHlyel99W+h+zA5DLhiMJBfo5pz
QppZiEC43oj7L+OcjI7H0fBWtlxTD5mU8rfrzebMDUWqoAhrqkgrvv+52AvJrEj3eeNhCTF/7S5K
5O5doww6yKHC08qsVguss7yuBvWYPowyRj9r/WwIixEmBP1gPQ75MzBWOAt9hzkXpEdBb/yuqUfX
LTNaZO2XDRdKtX6eBTHPIYNIZfRqj+y1v/UGl3wjUhfo7LvHgjqbFpdimcZDJE07ace0ur+9vYzU
fnvIzOKr9BE6FYm9m+sgLXlQm5RL4vsTnPK6dp29GZ0GoRibcL2lxZ/aMVb/W/2lCXNFI6iKjH+J
lEcz/D6NxRYzl90S72V/ThwbJtntVxIqRPE6eMzgS4mboL+vd2zf6pbzpQMiyrrwYa5yK3+hoI5H
R21yNMZHtrEpUDlZWHqqMzRwi5nZGOFEAu4d/LpqxJSJa+dQqgCiJEEIJUn47+MLsAtzlbvEGfpj
nbVz5Ows8xFljErdx0+uNW+ia3wiroNpqJGnZGBE8AzGrVE/iZjYUOhCe39RH47WL6xWKeAdAd8h
6AQN7iwj2t6bdU+tVMCTRJn64lKobIntqEls9lMgbenA10Vbsqtb0y6hJePQK7tOEsHospl3ur/0
Cj/Ms0SU25RpuKwseFHPEEqXUWOHXnGwx0hPm6CjMDTxqUOeWcxCUUCsc6tQKAwyAMDnNw3NFb2q
Xemglqcimzrpaa7oP351jzTA5YCTygi1cBTz7/WOrMeFaArQuwiDxW+HmVqqPhoBRriPcgVDEl75
YwFbyVY1q2GBXKzfAPFMcKx4p/TYXRl3vyqu6+mqPcls032SaoPzqN+Wl74g69/7WaOGpPF7dgZk
fvuPT/ACABPoh5TqGD6ZhDDvzE3G6tQ6oQgFl8gcTS6rZLMaXRjY/MbzViUFCLea3FItLG/MHQKl
IVsWGVLU3gpejdPgAUthzYxEgBFABmKakLR+2bRiCeroqHyUePqLH/lxn1eDHEuKG2oW9oqrt2rv
zInRHYNezPwDF1FdbFXzwdcLEZ45T3rOGrZMNyfFttvbvCwGXwaJ9oU0Ut2dt86UWevh2ikzh3Tl
wQouZps7gLpgwwlo9P6gurVk458O/IVUadt/ou6aXGOEAylHKSMWn5iDOwVsl1/uipPlp4dU7pah
IkCRA2tNDun/26BeXKP5VrcElPp8dI7BIzXnnN3RWNgeBsowO4MXSlZilnBiOsoJxCssmQYGNepk
xeaECa1yDxc2MrCLk6B4LVRhr8/0MDkPnP7nsIv6GCn5bWu7/+H7EvfS7+HdI3TKieCel+nB3usV
a7u2orcMMOsZ13OW+5rW1J8PsSBLp6e94KeZidp0wrlUphu4B58ru8Yac5Ker2a6r4W4/q8PUKvM
18PzJssKF+Ze9ChT1/Y9kCjT66xsA4vRh8aeVxC8/PWQzdVY+QOThH6hy9IKLhF1HXdsdzVBy+lq
0PuDG0lfbl0Pya4kxm/f7nl3dQt15q25pIBnnZyB7CXZLprrXZ1ow51ZwAaV7UoCqhqLdOOmpyKX
Ss9Jwwmcs8Tl79eBmdDyMpGw0SdQ+En2YvNUd7AvvlPR11sr3RHSVmeEG6eymQL5euQGj/VE/BuU
WwAFHnfsoAHdjbNc84WAowntlnyOnRG692uMFfJR3xft8Q/umMGX/Stt7FKb8kW7sz1WNIUmfNZu
xV4NRf5Z0oX1XixydsTQBYXj61srQqcdJgr6wIlEr0mWMNl+8VehuvM7NLOhiOpO+t2IgvLkEkID
rCqCOzK/bfO0VyqMk32yknUUtMXoJcKfT/BPqtPHhQBAur0UO48OHxDjv394q4ihWyn3deTx510y
C7MgXKW8beGFBxKuJQqmQ0LcWiPPRcIRzsWx+RBl+VU/qH/yCGoRPLrhEHAAYFnFxMh9s8uaGGKh
dbncNOuJLbj3IB43u2mKHhw1FA0cs31bK1H6cHwB2HGO1aaSJWy+7rCFkAHhkxEyP4zQYtn0ULLh
jz7Zb8CW02+XQTJaiYtXwcDT//R3/xb40XZXS8vbsVC9qf2JdLcAyzuHUUAPc31BXxqp0ny6v2kK
9ERC495w1abbYaXXCzxn0iOSUUw4HNjYCwenwTBT+IkcPGsWT0YbLRk1d6T6clBmmPGaviOU+Xhr
L478sUjt8J4Jf4EAKsanaGR3pv1tEhmoYmuAGLm0d5wx6icach+K4Ks84rqc5H10a86ugzuyIuZN
E4bH066Djw1xzZCZNIg/5uybrLmyoXTFkzJxpO2GGbzh6hcKa37Rb2uil+MyTWCrerkqcyjLhf1S
lH6dmJUZZW6su052ebBaLjS+rTyGYy/I1RER/JfLL4lFv1TekBhPE19uow4g7ypHO3iiYxhFK7E8
d/zt5x9V7FDwsYhcTrALv1KkMjmPOnsS2ghTCsSqPYh/QxA5iiSp993F3sPEPCzm7i4ScRILcCPL
liulgYiGZsWYIczY/0m2GeeGRmB2dySyYXNzRSqwmPPpfkKb87/5GCbRcfqfCEEG567PqAH7YJTY
EC/eFuda0D8aF91BhuBzcCT5ymMCltWygb8DAH4B9Tp69xBfLo3kLdwdMhO7gG3K9KqONcymmG+2
GWBWOdU35wl7SR5dHk679/cSSaKM+iyBVwlXawEIMZWGUQsGGDLPpkmkXK0pnhGPmMT5keSY78ui
ezr7GWaZPWCZHOGMUYkdZX7imGFrGLQ7RT/2KfMu0u0a7BfM4IvlAJiX+lbI0U/DzMg8AAqjd5+5
IaYi86mzqQ43LPQ1M8icoLNhDvWqvv6UiH2hpfiQa1Y3Ji+wTIQ0cG4WvR5olMKIsxOYzmfIde2Q
8gZIs2pTc40r4tMDkf1muBobEvNRNBpQqxcBmjP9sP26p/6yBOTfxdE2PAKAr6aBi32fKB64xmbT
a3tOU/ix8C8Uzp57zr+uLqCrSOV6HBYNcwph5NI7+sz5qw33pTVeAWAVn3v2U842SZ6eBaVpF23Y
28kRy1eg+8c5N+qEX4CoFkmCQxRkNp4m2++LGOFTkWpKyjD2XPSr1zh1y5IIMei/Q4bcHjJz8aKQ
8yhyMluaYDZPYE5PPIcUDYpd2gbv17ThU6v2Wt/EkXSaBFg0VRfCIYfOoO+Kvn39CNpvOpm/aHUK
QywGj2MMvcrXFOXdo+yNvqcONaxIADWs3T49jM6BUCbqYT9ZJHP729hLBCGBFjzyn6Il8F7EpR4a
G+kYKUIT+CD9Du4KevIrEHPSMdvcOj+cMaxcKtsibahMAVBShbmyI9WwAaHiJ38WxpPBLsg9yQ+o
WtORDoK+s3HHcJzULZYzcw2u/XyddDulmZI8BUSmMRVsN+E5UaLN8U9mtZyvo7CZhqa8dtm3415x
SFW8Bo6Bj2IlpccU7q2TA6dKCOPWIdquidqQjeIf20wndxAuewn6xBVYNRpawbqoQuCpG2u+r/Qs
zt2uzrTdFHg6IoTVxq8Z6nG80Fqu1eUimNo+xZM04nPAmZaZ1eGavmEFPyS+iUG22SJWl0t/O3hw
oYpfaOvXPhcUOLirx+eGAT7HlWym7X0mEju5ToxCwhUhmDWpeMhErVgQlZLmU8nQuvqY7RtCMGNt
pz/CUwYR2ihyzylLDpsWnjHwwN7QJO/94JVvQFPdSjRnvylnoK8Z9cIZaJ/UVyxOhwx+v6tLO7/9
AJYfZOY3U94Xge7X7TZ1hnMyaLuN8DFldd4zg0GJb78bRHGTf8dFnmt3wvDNQap/frVIXEx+y+bA
/v9TF3m5aOzJbjKWroBi1YQu5AhKSs3s9oeBUtbboVtoxhwvOGtGWESX9fX27PHj3G3hKM+JvVum
+qcfMBWkEra4CptsvoTehGZgU5Uz9m0KkX4gbt2W+KYfnIRaYxb9BruVGa/wXdFQwBOfB961SLwg
txWHHHNFzacRvCJFdROq1Ivgpjlc9XJG6MaY4ypegE4DbOSbbZ7cswL3ZXTOFvym8L30h5at8NbI
4LOeLH3B0GRUNUlCXWhe3yFO/7W7mZv7rpVwprMAULS+RlDGd4l5a+V88GCxnEx3fEcske2PrzPM
QhAonbuvC5/yxIrmhZMDSJhYl7rgPNkkRt5efdQgG/ViiDKcFhQNRqThXE15beQ4wbeMa1hkGFtc
Zm6+9MuzSymDeg444qgpNIh88cbnQ+rzLz/EHlV2+jmV8qZvgjpEZhMbeDwmDRtFp7S+AAU2dPSV
7mjq4k0WB0otzDxPkIuJK2k0LEyIFAqJyOV7hx/IYXhqrUrXlQEdiZ4xSZUEG72pvAVj+DEVIqPN
o8bK41fVAV1Xouv/p9PT6dYWco41OrmRd7fxY7qiHieIH9vtr6hsMS/N/io+zxvuiZSUvSrMaChJ
3hIHvYUlGiNzmcRl/gTIhVynkMIqOLM/mQB9np0b9aaaaHFk5svN+umoAQ3z4bU6W1Vaqy80UnsX
xvK8njON1Bp4FHKwjGThA69REVF+SNxO/NpaRawDt/HecdKh18ghTgzR4ug7wuNZnOpnBAEjBDdB
NxHXbjifIkycDK6U/JHb4MNXs0OhfXqyhqkifZXp1s4DBLenloWYoJnZLIyRgL2eXsE/G/oJyLG+
X/6b7H+cvmsmgtw1BxzGdxoinYqM8xp20FocPhld6/aNaoizR8bIRY1CUDorAdeWDJdtjNIh8rW5
wzGObBDw3ndMiDzSu/SVDb/r6SGvDWQob/WzwfdXuRU5oCvlyKIuIUNWlGVQBcFlC/bZoAR94Siv
48P2TQIYkLMmEatzx3SeDZvZtD1l2JCE50qbEisLy9+X8DltpS/Eeujnka5i1SAqmkd5pKHbF6s/
D0y52+qTGp7AN4mOt6ncPm5AvoD3g8o1YSf3u9SRNSLmPhqN6oqCljPrcTzp1YNb9uMtumJMSxzA
nfpXZdHv6u5VlTVdhsyhyluGhfwvr1ele58jkRj32uuWNuSrixVgWT2B5CgosNFlN54CnvWFZSnh
dLSJSZk/k465gD3XE5D8wnA05vypfSyHOtlR3ElyP3blBDOVPWPfqhEYQQlVyFyMmFliir7QHkXi
3M23C2UZs/+nl+LKya6Z5K9XKu15gjjgfhvjA/tnB0QNqbobMsgr4+PS7iRSvdh3xnIjodotbOaI
0ha06RbFY3QwZ+i2hsfPZ3aQ/JsjPcUVmTLKi5y9NmV2V6cCERheNsen+8eXNTdKHf+nJj4LRhRT
Jr0zDMQxYPH94i9+NWhqdd/0faMWtR0jeGmIBlqZCOr0Kd4eI/9oIdT6freZJYyWbDPqumorsfTv
2iSZcrhDCE3K7CT1DBQXYVX0Q/CxNdREByfOzEzxvzF4WYbCGbWWVjtLjKYbksZpDhlc+kv9q5p3
iqZ5oklquspAutQ7ebRQGQ6uDTMSN5j7OtW4gHkc8AZf4MsWzKopyvrBSqqI+3qDK3Xyo4mDDrMP
McskhImjXkwG+kHqAmnq4we9z1eIdVmx2eSvwsXz7WlI5To7CccTZDkOOESbuztU5sRVCTp7H3c7
X3f55LQ8M+fA9ZNkUP7dozYBp8mqWYzK0cSm/2ItQSxbEtTVdU7x59SBMtkuUIes0s6H6GyslwY6
YriGRa78q09eYIjDdSWq85MXvOFqa5h5tIqE1HUPJc3fmkWNPLbcPnfFk0SR8yRh+aEQ/C0ysXHr
J+D/eJJOgF/4gaRCutav0KYM7EQp/UbIw0aD4pWHCZfYsdx5OP/N2mq43REQwH1wF6Uex5IffB1Y
b5WFzakuk6AIJczHvLsRop82t50knq1G87Hu/DfbXMdr0xQMhXL0b038oXvOlznFu0Y+LFeJSTJ6
DgGqdigakEFKJ6XGRn6RBVJyjG2CWkocP5O8G2EUZ1Hh4d+N/2rc4RnBmhvQssKp5W4l4ELJgH7V
Nq/mKAQ/1J0DhI2RfgSAeii7asRcsd6KPInp8OI8gb11pvSfFPgb2Zvlc8qf55y51rWk2mpz1d2A
CcbBYKNDSCuEvIXK+ZbDPchToPGisyq0GkRYs6bxGv0uDvGBKAA8lFX122CCsq8LAtCuRsrOU0nE
Y7awCfYpoVdnkMNDuCduqJ95VvXoRYdXkeIJ8SseRkogNEV5HGuGujxnNyP9pYF7fOgY1/9ZxBrK
kR5VWieJ+X7KiW74uRUQwhB+oYgnN2aXzugMSlM+7Rf4JBvrrZbsPcpqQ/XXDjj6NlJVPA10ukt0
5qZr9erHlPuwwaIY5DrHITZtV147UHbaTtdYwxA8eqJknGw+K/EbLfr8cQA6m4qFDEPl2SdBZrFA
gRlrEjCz1BuC7Ukjsh3a+Bi3czoB48Ry2W/g3ppcd5OSAFl/Ai8Er4+ycNHInp0ZlwHg6p5UgeNR
iYelnpLZ6Z1o0S67qNeRv2nyA/nmj8CFvIQQPCIUVk1Lc3qLFyIOACV5Nm8ltCj1A4iIXNPlXTFt
sI7U4GntiDfjjZX74unTO0Yo3sqrIjxTyydTvcW1Sk4KsMWkYZza5X0GE4LXmhnoCurKoG2JHC3I
t9bhIpskIbUq6XjFD0VGx156e1TVCwTaycWcGQ7uB2Z+JHzpeWgP5+b/tV2uH+VJUDT+aI+bCzjZ
LgwuehTftx0q0pwV9l2un7uPbNEJ462FZJkxMe4x4U67nY5r5vq9lkVr83cPDD0OZ3Xwj+AsMYEA
aCleVYjNopKTaFp/r3Ldtkutz+MVZoSF7RLB7FKIE4npt7RB6r1I6j8v5pXnBKOQlT4aO4vt8pRd
Ht/jORN6vMsSv+4aDktQrg+tJ6PgkB2x3NQxRe0BkUnVZD3IYUgu3XaVgbActPrZuHLTLTsolkzw
O3sxV4ZJ90HbbFk7JquQtt+kiH2L0TqeIJxLj8pJoHosZjqYIs3x1gGM7J2LFkOq5ls00r1QMWBb
Wmnq2KkeUwwIKez13cdFd7fLILr7QAqJdPYRIptNuXfghp1lkrz2SAxf0OECB0tQRuR0S0Lq63Uu
Ub3BIDcpsUcG6bW4Lr/DPnC1FYEgEfb6F3GnKNt66dCV30yY/XCZQsQEyL1msk6KxL4/CAcx9WrT
sZFASlwUv5qR2F21GYrqy8E/UzVPoxOW7JWwokk5JiUES0nw16qPauesdszVVqrQzETp6YRTylpX
o+i2pv/U6+2nZ4XkYovrk6Ufowtb9pRw5WCw8uETAM8kUV6C99282Mk8fxtl3aS2m80nnb92Me1P
wju0TI60elN8Z7hJUcoRyGY6xmlCcm7OU6vZxoGHV8WyWxsERl0F1IF8+c7cSytJhiVj1NNlqO7z
ponq5iEjIdpYzWaD9GEkL4i4PdzdOSXm1A3GiJqsuvbqdst9c8xfbg2DilcQobI/PV6kZSjhQTX0
ZgEQWyojPHe+fM1VQ+iW/0GOYDsA6vfrmFSG9+xcRQIeXUYpyYRsSItRiUQoduiOAnB7Ir7Hxt2m
R8y8WE5PaPlyF8VtiJcFo12Vw66DGOZlMWh+yPW+uaI7bXoc0nVJZDYaF3fXo8y1C0lltjIBDTSh
gFeYmyapsmj1xgDyWDYTZMDeMQ0YRWV4h5XQEYhBPhM9DfuelCZieyxUsqv25lM1y83B1YkbKp5d
DEUJlssxgTEZdbp9oBDAlARLgJoywZ2/NlJDUa44LtpLp/ovEtzl1RxvLM6OX+VwhPojjarSx00+
7nGHmu/gn/BeK6J8pDgR1s2982HI43B2FLLGVFlSbTySWaSfxorRiNkRpJtFkOCa8NolTFZltjsC
YrUU+yizZZowAn0W/Uu1QLf7qtOkvlbRuYyK673WkTBzb73FhO2TAiMlJ5hOHSd5NZ1EtaVebusQ
ObzYD93wySDLBH/rt8bFhJ4kOXdgGf43aXv4LdDnfoCA8cNnypfvoigN4HSBPOAhTMUBD0yd442g
F9B9qGeJfp2+kS0F7NeffP4rmsXmHIirz6xDmE2Z3qFHsWEw/dcuMcgHnpuXna1Q6wwppSr5kHGQ
odVL48PHWS6e12LF6mlss+ogfibXqG+mNyNpA2vzcHx+NQDM9/E2WwH1mBB3FMQAh3e1sfcgEPJv
sRHUAJ7imnKdGMVtb1q+2l1pjUujD0/KRhL3fQZEjHu8CbxzBOIuvfpyQPrF720SUgOAg/d12G/p
I51M3IbTDNQmu/h9Y76XhNgw1Ve059H6AGfhmAtntUAFTEdJsqLpulZ0es/Ag3y66BIFtOVaKclJ
1oOfCQ26RL4qHXym8QMiK8cLP8iIA0RB4PFUEQDBfTSaUcp+bTOMykHy1TDUqMtd0Y96okLXPvY3
M5w59AMArd5SPcHAs0owsquVJ9HKgABaLVWOAuyPJt1vJx4hURZoEXlyf7FocZW6QtsvsA7+toAL
6hB6BXZ0UOfGEpnWPCatBWd3cf3La/su9YbUWzXNOfTxV0DFwrzeCV8NyBoad2aHdqoQ0pkTykY6
QvHsFeVI+wRprMAE5CSY0eLnZrOk/6fMcmZC7qc8+uu3oUF0l297ItKwJ4lNaZf05fpp+XI5P1xU
4/OvqyrMTModCzWlS/1vg/L4tWHCaSrDhfeBPEpVnrlsMrjc1+G78ZxdHggAoLJBPL1WlXKyL7Hc
hqL1zlaNHP3jSHWY8Wl77hkybsCx482ezdZ9CtUgNK1nlsxqTCN+By+AFI9W04RDyc6HBUUsjWtz
Ovpf7kYsEDmfdy4i5fDoiKwuuiYDWx77H3gZ4Dha84BBp3EJqATLwUhlLcYKQe7MEfwighXKmYAU
5kyWslLRh3cuBqfvREj7UKcEnL86bailIs3v1dcPtPjsHsk+CisrGB6/2vpFOHy0G/W7kHe211bS
qhNWoSTHlmkQqQ+GfzssQAC6wNL9/mkeffdGVnylDJBF3PIG2A2HolzP7dUAdTrUP4mX5MbiUbC3
DiuQYV7BLZybTSUNRK6d2seLlA0dbeL2Znquokud48LmSIKja5/lzsB+2RpuaZdWbKFLupMYKwyx
g14yX4lrAJmMGbocD+35WizyHj7+fKGf5l1+IyQf+wOisreGy1jfti09q4FzfbRQUCrQcxi/rayV
T6gWIvxPHzWs8DDOaxezXDGMwbS7r+rNA9uCrOFEZoFymDjIhEIMmDmyd02hcQW/62WMoGpkzMr2
4OwslJ0iVJe40oN5MpvHzk/dorFPE/CSyh8iamfLrg0YdpMlHFXWsaSYON3/fvU7lz3xLurnTrFL
ACCR2VaTXigcJB4b42yRbUyBNbWLtSnHDvXGIi1t+tlB38O4bOH1CNUOXHUlwWwUXAVbClJz4ecI
aK/e6Vm+rD/S7wjG+cYlqVvClBOIltAHbN5mKEV/OkKFJrrP+Gm7q3pahlpRg4LyAF+MzLkrCBUn
dgxAjWEfjoqNpJL1IprDS9tLYacW50mmFCHtdUG2Dd16IemxNStM/I+5W31/uiDQ8JMSAHLHVdf8
+zDrADRcnJNEPARH5u/Nu/6aAeugqHSXNknmAKIm+upVMt9PMQhL8+DHZsgUSfDz1J0c3npv1tdN
+UcU1QclD/rSO9LzGj9nlXdEFYajxk/VFDm9GZG6384v0g1Ct3yxQTZV4ZfOZdla5N3eF/tIMzq2
+o779KVxJkONk7vU/F5FzGXqihKN0HPiyYwuSGOU2IaAFSF85CFvlodTy/vJNfXaFD4/E+ZpSFuJ
QwtSS/+uCE97vxpSzXvAnh+XrbJCcz7UnpcnB/exiLQb2mOYgRWQRy4AKFE6pQGpdOUbrrhuTvHw
d3MmY2AuxXl9fouh9LyuTlg3GDQ4WHxdKqRsSKFA4Oa36YoFzk7Bc8k/m7GLZpN/hlIcUkjGQBeI
Hw3qRDPzmqB6eJCQ5UWrceKHlWd569Sf7ZrjEjRdoMT+t8wnxRA79ei39uPgNsDO8cRs/yQYbr6q
ur/ya1/lsEQ1RAkkFwGm0w5ehwh0yNmVdLzUtmhDGSTC3vQJb8MHnxjYOOqwTxswM2FjEaCPHimM
F/OktR1TSh/IYLnMSI8xClCWd6sWONbNOiWpNT7FyFDuQuXCKj7kGxEmdcWJyqMsiTOxt4KEYV1w
qosYRUbo72O43x7VVCTJesjhtI9yUOoAuGMg2D/ID80MYSu3O44U0UYbkX5/a5njBYlegmdVRR3S
GP5NJcH9Qwr42pg1rFGsY47o4x5Ovz4EZdYMUoMw1HnndW55ncVdGdDl/PT959pqVIyqx6+4gSai
WMtNpK9QayZA4qdEeVosrLJ50cblCBIuq3cyccuNTIvUOYby+siO9aKGCxQarx3/Z5TJn29qq2MB
sGUHyCw/6lnkVoX+5E869SZ28JjFsD5E1v/Ive6xmkTvHBeT/RVz7cYha/k1thsmqqNZi8CF2n7x
cvKuJQODcXp7pX+FgWinSmsyx6TPVm3iI5kIGfzCElmDcf/862OHXz+CkvQfdDltlCbY4kHEA5rY
tZl5gXIZllAz6nAPdKIab76jaCzGwRKjpXeorJH/QKsvu7dkNUup5JYUU75ETMf76gA9e4Yia2sL
/G4JmLGNCNGW1MW3wYHcjq5JkvMi9aWza/uXU7GVcJzD4mD+CSBvgDbEjzhUV+Xq7KSkfe43Rn01
+DoYxgmufBBZH0yJlr55oWOX8f9Efi3fibZYWf2WG450+Ro28U8ij3UXb/mhS9XICgzvfXvLdZAd
H2+utlxru1FsJT8jwv82ic4rwXCzRiJU+U05W6mfnsbmkKfAMpuTClR53aTt8piGNvkJItFopKPq
sgqrWC2Y0Rwq5e9OSAJ4SVDIXZoUkj77scLwFok6gVax9xtgen3l/r+3QzBWMkSEJgjL17BXWIbw
lzJhEfoDZcVTOK59FcEZqtgDkd3m+A/Di02WpazIuP0GENt8cH+xep/CA2JZQNM1/4NVqICtV2qg
teaejuw2ahkLIUjl01Y7cIj7gkndRIYdgBCdEJ30rPYQK1dGK0ee7rhcyrTgxdU12cqLGifg50NN
cEJSxtz+2mib8L29ywNrSLsNBSzbh4+Sr+ToFvyLgRrVZZQbtRPVsY9iO+T7yCaQgpWnPdHAymDt
k9taYjqLSygyNsCoqBkR2a069kq4hVKxMVO08Rk7AWjCQt5s5Dnq8Zuek+wRwwRWfy10wBi2+FyA
4oRP70Oq3JDFgzt1sgiv1n4aE5E+IltFSCGgKyiYSYmi/F6sVd0rscNgOROoCmeNmTdUgV7yDrUW
cI+Xc+LBmZewQDq/uhK+Zi8pZ3ZcAHNTwrlSrNYqdPPv5dSw66AkqcqJRhwQzmuY1zHnAXgGyxY3
eZ5D9oj4JsUds4Jtgwfl08XeS4A4OAdDkNffuLAMkC57RKgfE/Vc6eEcaaWltsT2QQcgLzGRPJzp
WqfbYWtYZHc2WwbehIpdubpyrl6QzOPEIrmlq9uiE2ZnCAI63OePqdYK01q1DV16DHKAQvzMjybW
OmAnOYhMZjLCLsGqky+kPtmzMmsQuI8vRpZqhZkBrvM43qIP/ZzAm2Jb6WCa2ruMG3tPNcSe98M9
MRyQucDlhjseg/o04tfe5ulKS3/B35sQYYY+fBbKyH2iULmpnXe9HcNSLuclCH6osqx64N8r2Q3C
nCb+CUCubxI1K1WFZF1vICMfRxry2IJp+QeSSBhGDxjg+lUmphIMUVlg8Bn+S9jKNIkJgEKA10Du
DKZGHO6OEA11ajgr2jlY9HHy+sk6VijiaxevrNYiUytAhHh0fM/+r1lgHtwL1VNa8l15DzrzkR53
sjryOcH1PBurqxTzohenKt/kr96pR1K/t3yDV1rZVYlRrBNZd3KVeLsY7iGPUvmvjR7O0yeF918i
yYqeqQ4QeMitN80ltmHyWvMk7opxcGtJjAB3j8EuYh1hJu+6FyDloG4h/7kF7nH2JCh6fUruFs3d
fkVaCkUb1gjL2JwobLd4u7xFhNW2Msj0s914diQ+zAnzrQNNRZscLov+iM6UVzFvAKPzalPMn+jR
kcvWLdCp6eaIOmTTuYdhpipWtnnuZoPasRdrEPm4B/FEb7NhuTJttCDgce24vj1CZkMFddl4YuV/
2H0lk4AvGmTDSoXCufUSuoZHHcdDBQHGK46abroJ0JcqbZWZEwOaLF8W0KyteZ44VUeFUSKVOEhw
ANNlyKR9+HzbNj/saG0PF6tzk6dncVYWFV/f4MRDRW1PsNJY2lcrPxlAeDVVbNE/Y62TS08VuiCS
NReijvwu4DJH11XhE0coys3NXreWGf1ehEW1nBlKR/tJIdJrEn4JdGagEuB23i0M8S8OpGOrXC1/
Zh9Jsr9seBmqeapbtBFoTmaEpR54yczOa0PzCyIzr0VvvKBLGN2gjQQ75wzxc+mLUnFYA3ynL0DN
cDyM/hU27QNae2CFyBLKAHnkbv6d5wJNG6QbcKSWiC1PNgFAdwoC9QiDdWQ26u5AqsmV9ypOSJZT
DFiriX4PzCfcz0qO070CItav3ipK/DjUNPrfM7afcGQY6/SN3yPEkrRQUICr2skC929zdZcE+m0J
6tUmeEPnugTmx+qVbfDpdfSDirF7W6EvYVeboXlHB4J716fmKx7DAzYkDzmu3AKKAGRUIbxPxyaW
1l7avHk9ShLoXPESgfRFh2mfQg/ciEuct22PZOhG76KwoiAZ6h5059bLOLqM2C96RWJI+pLeW8aQ
dp2GCE5TS9FCuZK32g8OcxZiPV4AsbzI6l9JhRYVVHqEq2XMPAhu3KKBL2uHysAsl1Rj2nHOatli
W2uxArEkBWzt+l9Fu4QO6Y3eMcZg4KvOc+6GDrgzbClkFsuV4wHLxc+W6OUDM6sByPY2F4c9MtjF
7pjmWavK0lrcymeT4VvAPcLo6rpNbLS4QiqOi8UnLVCs7G1ATLaiJN/QeMK3XNjkgz2dRisK1qX3
ySj0mectcc5tb18TceizOtIGc5ODj2JviyIy3WLGUSofAYA+6SLfqndRWLqli5pGo8QJcSlzEoH9
Yr1A0gXiHmZXFiPrPRN5ViE+oAvVF2TMmU6ddBkvJbZWD6hoVrCy7bYjlc+vjTzxsDmrbrbxiZC+
CwJQe/bWLvfsjEdN9zDq/K28EhYzIpssn8A0e8vSBZAuF2RD5PEiCOhyA1LYOo8kjGvsLTmipueV
k16KAZ2W9ssNQT5ic/A1fVdjh811f5l311y4C0UTFLH5ZlWY+3W3Qrj/ZlmHdS9bo46M4celzw/h
ay8s8eR6guFllI1bP2HQ3KqvTfK7bXTEm2KvcEHYDZ/5Ff8i7sKDZwJbcnPKUpqQy31i8Q8CuFfI
Q7HP8+bOTkPdInxj8Ts7a5VMdarASgEXlRqMyGngVqV5rVo5g2KPr9LoWxqQBbkAgrnn4l0lwuup
X8G3Rilj3WO3lRDviR9/eXeYDvr/9wh9HDjcnmafCyFXy5HWRrzjiLxLo7+Hk20keYRAYNIxCXHW
KA1ZYZKdMJQa42qWy4ONTHn1jeVusxCWtPsXliFuSRMHUynEh8eDrBh6nuRPs7fFUTd1y1W/WyXu
zRC8YTUdwggWXePw78+BiDSbzXhFWmKPNB2MvLq4OBuRj51Z0lVU32xnQ4+HZg4jl4ASiKh89HFt
J6m7d1yxJC/oYitgHsDPd4TqagkxUKzUYUjA6NX7nJtWrLCbKmSe9fVJQA1zEibVXxIAvc+enaOH
LYadK+GL4f/CdwvuKLEiW3auQt+mk8d9Ha3baks9vLe3Uh+ZFGjxMl+HHrsqJcPnV8qk9xMe35IC
O6jSLphC+d5BuiJf8X8r1MA6kk04LOaskupt9mZpGPztFlMAXp32QT+YJ6KLzKzpuUV5SfdP2kPr
k/uFfIMtTYlcmcpi2qEqwyVBg7AUKyN2PD5XjL49tcVlKVjJRXLoV2SGEX0Xv3+fT9fpVfDFluMF
XT+rew2XXi+jfwBnM8XSRgrpxE+aTL5dDEYK5V3T3ZGD4+uYzpIgWLI++eqRLmeQbWwTCznojCgj
0IbPNE2EmPEPj8vQ45BjCn/k+SZohEWj0wbBDfsN2mzgRU1cqVrvgdHsgk7r9ZCl8Y6rDrNk2dXd
OctlvUqEMvDt5uevtX9cwboSlXJ1+zxlUDGZDeELkVrMzDr8gDjcWqf4Bskjdp2I29xwi9o+dLyy
6LJMf74t9/2IggYX26zN7VvA6mWLbus0wGKW+I/XDyCEpXe80jlJxb72WSW79ADaqWCP5x5VF0N4
he7awAQySQCD2ZyTB99nhtQ1jIQxW2f+hvdOoV2xhCvrLeCcqLjdWXyZhwzPgbBixlNQ6olROmV9
9JL3uB/WqE74QtNdMT7rtExxBaY6+GZDYpEwSNdOSJsvvjeOT+bPZdsAzm461056kIqubPP3cawU
3NJshpG3KXZZD87UpxE2xM5VSJJ9e3DtntL5tDz0viaWlne5sysxN1xWMluss9UPtxJFRwJYgSdW
wIphl3vGSEPu2ocH25VhBnJbE75UH7KfS+9ucWZwX8rcxfOaZCyKdPeHmF5I/8QYzt0z/V2TQg20
7IxTLoz79KukZBxB9y7ULTfRUMeA5o3iT9n2KIZCTSfPncQ8josndmPLCyNHkbBQXPYRZZpwi3Ln
XS19Eagtjd+OiHMlNprRotWI129o4tkNiKRzRgPGk8fDHUifxp8ST+UQ2I/fQqHCmfFMFX/0Whs8
+xUKLC/JpWZ2ulaBV5djL7Acg4MX5FZlfdfrongy8mhGUa1syPWwICtEM09HfVTSA3IWHmltd3sl
VFc1nwdI0+EWdFodNa01/7g+OMcNrIDmlksQSjVxEgZXN1Z+iiiFHnH/ipWgumIaURnZxb7OLGVh
OxgkruvM43bQBFH6oW5KuvEpiQWNrQkO8SYeSbdIjAeQrc+K9NCihI6JHSf1lTMus9oewF4hqB9p
nn0ZfjgBiajqTfL+x0rPK40yWWGlB7vz75ntQniP+RgMiR2j1yaWHeTwu8sgZRVTh7VHTmq7D1Fm
ZFoYgZOVx+ABAGVho2OnRx3nZ4zOqkkymet521Et9phUaP4x9nol5iIbnZqAE0nB9aCz+g7zNGF3
vZFCgzKGkfdwI5jnZXEvRQsKijWSDKawon9UuNCH+sY7SosNAFRG2NJa/Ae9c+zNJG1xRRQba+fX
gExkElWnQwGk7aBHvURmQU74La26sXQpsGecZMzTY6+oCKnTVBMUcQ79V2P8lGJ1TGBjowF3EvIb
I65PMjXfU0UtTTdx84G4FplcjN8F6urMwJ85UXHmUG3SKaGoEyrliykKzpiQceUXCPXA3KikPww8
CScUFOU0U2xgNtd97HGmE+E4vyq9zfTNcXB8jhh1ThD8dJ9FnppYw/q1indZ/iDk0nuNAbCBZreQ
Ue9nf7cCiR9o/xv54j7IKfeNeOTdGBANxb5dRomuguCLAcOR7gXXa54x8i6fQYX+gD+QlNTLcIYS
pS3Gfy9eayULyHOFFs8FC1dW55gKKfqVZdZE6RWtgSzFqkRDwf8G72ow+3Dgik5/aW5Yr+U4p9+7
KV1t+bluricICsc9Hgy4+XaotdBad7aVFCf/esbNQTPZejOYkU/YuaX/9kMAjsEm+iQ7yltTR1Jz
cTsBhUhgaxZDzm2IkBSI+AmxnQLniUug6FqI2tw+dW7jzzMaIgD2n/OSwe3EJbxSWDd7yjRjw4Pw
8CA0KWJ1Pzla9brbY8ls51kmCPImxKPD7qFYq7h931iP7MsyGoIWZIFDFgi2wT2D4MF0jaDiQ563
nyt12CQ5vLME8oxDa3dPEOeb6ai0D6LyDA0NyQBkWRJSe0bY/3XAqi2QTvBNEO703kHTkMO5nsxt
puAidD21VzS28X2ArQnSwuCkX0JYCpCHoLzC/SeQ2BtTpefWUOI7PaOH/3FUDROmbiWPC05A5GU+
6dOCDpEqNSvE/06t5XWkA4Q1esKXVtqem5FXFnbl4sy5sm+zkeiuuu4KvUR74ktpSqfDAWrxRYOC
zEIvi9THjkLfnO/3zuN9mz6rUIgfq+w48jcpo7UQaAb++2C3fq5K7MLJzjxFenVvcT6CEW05uvuR
TSKIp3D6+yLxWizXc2+Tgo5eJRCqnXnE5DKQuylsCeiJu+zvdTf1e7nbrtByv4Bc7LYXhzE8QQ5V
Zn80PyexT1vhfg3qhFuiYTKSYxJ+lRNQnWIG3C+F5KX83ZAIfpf995RuEMOuO2ron/cfxpNugYY4
akv8DckqcLdCpzmorwfrl7XsCCGtq1mGpuHPe1G3OHP4opbb0CR7oDWC5cDHT3yEr5uW62GRuSsz
ezdfJTyPcxnE3I1M/3dUvI+FRhe6NBSnwiWWc4jQrx0rC9rIxLcyWB7Y8KdEBewXGNoKd9zqPLmL
KhfKQ6RKWoNFtvig2f7JcFs4sC08zMDTyT0zVSR5J0evKd5MZcv8E8R2o2lZMAAxSx2r5U4pCTfj
duE9sOD/BYztr15s0EBkP5FyDo8////EOXcQs6FhiQpJ8pccKNjJ/WpNk0BO2WlGhxBurBI2tJWi
7JLNOfR6Q03CocxM1c8M9vRfkVNNhh87beJjfNiqhREHKjigMVL6pwZiIFZ5vX/JJpoanr1q/CjB
BJwBMeZgagVnBWrQtbtsQ69FLAxBRMFzYpR3+PLf1fg+8Pa/p2tXvWnGevzUTkaq3r8MGS/CA1Zv
uRT6H3xLa4AUk7g5A6H9Xm2jDEF+XCQbxELUpW4fiixL7k+YxPJ8shANrCA+qDCmzk/CZ8zrx9mg
XigdSK4jL2n+WX9vfSzs//d4fb2G8MapNGX9EVT6fMmRg1EaF+cC5vfQq/l25lYryiNvwizJsYVg
Z6YFQpzpsb/hftppAnQBbrYna7IEMeZIxA74ez9b8QM8/Is44Vp87cYKzhWyiJmVGdhHYSbghZC/
F/NfqXFLzQov0hKxnaC6HnJD+4IuGqPp7+oArKY0hNuCGexKaCIjhAN/6uvSWiv/E8F3gmORjMZl
QRVIqBotzRO0Bg1OC5fFtJTyBKR4oXa1Fk0gwyxXcvCIQr2U3L8ITGHQP4061/IThCKLqM+sHLF7
25eeutdy0sQckqPq69HTeP49iIJLAFW1AOvNTHDs46P9uifWCEQ9qNijxZb+3SESKB2gE2CnZdzc
qAecCCfwGVjCkC5gEfQvhkENTFUozrz8TeiX7DGy1tM81PJQsfHk5lXNwXe2V0ewh4BCldirmXeh
iQb3vmKcAm12AkqhfMS9r5cWFuVO4ur/K9zrtnkpcvIW9eWhvFWZXhNnPC42NROEzB5yyyz9iaUp
FWCuXPPaSZPgnA7uvEFeYSd6bPWSYz/LC6KeP6/Bnh8CHspQjFly+x6hKP8qAK5y17hzn4VRbe8r
Rpfc6XgZmE4mdv2dC58Y+UreodPTMNuMKIESyIZBrmZ6XrJBrme2oE3/mLxEOSiMToJIfcIZn+1l
mEVtIM/YhYREbJx26mLZkZL3gN0syjUCRz+h1sl8iJGog0mCxcqvVzIV3PytmseTW5tlVxjlWh4j
WA7HwybcZ0+0Ir0IS9Y8BBbaqSP26XrmRt5pSIoH2RPzMZ7Da05d8OfLZ/Wnppi1iv4ThXyAyYSE
F14t3Sjkff3VpIEylunlPpb0VNifQD8FeuYM/aecPiv2zl12nVcogMGMDtVoAq6pfEABCsQBv51a
lLtKlRO+8lzbfkwj05mbf/K2KDkZoqCZ5kgcdP8WVsE7sopI+WQExQoLSPNiiQb87zMGyvIzLQiL
ZpjvRZc86iDWEDGlsc3xo335b2t/Vp0XRdS5XEopKTkkxXFMu6vUt95q8gVMQ9EXtM0ZlkrNzBIV
TgitojyCluoxiWUmiaBbBhHn+177dhNX0BB22nzUMXY/mkNBtI6n6kbWDRR3sJXUQdgGbTY24R5V
oypd7q4ZzHkNw5Gyo2HUTbRaYuDL43Bfj2YeZG5kP8FaZQh5gtYz2WnTRhSF++ojdP9GNAAQLDo5
yK6IPMy/OrZSMUaiSZLzrE6LNcLYU7YjAA/4ktTtpigAlQr4oYm5d/w4TNjaCFVFkiYPhqP0M+gQ
MR6BX95cVD5r5AEgpfDBUo2WuIJm7bP88vMFKCeuG5kO1u3Vhu/oDg20Iejyscm4ps3FSga1r1jQ
IY3v6LNejO/1lR2DMFIgwIwTzVnQ83Sz3NUrOSMZeGK0pLwSb9vrgevt9x9wkKl2HegvsMbBxRjU
TTUFx8Yno+lWmDaVF2DNM+zj5dtCyA0QVuoHwfmMFTTR0jFYbZziQRhqCEgOD05WdrQG1not0Ul0
jTHO+1N/9YuL9zWm3fYVtyJQiPsLkCzHeNUDTAboALBkqM5Z5C1d/s+s0Hvu+4PdRjJD0gifrGnb
sX8rzB3DCv043wLjD6P70+6J/Wot9JX9mTwo58Sg+YoNUFYZX9tX7137aszc4sA64VUw+NiEvTfF
1ol100uKG4eYLQdNKSHcokjzRXxnyXRrrq9GzyhxSLLL7MPdqms4jh2WTCDlaWHG0xL6GYGKbXkr
CaufA556KKZX0dnv5/mPFoQZ8nd1djsC0ZC0MCb+QbwAot0Zm8jcu+5Mj3rw3y0wKWMLAkga9nFH
ge2hJLDn5E/2WSEIKE7+9Qwte0z2mYDjulGtg4taZew+skFvkD8lEn6Hm/ndsxMcdaDFBzRHfCNZ
tpbX3rCpV9pfl7pFlLncnZBgfnUoe1pZuSnz8l5TPPjYr0dx7xHvkPEqis1T4ou3MPN191qkpG3N
t9bxIo6s+mbeOWrWKRcZ0/6f/iXDmOxqo7Hjp/q/Oaz2yB2YF/YMRKFZ597bEQP0L241k3BsvqTJ
g+V4tq+g3IOTlx1INFWovksK7493Fg+2a6kVbHA/bpRSIWwzmfO5UKLsjJcZJQgJATPxRtCv+sF+
um2GgWK6s8TEmkafNMRTNG8ajUqEAkEVHZUSRlryNNhdVitXvB/kCj4phkGYlB2cyGoFnxwZxydo
HVvYrOTATOPebKxsPLx4NwOfpFqC8sCXHQFrHT/KeGisOAf29EK25NsGySVpxKwxfU0wKulgw1dT
WxUr/GRPjbDhxbM2YprDk0sichH3Dox2pV1/EDU5gh1ft1xl9UEwCpnajnoGAO6gP/ZaHkT/dxMM
Pp+HqVw9MoZ9EudPDbrP9EVFVcCKfH/pGRARNdeEaCuIIV0N/bm7xmDRuV/bwGYbVnrWq1mlgVXZ
hqsgVcOTulu9d2dJxrZ1QVM6Hqg+JY8dH0Xl8Ff27ojljfylxw/6Rj6ys9bpA+QiZE27rgeE4GeI
G4RWBFvQjAev6sCwgmEoDZvHXG6OMx6ZmWCHOMVwxjMigzcwttEUWuy5ZCargSOo/04Mb+E7kPrY
j44uACaere8y9tCxu+DYRQO6ggaQ7nVuHBT3pfr11spzJLXwPcVkWND30QTcmCS3/62JbOuipjMW
G/l+04hUJ2cFW79QE5Qw7xK3cENuGeEGPvUHI9kJ797r4uC4Ib+raSkIgSivIWyOms8Q3bjGIq66
Phknkrpnyy/zMB85C8Kd5B9W+pxlOmk1qRTT3cndG5KHXsnOZ6RhYpL+OHCiJNfpacjPENqHFUoe
RCTe251GcsqyA8NAlIKcSsdZgWYAn9+AbUE5yZGWb3dMqgoLiC5wEdwAvqJ1zsNjTXloXSqxUdMV
wnwRd4IrQprfWpsXhL06Yv8OepMo8B+uba2dPMdNSWFaRgnQtrgKIH8xgMOLc3tG3r2+/ePZ1h/W
reTg2sS9EjIUPDfAEPOWa4TwzFsJqexvhbPHKI4iel4jyh3NbHMlyEyMxDA20I1Vd4+lQ7yOFFuK
i53BvbXuS31PN6R69LdD9IWrq7wHq9SiBC/jEqeT/omsWE/X9Fvvub+vZw4GS9q67DPzYyQdc3R4
6yr8feAgp9I5PxZZSJQdWEBxBDbYPOot7GPiHE2BX6SXXtZnM1N74TcBe8yCyhfuWlkbLv6CjVWu
uvFT30uSbXybE44YdE/gqAV038YPI135xibP+yHAh7NBhmF10aLFtP2G150wMaJcXy5MXrZmyIl3
3pKKK9juLlx9JhLtCBS6qdwYUhmE4u3l8jFsYTiLUurITMvukpX31TFUN3P5GRt1gD1cbRzmaq6I
4hTv77b/tEOSTPioxOkIGse3vKPqT7sDLVhyftY2O0gPPQyX2qYzcUWl5uieqgWqPBOZ5UX/CXxS
oouYsYBDb9M1XXSkkw8gNnrBojmjigsM6BdQ54JEvVG/8IBeiS0SG1RyWoJyIuHN65P4tDODWAZf
9GwYRNS8bPpheifeGUCvKedlXQJszczoYJoPCwyfXW7NvFeHRqb0QQwz6OOkcAi96MDF0M+lMojx
+tGnQZU7zUAdwt5cg8eqZWS7JIebjdEcYqw0eYHvNxicYN3H1aXHEacDmFzDiFVIKClWsXYbxwLO
XUvbIgFLkNkf73E08KH5zn2C1t2hjOoY/zKlgzMN317TLW69K79u2cAQ6V2ot0kmQJg9FWEUZKm3
3tpL8ktrbSGRJ4VkxV83GyIC4eBFXTKZBiKU2TNn22eOCqAzVKxz6ndGN12/dHTTVXudvyOSySNP
OzWrSeE8jhIKA42tWAnLcowNAtbpzcmuBElpTMzZX8e2+MGRv3tNHex+sq3IiauMMJ7upHQu7Gl3
F3a+aDjkBVIAbg2n7tv7LD4+XDaMUlgq7PVrvIpG1wRJ7art6el1Dpevy/QFFMd52f7p665Jx7Na
kDxWb5JW9DcSzQXYTflNdts7Mf7TYmf2dfvrvzBbr0LFWPI6xFNnimi0PKwX0JTb3S889CbTcNEk
C4ABFRVszegY6930C4/7hcAzSmC+PoJmLHtCy+DJ/KLvmw8479L1uVH2KMQYYY84Kt14Pfc22fVM
1dxqzSZuoUGtKdFx27HgiclgN+stBjKgHZnNfu4py2dXJJWn/YZMG5gLSIRZrlPeb5QeSTu5mI8/
pXFZONIg3xEuZi2cnKVQap7AWzYJIJXo70mCYaqT1JHjOT2ihslALxVluPatm5j58VfwkV+vGE8/
wsIfrvJectF4S+rGwtEe+EJQb/KUvmiuKbSWbUHq1Raiy+/dq1CG8d/CA9o1Cfy+F5IdCJCVQ5jz
rzTs+8gJKdt1ixp90+inQ0KasrejdJuO8dSxmJSc8c55WpWOGscJaeK8Yg/r/+ZyIhWpCDY3nZg2
iejpzDwBGgDffbEAZ4D92EEBtaTaP5Ehs6KoMDA2dbwalk6KkVpZrz/Xq7GtH1D79Z8Yvbi+VJeg
179wts3qeKQWMpC7E/MMAEKetwQ+TDqZw7DaVUFQ/xiJyuCY1dCu/QvSLAgoyCdziARy2tsoBIsg
InIAvmU57AVAstk8aeNyLz8WTmoDskTOdkvlsg+8xFpJ7Fe/h+6csum6Ew20ju791kEAK0xR2Ei4
BZzLhr5wh6hwp187tNCN/5PdheXyTp6b6GVGrWfwr/ICMeNzyvnzUhUMYbGvULm/Zn4PstK+ifWj
sVde6CrnvzHLDnO4UHAypPiZCIB1dj418pA0ZRxmvWESWvchZEM3DNmhlCb+sN8fmBP3d9wBifKl
b0HYXs9czGVdOsavWXiZZcv4Jn5IHkcofBMVWDpU00ADJ8uNfTDU6CIYHcMp46pNHxiveey/AcwW
Xr3BOUH3B6MYnhxV0Y/V4yn8r5zKtwuxb0vzp9VK85dZYp801CfXrW8mFNS17aRv7sGcHUWGZv2O
vwMLXMDuejNTUs6JMft1U5YR23tWBRlex9BLSXFsyXLXXXda7g+je+33s2ek85gyw30rg0i+gEE4
VlxjkvvFzT0/IyrazqOGH81hcMsps6mgiuBJjwauOZF49FhXrsWL3e+BS28w/JaCjXpCHFaswxDU
+zDMvn8r+M6DXxhH/jdz9F9iMJqazjxZ3Pde+lu7D6PLGcqnFKlIllBrjKnZz634KzH6nVkXNEuU
yfIFk46iplDTYveydvB4kPHQTqxpcjyEeu/jIi9TQIcVDvIxfawglTpmqh2NmHSDPh8IYdifYt8N
m4bRXG93ury0JG8z35lKKS4DcUMBLX2rRCMWVR+3/Vkc3QddF8ds0iTiZhsMwizndMk6XA1zKFIO
DZjsBwSCcSirrvboiKWX/b+heKnKrZofvwAz+QQtcywQpWa+35rI4AmTbQBxYCVXzkGyk9Bnxai3
AYFQzKPfJTz6bwEocibBjC8/O/8W9KFHUlEHt6gJRnD+c8tEFQgMU+yDc22VsJiugYCK4n7NFCUD
oxh2j7x4Ze7mbLoqRYUCl/i0kfyotIfxzKleRbzHFtDPhROKqtXKP+EEfHHU1EzPfV9sKLgVqwgz
leQJbPtbRUtGUAcADuRCzWJQSj4ultoojaz8w4SVStfdRRaebtEww6IPqkDWRynbpZqrhSGOtwh/
UyM5n++RpjhtAFd/RwLj9K1tcqU483WdmqeRw6wOTNe2xGE0qk9mhAjdzPrjJBM6NKbYEf3LCmwO
K+axCPiAu9mjMfLXAfN+YuFnmBqLpLMPeIpnifcdpcdTEfkzwDIjXw4xKXG6oDU0FOySpYy220hO
A7cglxao3XG61J3gwZjyMGSBR7hut4SigM15BGzsrj5rXHqJitqQSBGmyxCInZpTuR031J6D1tJV
Oe8EOx/3seqIKSZTC7e9vmbWj1rv8365UNb2cGz5Bno+71Da2k/Z+Ronkl5U6/vr42zDDj/WtIo2
x/2XFlWoOJh2CfvPOIrtliyz3mroRsnrg/FlKgHfXjuah4zlNybY1gGfmdrebxxDrpAUrPxe5+5e
wSAWEavpAQcocQ1ygZxuzzjy9hIzqNG/GL2mTDEc8dVQzZeuGA3Yq+0FNQnEpDYLsQxKwdWFJ121
nGPeftVqqhwusI9F9Ib7sa8yxhS2YHQaqqICELOShAoxqgfJAs/vTF7howTroXT3BJK57Ot8ye1/
hFy2MUCB34qPK29c69EwXjUAVsdolEKX5Hd1Pr8TTeHWyCL6U/hC4ttls42aqfyMrxrHUYD5ps7t
44J7NDZzA9J6oaxJeqxFGuaCqkNjcW2Jx/+4IOH+E+uy6rZOgI7VGN21m2rSi70UzRtn5ZZvna2o
0NBGlCC1ltdKktBkvTGmcPswGGRz0iD2GKOqV1cVDPpCcdyJFnronSn2pnez8/RGmdCsl34ewiL7
sDj8XtFLU0xdPyadorsL2Uaw9SVKe9xl3oaWzRw49eVTyIohcop2hza2FjpJ1HbFH7xCXS8b6/rJ
FGOllqfNHlXkKB+YvW5Fv0ul6JO8CzeBJJC4rP1bf4xvMtIJRu2pzi23XoaDIy4hx+WJ11KPkMhb
zNFaG8BwpZRr8pemS0cLFeXkrkgbPaYSz9h0WUqsysZSNKllNB0ByHLTkzCr/iP07oFH0xOWGnQP
0B9BpvuaScCIGRX3R4H7mT0bTurMXIzdT9gpbvEublcZYNOGTlD+mDS2iGSNnqk7u8Eyc+fSiZiy
EACWYPGZ7fnIgzNS/98Lj09ZhSsXIxiwEA0pIoHU2UQ7VTs+l2tpzCXCUXYSS1arao6WpOFfObVE
a4B9q5YUu8nNYjvISD0U8+joI5oXylJhgxCd1zYyPA2P8/l3GxJ+jB6URU5Or8V+FJ6it/nONSQp
QVWH759cKy4NB4ob9/ANPc7IyhJ7BeyicterLJ3Ep8VqE2q+r/6uciPNaKAFDcDHuPa8F2yHO9YX
Mswhrk0N2+J+LtDdZ4knbuOUlqw3EIjW+M+XTtolvjKXnFf2UnR1bYleOgZY97SI+ZenohKpskUJ
fqjNsmhbHA8tWukvEQF/2nXMdVUUG+E4jDE1u2qafEimfu50oq1OwEXuctQT/h8vS2F7dpYaaf5i
2Lft56XDhCDXwBhs9GhJxxQaC7JIUNk4PLupiQl+zpqKOoLfRT3B89IDemr8yhvjj+MzkrrKaNgk
rWbdPGv52XodNsU7oYBXrROOSclZJmZ//8tPyCUaMRGq5C6IFnR9nIad2qcTuI6Et5D5rdxNXkF8
OjctaUpQ9k+dHgntIxh9/as8HBTFMWqFQ5SRCj4sTqDjBThyWhij1eyxW1FlooGESUAcZ52WSbfi
awZj9S9JUvvH1LbNPxBsc0pM5or5AILTrzGxj8ZW9BVAafUSf43qNTVuIiqTqK7WaqD4bWpFf7oW
3niT5okvjA/AuW5emoZo18rNBIrM26Wjcph+T3IIC9sKK1jevQjrBgG/8DyL8A29mPqIHblZptxZ
tT4Teb7RkcSnTS13CBqKwrWrB98/8TXU1YxsgvvoqtN6m9UdEr90g6kbflr+nS4aB8SD0tUHbJve
a/EYsC1Ri9AhFN9UH/y6KoRuQz/zQ88GW+bU9ZI9XKXF4SsLGHj84embq3/IVSXanz+zIyud78+5
QqzzzeciPHZOvuG5cCFUgpBz9CqIaHhadMW8kgrmF4zdBV/NfRAYi8HWrgwZuZfag+7rI3yOVVeu
rIW3bOJH1GMW5nbk3mKyqaJwDmEZQ2xpBtnQkCpLVw+3Zra6HGxau2GfBAu2Gy6QbRNapIi02OqJ
oigZ0JzqyUJogUJK8DotBM+0myoHc6BbXas+OaGWcTVWI8fhhf6Rbn/2da5/LxhVLBOEQEX7ji48
R22q8Rycks/3IU3Ux9ipbwxFrkLccHPr0EUCW5ooX498dNBYmOzQBIFTDg+i8tfOVKbDkhIAyKw8
GS56/O+Hol2uOeBQryhU1FHoCAr+s5kvpDJNWDKm69rLQjr+J/QGZieoPLdkITjFIuLtLIXggAmA
+svZJgQck1EOgQm1oHV1KDTw4E4Sx6PWZdy3GOI66tML9G+we5moq4X8BMoUIrXvISxrkE4/fSqV
vdGlVy3QrLHYQr/80CAFiGYaKodaWPmgCozUJB4regJyiJwj7w2AjVUfkuZlMkjV+MFpAm1zv5ML
7juge6VkC+TrIJ5IpZDq1cXeVyUYFncVC29wSfK3n1YQXLNA1f1P/lqGhw4g4R4NRT8c4rPSahXA
dwN5auUdwaExGbKoOdx8lua3DapqMi5sNzsAyNG9V06Jyu3Oq7KHyhVzT74jaDQcCWJvniSzFk2K
C9Bov50i63A7ZcRcmt1mmBirnc9kL1YV2nHUN4clXtnG3RJsakPS81WHG/mJY+8opWOC7Z/iP+mh
cJ/2dAUnVedy+E7DgWrgHSAdWmkt08SWunzuwKsAeaC6B7Dhfh88ZWFPVuCZBmzr6IRfRWYdH6fG
cJNocBQbyoJIGuoNlddE0X4LPqu8HMDCU1neIsp+oQDf5A89loRLsZ9scHeujHfmrdF9fZ72N//O
/Tn0TuqN8zeIpphwdIOltHuVchLNaQzI9VQtez/UlyWZEZFGaVbS41ITqSpfOCjc8+roICogtzMT
NEJEPUMKg3wYLuJewJhSoA7uNIJ8UWUi7XG/vKSqU0lCDxqwwYHdr8+XDq423ilOQENqpJwwOJNT
9fXiMC+IdOUU/Nw1iGX1InKOil73QEqP17wpMawVKYFN5IHJMpEUvsdKWIVWgp9pmxnUGxyNFtG+
KyUoq9g5LkqupgqeoYYHbw9XAsefgeTbo4lb6WdVPRHoOJGkH1jh0dSk5MevLFERmX4i0XvRCAaZ
cobDr7vIWkZ0YiKVwMJmoe0vGRa1vapxyBTLc+zlpOwxENhiSKj5xSuPbayWYjpQ83F2aksRatAr
YC0nfopLrT9eM3gOXycACJlIPCLh7LYS+rE48YWk3NNVriYcABnrn5oXXGGKJCWlC3lhUJ9KJbDJ
0Y74sOfgthxFdXatGdKJ6k3qTt7NFwr4oAq8h5pVic32yzmPlXXWr7904x7uR2yomKycLoM2Lbvj
jgPuf5T+0Jsp7QRsDauqCHYAHBJJq1OVLsM+7Fwcbs5BrUoAErfA3blbA0FdYpVW4tdluNlfXS92
/snjO38XleMLboPDFYgPsJC+GmHFqWywBvjKiRIBDi+Ua2UtGscWpyrgkFEkywj2BWcdaBM3p7XP
vfBKky03ggNZUrRHhCp0fMuIkUxGfyLlK9Jd8UgK+3hzgAPdtNfgHLmlpI9pgjbRPM0OIx9+fnzg
HZvt1hFvt/rC9D0s2yQUqygG8e4OUpP5znLXYzsLZbh5xP5ZH6jmMcPj6VYg4bSolpJxKlsCQgE/
q3qbtwxlJD+p4xSfmBNmRMY3v3QP8MO2Hub/Y5W5QK8g3Lks+fRs7OYbcAwlWJy+VVQ14kxHOoDX
HNc5+KRNPf8q4Tcj0wacKMyql8QjmhfO8r0Ogjl3MvSKP6m5tbe9lZF4dzp6nkLLc6vcki1pdlWT
RoeUbFxm2uvUW4IeGu3tXJfzRSEadX9FS7F/GltnjtRn9Fep4IlCe/DOc8DSwbumzNa257RqK7hj
t7AXB9B2kDPm6w1IpYgf4YfiQYEWXds3aaDayf8Q6Plp4Fy/PTxybger6mN8qUORmww9SA1SJHwC
OK0gN6F9fPESQi31IeGFcmcfPWkJe6BWKim+2A4hAGspE9ZZBPWq3JPmqwX3vBRccTEvcCFFm735
jBM7kXK8R5nJYBkVH5tS98ks5pBzt+LohxkQS9ij6AiHhSJVPAiuLAD5ctNt0o4l/BZsI8mDMT1Z
P+7gKOI8lf+ZBTbQ48+p9f5KzhQ6LuM4LCbMYrJOiy02OSfhpUb63ZZ/FgvWJPqAm+5pWoHaacI8
5Ah+SmamLei6j1wdxXxQn1IerSny1T+08o7rQk5eq12ndqg5obusWVlw+/pGfXCAjhLqU6bwgNmD
b2CXUFKpnakj45T5n0Y+WVlRLotksXtzjmlGQu6aPwnr6T6Il2O6a+kmUAkxL2xOVr6Q89Rrg63K
plbNrIlPMe2iW0idbvRd/SmfhfqTZcMDAwihkn+ZCdp33IJgqipGv0z92FSz4QfCqrNVdWpIy5hd
4nquf3CVa4OvKXpKL+XTiTSvKc3Bcq/8hYV57aBgfKjgvD6wwYlahiI1IQBERmqc02mrO9OKeW9P
qX+ubEfySW7BZwMc9gfMYtCkg1lJakjqr0QxNrqroOeJHfk9ujeEFsqogKjY4Mxtk128xTugODEI
CG8fh39hQ0TGlMgacd1z17vf/hJGgQ0buVVzoY1tcxNkLtjoFatUBA9EoWgz7rQlO+K1CXVLRSvZ
aw9wgipbneYG0tKcCB+ZP66j8QPH4szVpKPfddbc13PxdlvS7puSOIMUZeIZgj+/weuKHtSdmzxU
BIhKUFtn3v2lTyqwKhG2D6ZeEkw6fC0rL8p38UajRf2cXJu5hF3ocnriN5AOyXcFd5CWg0KTKOn0
9O1uVUvYfKtXCfM0DCt1n/SIVtTDiBflwHadQ9yAHjJ0xwEgqxlJqtBrZ5FwlJJQ6W33KgkJ0BM/
1I5THla+g3CgVCcSll9cc3jfsYZK3heKyF2GDqHa/+/7LesnarkiT3QRv38B70cwhQ4LrfyQzOCC
UdzTZq3Ai6mQTG2Wbw4g2KGoQpOlHw9/h59OSvmrr9p/Iw0cDacALgdr7Anwjg+1V7sYhXrQGwf5
OBoV/voKuOSSuvrrQI3I/PXelBcakEz578GoSmExCfb9l3jukEzJj9Ui/xeQAhQkJkuKLO9A8YLU
iddG3IiRIHpuXeWyRxB1veRm+0cilUWipsp43NhVqKGBGDwfSRZqFxs8SNuqZusYq1aME+JLwJWQ
FXbQhZr36J076iPvfN8EpkJmEpJ/1rO4bqeY6alpzQuDb+iXY1zvkdQw+up9RO84+nOsOtzvm/jY
vNZcuHm5ZiODedT2xP0PySBYQspBEM0sf1Zq+9+Bpm2R/IS92Ku+op70lGzRNGumNAiHMX7HiICD
CCqrQUj0AMY27/+6mQC0dv7n+22WiXrzfV4pX/g9Bd9MXmmTaLP1KY9hUOqXtLIH2WAUDkvjziCz
a+g8p4KCbDh/SMyNMXoWLd4t+RYpaDGkZzIQdu1EpTUZ9zNhga6DGCni+uL1b/TUC/J75KUDdUrt
AENWX9sIC2HhHEbCkEU8ufyheHRpKdP63MiquuGzFatbG7kspPPgOOysArZIcVEd8ENYxEgU6R7x
NvcHcq3qSymdhldgmlFtjZEavVVHd8eBhHLbW6sEPty5tp07IAGk2sinqPZtulR34y6Mec6Pw5lC
I2Xa5OiUX5f2idr9fEijrs+Ygw8fEBSvUzWlOdJGq+QJHK2n9OeNXtouI1LBgNxitvgJpIWyGCOs
uAvVS0uAdTCMcRsbvGTRFRTWzThgReKvn16phFS/oNcVH7fv2ACkMkt5WE+HIp8b4QDcYvR9gDK9
WVD2+u4epJH7y8v4l+vlSTZ7N4Zas/Ydlt1dL16cu99zZBYEJdRhE4i1MoIo25cAvoaNwL9pgx2c
98DV00c1p5HLvWJBbZPErkuon7nFtN6LmLbLZXgzSDBznV2BshkKTC2o+/BVXFo14ei0Lsxu1qxv
+pXpshQKn9OpjGJKO7lJ/jas3J+DpgFJIMKt2b9xFrf2zWPj7tfvsQY4owRlpqqSKzFO6MbZT0MS
o9hqVWDI0R9tad6Deyp7yaav3hB4l6L3lZNNxVOhj/O2z4tIaQnfUMgoQQur9V6m1AnnY2dHZd6k
f7v5kr07f1X2IEtmKCl+ryq+W8Ph4IXN0cuiMIcgzDM7oINNWoBwvzH6qZzfjHejDtDvYx578xG1
3z9EBnoJv2LqVc0/VVxeGe9S18SOQnt2MBuG7L1G3s0C3ErIIUpyvX0wuo6MhUA5hkKyD3/rO+9c
XczxmrEv1heESludBPzVphGOkhnuRWOw4KzPGC2/d+SPs2HPTziyDpAqZtqZBPjQm+DWhQp5TKnH
3TU9j4HGMTRqhiVhYnnHtbs0W1/YGFxGtNCo+e9YTdY/3Mn3n3QJGiS+RInNEkZyGx/ZNCp0zjcb
52mawb48xMxGJxUtt1QKxqikC+hQyXoX1fJbjuUf8LgSCSkpmGjIxFWlK38AeJHtwCGjHu22CMV7
hKwzQJFEJu9yKrVP+TKR/EuyT98uDtxZFW0GCE4aIT6ZupWBsD5e7I2LjbokpgzbQI2my+O14SbZ
PhekLJoQP7DEZkhuFynrDhLEgCXRtx0d07ptlqK9jFjk06Ygw5igncciin3bb4yc/Bm9KM+MKUtH
qyMBmks00cm9aGXuvNgwq/1ikzwgjoyZpv+/6Pgec2PmNahrEJWf7HPsVocc9ct6RrwReQTsfGJw
Ge/7kBLd6zb8+exraraqrXZJQu6ZWMNFvZfR1lMoRdqjT1L21+PgMRREQ0jFrtNNPlnb20w7HGje
563t6MyTWoqpWm66j0PWJetbCBfTOJoJB43s772tk+F+/Cp6n+v4/P9KnS5XUZQWV9eNOI3MJCfO
FoI9w6l8v/8mkuGM3mho17HkleF7FDudl7z1Ovh6M+Mbn/QCkTmQ3eFHdcZh0lPJWGjwfWxuSRyI
ImZ29OFvZG5w2/jV+M65XpzWdwbUi83jqRBA40HsWACqce4Ocdlyl3MZv7a6Ne+WND7oCLm7QLKL
s8hr37807CsdH6lhEsLMy1gKMVDqpA3hR4ZLIHmXML2QoaKD0/S034uCZaWQgGBvuBgyLME3tY1c
262oI2NoS6oM11U/0F/KAG+5ihfq8pAhNGvEqw9PltXJlUBKMqoRzixNsjAQCTbZg1fDrcgo+Rs5
vXOPGUldkGZ/iYQlHnof7sZTxLKRhhgu1w/xPKzBgzK8X6vTAEhCiw5IG2dcnjCFUXfZI5TnZ4Tp
r23WKKfHS2AJA1jxBeYO3uxvXTlLXzypDAOekYXxD9861KgxVONLBjYWO3vUBFFkhiX/8GZ++PpB
iQ9XejaczbZM3a/dctABiRtsWNm98HzaDEXied02XQU4+LYmeuTl2KACAFqCV62E6v5J4WMlXb2M
fEVvFVKQEgfOUk1WwWqHh0E+eadayN51/VENezMrYxuo9vALmKiEARSn2nOxBmaYObD9KMa+y7I7
q+oGg2QxbJjcEZsgsd/9HAIDaC/wz8dYieMooIu7ZJmCJmwUz+mxNYEaAUlCRiJYmdD82B8eqDU6
D1sZ64ALxNVRVvFldX2x8wirRM24MYiDmDM0tU7QFfGnA9u4eQ/r+3cEE/v6C7hgRp7Qo/Ii6Cxy
8yobVOoBB6HiTMxE32amY+UVpaRWPpzTSwZY992J4+Msc9YqOV7nAGSX9eiusRPCTCgBjMAJjDbo
sMaSwxsCTe2aE4tJFFukgM1pPKD7srgBwX4A4Br5EDdjzdZMinlEWF8lyiORp0bI1AexhOuGcwUd
lYC99fY+5AiK+PsUhB2Ls4PY6eXF+vOaIEcF218MRuRiJjhqhqHYAVswV7i5IP/OCrssNSyPVTqF
nVGM0BUxdMDUwL4OY4iIxrN6Q1bVERWrzFax0GAV+GXCS7GxRKmoVbfqIC9apy1rs6rtgO6ncjyQ
aaq4dM51cdfXnUmtCSKELJuvaPXFhmJ277vJyJgzKnjjOMDF8pAqwlYYISd9AJnepE6KoDnRHVxn
NddsrsBvcLrUQnLTatsu4s57Ed49Qyls40GWZBqBqCPilzgc8O86U+mRfbp70hHZq65mZ9up3PFE
DQQt+iAtk3rjXv+xQrgz5zhJ5D9eFSUyyPfx02xmvN7LKvDFZxi/OD6qZYz1KBbAWjt8Pj4vLXsc
20XxQZ8cVHf2zFQCTQSuTGlY/+IyrK7dDmwBeuzAN6NpPCR46b2EqYplArVuID8RjB+EDTh+Xfgn
4Oyji9v9z0+cCmHjCGLtFL0P4UhBGIKKouK7es7ONx6DTixqDO1pkRsQoiNxWdz5PJ1LLgwmLWP+
oY4HFz7KSKGjwTsw01QdniWOCA82XplKVg5dZssN82gytpwr+duyTXDhVdPSeY8mcGAudtEEG8O3
u5CQMvjeR1E4AGQfwFls41jJo1T+2gypP9JeFWCqQ45TDXYUv7PQeHEzKnKeIYICejOhMCZJPk9B
aIgvOKm6LeLfZZu/Mkhho2k/LjXDWQ4hOVE9kl3tFRmp8bEjXsyOckAmjxwHQa2koBtXrJy/X4+t
dNB3wHwK45UXOSptTUvFHO84tMxjFObkkmJ1aVI5wjDnOmreLKAT72J8ZOBeVnJErwD2sr/gU6Du
hvrmi5q1b2T0N21Pygei7CE9MZLsYWixAS5SUUEINJt8Q5lPDH1gTcRBolAU6dxjtEszeMfPzwpl
xnIrQfC57pcoleWY3agh6OT8ZL2Keu198gpjzltcu+UbPx96JjfJw6+kZT0Gb0IKvIxPrfUynj9O
FcbRT484MezHY2Z+tpKLLCQeOfZlvhuYJF2N2E0BmZYBRptzspmmCeLeXS9eyayUqz9aFRc96g/y
bTIpWWFKYTs0CF+TP3UPSVOFwItTHsJ0p5CuVMho8YVmmCUu69C4NH4UgdTB/LgaZJJM0pfnokCl
lUiNlwpJsEtYcQr57EX9VFOu7qgTMRqhTUVHDXW34eXLjD7H0i1SdGAZuayKHsCksJ9cj0VFH/ue
rQ5v7D+zqkXQRHW9O5ix6nEl/7YIPIkuLu1CjPM1ECgE+9KHmoGRgM/PHC9XRwcfKvDYlFOoMewo
IXgWV52UJCIjM0r0X6k22BOpECDTPdNUvsM4AjOtRftQlR8i4OiUNiMMMNuE1HAnZP/dCheubIs7
v4sUx4cgSgPlGoTCBivPbXjogcA+Lh7nq4JDaUunjfIZDbCmucsr3KWXoax6M6a30d8I0gCConlI
gZnYLeT1e7Q2W8bqtRympjPH0PAY/Phl2lLbDonydyhz+WQ98LkZBLSvoWGGEI5dLQoTLD2BTUTr
4Ejz1eAquYzgzsJxDzTekYivM5+7+nCBcrPfb3fffsXm6NAKiJP9BrsiDUqgYPb37NJYIkBwv7JK
fTu/TiVEf+Qw1pga3fLrVwKrwKPo7vWRehm3S2tgQUMaJgeTG6hK6QxWdCmS0HksKW/yFPVmF0P6
lxNmla24TWVeakZAQPXMADFCc5evFqSAKgs43jyni2LmHcAbfGP9eFdswtO59S8n9LIpcpVwmyJF
ddZCEJX8abr3edElHrAX6m+jRZixDHVfvg6xNjJLOtpxhJt3zWKezx1A2qH7OCSzg/V6NqiWmv7P
EQfGBsqxjAYQxjvyUdc+O2/wq4RFv81u+vPK0S3t/8kICQMgCFlfWnd+U79j71fI3sEAGJ2CPv88
c47q/uFsk78kVIe6B7dq6szvIArqBsSmuscf/WJ99wErUo1G5aIUTQwQPDVspMo51CwQ80g1t/RW
6JNffefpDTz1opKbTdh2O87+l5cso5e8W3OWtobvoREJyZvgRwVBMYUnvtdUAdpKGlansKDP4g/A
ETh84xOT27CS6ycOMOqy28n4KLtsk6kO97wIL5w5wyjlsBlj3oKiQszgN2M5vAt3Zfac9AYfxvk4
d9wSW7V8icC/64/kOn7V/DeFDBPWzHZy18Fqg2gwQnblB9seXKQC1r1zwU8TpXZrv0WspME3zgQk
aJ8LLcubtk32UlirPEy7NEECDFZ/5fKKHqJs56eioKH2uvV0z9yhJiwnvljVM/7ZnbqjV/d5DvUI
rXYnwk2UTO8uzG+PyYRLTO0/1ezgKverBGykgBJzG3sHeX1vWlhyRzsgpHIhCyL98u9GBE//bV+F
ruo2eloSDNByUmk8N+iviZZFk7wR/biMpa2k0udtGjdQYMqRbZrsBmqylaTwphrhgZoHkfoBwosd
PfbRuYr+QMjvSB8bWbWnZC7YYmkYQJmZU8giV3MV8mX4n0RKqD/go4c/OrpDRh0Dt0ByR8MSrTIX
PzdyPzta2E8rYDcB66wdmxLI83OT4i4SgLMQjGP3Fi2q6FA4JYejet9CxZw4snW7STuS2dtdJjfp
M0/MXlIqvRgzNgVB1uql60/uxJmiT3dlZAqH6tpsQ/BvhLcf92sXtAy3DpgXgxxTK9dt3OS4vZ1/
aA1M4vUkoStULwAupAsmQhxeO0Nlga5XDer2LPx6FBxOu0O09HDt9X4FXdw2RvPQE1/FLqyer3Km
RMTViHZ1Bnl34mRN6ZSuMaP14Ynu/7H73PYXVcMzr8rukxr/75euU0ZPFymgWQ91ngWFpKJtw1c7
CqrbLcP681/Bl5SBImepj3IeoPNu+8QRX2Fpr4EZQ3HvAoijrdpodYe1xkivZqWR3IYeWGNmaNcr
gAWguXNf9EXEJB1wvfosoFCZFK3Q1GuodGcCfQz8DKygc5Cle5fPno0gIroWBSMz4be2xuDh33W9
3MbPCyey3Fh5zFojkTgm5Ozk4YEQ1E1VyR7rDLf/aFtp0y978bpRZ3uWT1uFm2OSo83EFZTNtq+k
9O9jHlojB6dLNJizdu6en3xvr+sHuM5OYgSCNQ7s7sf/f3Rw2KQorodDer/8LcoOTmVwLinwoZEN
kMvfmhTSPVFVNTs3Z5SX59XfV4YSuLubLbZPc444L++sJsJXJ8De1UM6k0LStfiup5O9a95xjfou
dDLHkW2Ae9sGNoeTJRn/EIyhPkzONFMGCqixNBee4pHIZkAnzHPKL3voUpYwH8qR0xUnQdYzKbpM
L7f/PNWl0jLI9/A2TilNSKmclTwtSsjejTVM/M8CkEOBGiChPV0+o9fMwywfl5zkNhGYUGe9mJAU
Iav0vPcMwqHrnoxVhdrp2F25MBH7iHdIHwyygcBcLU+lsd+wKk5G2PuwZNMD7YA1BRIB3E6Ee/ky
/Uc301sqsK+eH+V+jXhEc/J9mckZVv3pdBElUROuTNTsEr01ZKhLfA+pez+QuxvsroZj1vHzT+ym
r0duuGECTFFdo6YlYSgzpzE/XDCgAm3S0NZnWrZHWude7jeiUM0kfnMDB8wIiay936FsUGYxQPcB
HfW1YnrG0pYv2UB9pgsBxoBEoud0euN9+WtMIeqk0mmir3aO+yvSbi4iAQr4bVZUBSt8Tqgz9CmE
GhcWQb/jP0SF70afYMguSWqeIHd8gY1NpddUB42uhVKMRQOW9ZpRP/AvD0VCK8oLKIB4dxIr/T7A
reXkWo26ZjrD6yb99H/YrOP7rQdEbch/cAprdlj29fnAcE2MMKON6bx4NC3kN3STO88be36qLRwN
EZPur7w4eQUxo2TxktmypSh1KCGgCZXeYHUSVUCgkVELDPkhZVxelNgDvM5zvFaq8xcyluHmv1Ds
OmFT6CVfhlopmWx9JEcLr1JgTVhbmWOzwLzVqP3yeDNRhvSj3gBhEVzGG0rI6VHtJPVk09moSIIe
R8hzZxlAEWdme3D1jnSG6Et4Z9/05EE8EFvKltTphABaTI8CbJskaLTOsPaV5u09co1yCLBjUDl+
fR6JGa6NzV3DYK3+x8ZIl4NrBXWLtdCR5YjrKJ4cDc+aZuc8yAvI6x2CFxxUq/TIF7k1ltO3EMVZ
2gaYpDKLiT9PAZ9hBIV6GkdoUyLE9iI7CbasqLdygvWu1cf2+BdroKM2zOh1qgN4OzsdrmwA+RUO
KAYN9useu4nDeoXedlWMT98B5j2DIqTcZ+nMo8hoxpnruiDFuhl2i1MvTF8qHl29rSQJ9SrC7Sw2
oZ+Y4HwlOHVAC6T4J+DGKqGF6keqdNf3PVsjYW8RXBCMOpF0BVbPUtX7rS26zEbaWakoBAm4WBm+
vTD1VJnh/zHLS5ZMsRMX7F6qBWoASh/RzYJ8fTeoaFaXtL24jzafbAgYBJCCaZc/cZcGq4GqtrPt
DTpxCAkdP4IuxEWdX/QaTF/4xSxSh7X3hkkU0O7purkxEFEnkfiYICU+ikwCDgbBGHjbR6aXIebk
PLT6V8jQ62j6fPJ2YJE0cQd+SlQMFcIBHg6kbx0eMBNRKV7kwcvqrdpg1EkcsautFPIPc++Wlx/k
dad/rcG61nkpibdIQTJov0kyYuHWpVZbsLKar/DnUJOweAcL5/Dkf0Dymlid1kAVrglOnBuehUoD
m4wwwlfrJP/wBkBBebrnZrJx2In4prJHtUpvv8MZWzCRO3KUJt9FIc0gOb1QPy6RnDCdD72CJHC1
IcwhX++kVNCglzFutb/hMD/PFLj6WSbTU2houEBL58ND2hvrnW9SNaHadWofLXTQJ5W9ajSArXG8
1ko17c86O5NTmLpFfoeGAa6cIS2bF4YpcxQQObB4JnamIfLpS3OjqL+5D1IZNxnu/hpj3OEitiO/
YfQd7B3ODGQCE5xaN3Pdg/mXDkB6OZylnhZGiXdgHcK5Q2sUORZcV3EFEsnsbseBbGnQv33B7sX/
XlwBJytN8LXhJtU9ZrQTQUGVb+tXqXenMDmA3Y/kV7yCqzZrfURI1jEgHi2QE5l+RmWCT8t3ZsgU
mWxWEUDwF6poVCJDi+DWq7IybaAr8LgpqnY8TLaMQ7MbK7F49JJk48MRC8dM8ZZhUbaDhkYzHo62
NqVru/x/AQp4Coc9+lxX3u0dMFUpjJEma5MGpVL+0ALon5Eypy8z8G7dSi4UgccH1RCdHCZ3rYBG
Eh9N9Co+Ea3qTSEkTwraxGo+VrrjLSM9jnA3JroChPrl5qLFfyVqnTBbmcpQSAjp1sGpZ6Wf5z1r
sHHYYCAXA9wJTp4HTaY8LM2jRLdxj4qP6P9BcMkmOhsi1BQhTb24PFlQwS2bevhnY441JLJf2AAX
tVGN7lHXrR7V9QeMCAWaae/RSEgPxoz49ymRtNoX4m6PDftSHbgjuufUtxvii1RKepm4Q9/FMywA
wgoMWtFhrANMyPWkUR065hqcVDD32imAFy5KaLFTm+aAz2UEv6YmEyb5OLM4OohsQi0q8z1H1VhC
WiwhPqr0xX0gE00RIZLJys9p5vot1eGzCQvALx2g1xZSoXQF8ElM3cYPfXX65NAiiLajZz4C5GUV
5LITUgJ62FHB77WAqTwLI4hMbrrq+F2acJfC3HtRg5SOxXJwllSdxc1LyuBxxSc9J9ud0YSgJBI2
4YmaJkckYb9YsUMZHFUGByCrMYa5KN1qqqB7c8kcc67L9eqLYGSjHPkH8suNPFDcgFJ0dtrQophH
XdNkO3Q/WlCrI0xrtiM3Ko0z6stdBgvMmbupaOlhRrHv1R9AH8Cn1t6EnWA3R/buyzYIMJsBVCsE
q1ebNOn+lmvF5x5KkLJYjv85XdFU7ea/Ef0TvAWXaOndg3JkHrEOSwVlYCeFoBpcsy3wNTw1WGV4
h/f2ciNCjRxM+i/O1o3Dnt3FgIH+VHKYwL0RO2qBuoIJv92/Sqihz8NPA/YY2BdygfBFrnTzSzR2
0m39++f5sRh25U7E5W4jCM95ZGNUpkZVPx1hbr1zVwCgmUlxhoXeweNIvf+pehZDw3YdXvJ10k4y
H8W9up1M2guuagwVslMiYXIBSn5/IVLe4PRL1+6W8GOfEkSNkxGUYzsQCsy4w9vxBUH/3X8oW+Po
C0k8jcirs6QI39dHqvr6AQ6w2FLz+qbi5oZ0+SmEqz7y5+uLupY9Rz71tvye1Z0Ghjfv1YkddHt5
cRyzeYN2SoJKQVtzlsRER6IuDCIXSr7q0kMMDwBDQ9JhQGy2I+kCl2/la2bgzoL3/4LBoNeVM5kg
3hScZEHxKUgHrQDdzYb0/Jq0I1GY4XroUCKCNNOegXknOSkjX6AMJMcz3LXF87LD4LMsbbLLIQYS
W8gqM5/htznhD2Pj2dgqMCjnS5CyQ98Qtr4KwEn60R7FatyxJotoe71kpw3pCvI5x5qAgzAXMRge
5AYOO5NV1npcSFKuMJj+PnBwmT29TNxdasJaC9gaDYDCghKkPtRNyWYjH94J3Z9sozVZC5+E4jus
nspfq8fvwEoc3jUddKCSEBHKk199Dir3V4zx4bvXslU6E4Q14Q8gpmosYeI++iYJ9JjlOzc2qJSF
NhgYUf0XW10fAPdSiDnZQRO7a1RybwRH7QtvGlk5MglTVUiz/wCg3Lxq5qY0GUhpvV2EkOYHZBuX
Cqm6ae1EK4nz/oC7Y5WxvSffld6v8SUhTQFHQF8+KP5SzDbgexr8g0fbVlxxBn8Yl3lUNvw5JaVL
hEzLxVmCnpTvlvujAr96VL44JEqGTqK7tr0CgMTyJFErSQWnCYOfztJfaOtHP+NhMcJTHatf3+7B
wk6emhibN8A/yuJTjibhOx8BApYGgzYrJSQ3PlfnTRpJV88e4IMyMq6RYJcpduaoRFpsMpPXISot
rwn9w0IndZqF/MJq9DSPoM8ePWTFl+pQULz2ZrKNLwD08+VyxGUqaWOc/kEswzAwrZROkVCHll7i
yh3bVMjBVUPlxco0/VwKBqBXgpKyEs5kHBltxZlSP0H205F+RbhMU+K5M0nZz+G8mVbFi3976f3N
Vrs5bcFdLpQuaxv7Nm9nqPbuxMTdysGYp1MQEe9HKPyk1TS8TShaD8n3pnH3DQFd/demuMDr3jzh
puNPiKEg4saM30yOgW1Ts0SVBwt6drwVdYNRk5cGfvlLRKkvLVtFtijNQ1yJHNrEdshvpBiZ9afW
35PYldWwB7zq/6ZkKRGic653GumuFv0YUYM/p2CQZsAdHAZNwyBGXwvOT8Q1gB/H/DZsOq9ZI2zb
NZogufGH0KLqk2P7mdZ4TKJyRB14TPM69+B2aX0fsEmvu1t8DmG6tOKQYtg8B4n1HMS9g7l72gUP
Dxay26GUq/meawQzmV3tLwBrMTHJuK/V6wIwrftGp3HY8xS2W0lN/PC/v9mXaiWOh83FK2PCgqy2
jJET8cXuX1K+L5/jTQaoSjIN51kIYRDsPHzJwRnxJ3U5H1Gieb+X05W+olsWGhIQc2G5VxXM6y8Y
J6RmqAk4xZIkfnMQYUYVXZzThLRXoy/U3hA810ioNSMKckpu3WQaDTQR+WjSVii3dJRjN9gbKcBu
DGS59701dY+IuElZk3ZVrPO29/u89P5zEVgfc+XJUijfRSpjK8kCgA4GK1AMqYD9vdLzQcZgTlh7
0MEggjg4FEmhml7sw5jr9YfHvgxUFu85W93APAjGx8eG1tF+g56Vm1223gWJT9otaOCqVpW0XtFv
BFwTLgqiuxx0h3W6rAwemPIT1bGZW8O6d+jQwjLSGNKRQFN28P/sP28NKd/oV4/GTzkboOXd2I17
QMTeoFiBTQAl7AOOspqlDZCpWdOVjorG3142R1bnsnIHM91PsUkOoPsaYt3Hp4kjmbFmXc3Y2Il1
6rP09O03gyOhkwAd7LDwuLar+7ljged4Ta0dsLJHtbhKs9T7iDdXsXygSn05sT2avFayecXYKMjZ
ELtEHy8ka1m9DjCJYvdwRm0qS9avxyK/e06t0pGDhWwdKnpgtzzcSGoyhzXHi9trACHFtTGe+SuZ
WtntJdXLVmr/PI10reISbLxBLvjQh4Mf/yaz2K5c/VeELo+q//3JK48/wdcFkZlZcx3MBQVLpV8M
oL+p5m1wPWbdSe3UmgtEqKF6UCk/ziWs+kWqaUyyxi8mT3OX8H5c/60wQNBOikg1lWw/qTkdfA6E
FZK72mUaktE9zt3nzito2eetxLBSZSQ3q8daOGc0iibONjzNJdYk+cmFBya1na2N6oh0BwzcB6qW
hIHzlBhFw7CAjH3z1zeJ0wBR8Q1MZDuYNOTUVdkUxuINkMlZ8WBVqagHwaX4QFLMB9NPP9zeyZkE
5t2yYvCT+PP4WTv179hw+sD8o6ruZx5tWzItLqM78kUn6nsQGrG5BJ3dUgcH9rCX4sekqrox3ojQ
bIW10+buFbB295Rq1XwRe3ThuboWek50H8NurAIyE9rjGEaVNCFQqWQ3Vg2SD/Q9D4/9X+mVMUst
D4qvjAYJsWYoZoMwav23Z/6/aMIgPpTDFcOQUokyLzcKQ9asnqbBhsZcQbY1Ivg/Un4id1DfDLEy
WEPxSDDuglv+N+wOopdhs9Eqv0NNGpT8/oOhEdRr/7mV3KQquV3cNmZVbxat3feBXuy7e770y1ts
flb9PYGzlsFaKS5fDi47QKeqmTBcruS5X1utsIadwEOkoYA+bEVtupFrd7A0YPUGQQ4Bf5X+15Y0
B/mOQPB6e8lE1KNQwQ4lAU0R19rq+cTDSxKWNuse4VLAmR585goWqxzlrUa1KHxJ1YkS5OKrR6j7
EQHT3AYTgLTF04u+E9yvwGvBGI3vLOe+BkLNisa6+YbSmyKvuckLeSmLfIQv6AJxzaht1qhq+GNZ
XtmT7SKWjxwcHYdHR4AbUxBaLrsdqEXeh4pEzvDI4LMYCRtBn9ste1Ra5zPp0pNtpXr0WM7T1nT+
r6WiTHnWozwz59dH+2zTFwSWfuY+M3qAVwOFzWHB0v0zBUNYQcvztJ7s5XVlXnCz/hwB/RWUQrkY
WTVEah0ZxGb8pmeBhuumD54wCBsD4+70PMGs3UPWGQXYMMsEvhQjNpebe/ZnZDDIs6E69aArQSO5
x/L7F3IH92QuegWuKRhjjqeougHfW9MhGUMEC88KnF2qL331wMuYsBlxL4zMhc8uYYy0dniZmb33
NWycq8FSHP6GqisdxJ1CItIKgmj1jiV/TbVYnriDz3j8caoZdveKTiprB8B5U8rp2HGmcwfQLIl8
J2+BzEvqLc4B2AM3cK+g83odzqgj9d6M5AIRT/DfwuRfQr+CfG3FReVj7ykPGif3O5gr8Nfo/Jw+
8SgYh9PPOLKOCNDgjAKUV2GXlYCL15Nt7mf9cD0VR4OeA7q6KK3QTRaegHeWWq10v691Fd36X07/
IzYRBEXIRQuQyqJUfsXQ/vwFI3yy13STX0vGtiOU9zNsghChP0fekZjoU6QLeHl6iGgAV4YHwkS4
N/E1v3IJxdX7IHkmyo8/7kXylDzD8LRH9scfEbZIxgXXz+rxs/DiY8h+jnm05foVM5YH4trAe67g
cHzggfL9FdPE8x5UxgP+1mC4+g/wUxNgQjECzPu5sOCiATF2LLU0CMweciZqvETdgQhAj/g0BIoL
lyKbIeM6VuBF6vVXbwVVyjc1bhGC8iL2mmgxB9yHbxfnoHKa3dhmZ0QsrpTu8YDOoUgvfIclGIXY
MJNFPNJGGsYsD3P8uCVrsISK0i/CoZkV7w+2wo4PftzmB8CjDK4iIPeLhQMNxU63zCQY7VQDBctb
JNdFl4I8hBg5DQnlkifEmJxkxc5nKXsHhnQgTCvvN8vf4b74E9tl+uk2uQREAFFcbrYuZJPlVv0F
hT9YkkdAA/zRMnzz/nDMFBoklFBqfaioQCripAxcwv1u0hN7RWTw8A27wYhzFPxlMWfgyX12P3lG
pJMzW652q+MPn/KtJMeAZ8F2hu8CkiW1jVERI01w6JsJNaX3nq3DluVgK8xHTtm6722iOaTdWrFO
90VxjvyxBN3UMoLqM+oTkUsSr5PU+ph+7CTMmvKiQ2a4zQvTiSK6Gew4am4N4fXrWGtqFo68J4OX
ZT00yd+TFto/evyoQkYBtP9Ecp/V/oKCOF9cmN6GEU3qah05V+uUo6h2ZctT1EYpINHLhPxlFe8w
2gllSCMh+2egXgNZ12Muv34ZiliVbh87kqJ6VVpoa7r4jRDY8UGe3ujNa4sWnqBlJxnZDpvoyVfO
46Xe7vn8f2tdwa4h8s0u+zyI2lfmzFxZ2LZWztjFodNrHN1Ck804d8Hi3n1t9H4t0s4wgOoa+lX/
OPOh2iWP6WZpX8WLbeuVgBSL5TpDG+YdQFcIz/k9PvxltxYuh36JxYhCorMt6IZEpKrF2bawR+WH
B/WiXdYgrWSjyZpkV902EMPms75rJF+P9LJASo8avqhYX1PQ6u3bCrU+i0l6HeF8UZOowV0Zekcm
WC9P+eJYCjVvYuFW/pAia6S3qobGEP7FrsGdq4VYlKjkzaVJn/BG9MryqZYNU4y8pphoEdYIeRks
q/DAGWR9bF8HAuHsOySxQ/IZeuCQwHh9BPU1Neln9OMmHXm4TuDnPMhiGsALzHFZsZDAZe/aMnxC
V/YJMFz0lYEUNe2zZnlbX7XOuqN5cjVpwnLFAxlU2VzEHy7Hz0SIb949BC3nHHL6/Sb/WtLkGEcP
XCbW2L7pw7JNwxyFqzetOaiayALVX/nqvLbYfn8dE/59yO/EDYIey94Ae2l1nG532PjCWjRN/Z39
EmHJbxpZe744uNA4jVvFKbVgK61OJrRjUVA5M5xclgyom/dkRXi4TA/kJSJfcUXI30P2SK4lr3r8
TkbB+XgC3FafE2TQ0pmntDQ0kB+BaeJhy+CNR0yPeL5uXs7JlVJsNqlOTswyk56NPkq4r80ptmXa
DHu6uoCNSMy+IzxUiJkst61inVvuZJcbv1JrzxmYHlaeeZFtPIT9JMvBxa+XwlP9uLs2raB+BRJ3
ygjpN/s20JYpYjeqVHbJ55MpJO9AjtvZU1kvZXqKjmk/LMBE0ZFCrumlldn43Yf1XTkDDmm6KPx0
GxlQDTOtS8JV8gl1QdIuJg+ClHNp2dz1UpYXwOiCFjkBQbXzwraEEIqpf2lze5e+Ekz34Trp4CON
vwTQZ2g6/fUEzSvPUU3DOpFrxke5lpHVIkdrd/rTdA7oiqUUCVbMHoRMoWruxqHAZheRMktdrAHm
BC5GLgjcPH7dlAITSJZ/yg0AnP90i6EJz89b+Whe9Bt1QJxRHIsL6a/pTMSoFtvKBLjWH5xbLY8Z
QUcYdDp4DzAujNaCJAwZtsQ8gayukU/sLLJSKiwyrtYfGbtG37MG+Q31qtwHH+58MSSHIVQjmCbr
7jP5lpxOl1bxpOM8q5hZndw2gPuwqRByfO62BnqF7xowUucs4QL80RzLxHYba9xwyt+sg8NroIJa
4aiPoknPRsPfgcTlXdjxM60rSa3VtGejBT3MP8cJfj2X0n5W8UjiZcx0Zwh+bojihKSNhyyWgtNy
Zf+KuXgvy/u5ZV7VJLSwslhN2ThUfCGZOdLSvvFbhSrFM0A9jMzg3mgF83mQ/vSOEZaizm2YEkCi
YJx9EbDz02TBbBk9FDLFV01BWjppaloujifi981XRnJoXDZLnO0KUjtST+KwrAd7AuR+w5fwexf3
skJYJmpZlvHDQjHMhd2PPkU2EntpfaBhSxrLxfxu/DYd5H861/Y0XNnhYdkNLdtJiGJhysHRqjr4
HlpxXsVY2ePhwfq/5a8VfvhdMbehgHWxxdTy3d/2+K7TnzpBSV9HW4x7Ba98Mj2toOFvMEkUpxpd
OFHYQDlcvtZohlLWM1rWD/CgGH6wUuZnHPq3KzWF8e5G4CV2T2OCZK97PpzAhbYRE71YOcwkPLV4
WDWBnU//bmTjiAEqHVvKC3j9FgE2ScJOIAVChe6XWXVzpuLfPXgjN8lGuDCBeGZGF4PB1TOGvsjj
FjTHJniLd2xxcqfHpSWKpQW3psMQixDwDWmV4uiNn4TyvZyFTIDSbsKfcJtL9OpIaN0c8s98uHqn
5hH1LtlY5nLoehiOOiQyMCFLR2texV6qj1A3oupM+vrtwBHZcB994yYcZTl8KywU8YsJow0IZgs0
7ERvrAOO+DxEUGkU4Fu70ufILwitjfZLe3NzF65gw7wEVXmmWZNOkQDQk9YqcbMaDTgJSpfiQcQ/
7g8eeRoriLKu7m87zD0SBlelI5NURTL39QLqB7XwpAPZtlsza0hKTbOtbmqRCHXHGCWPXd8B3rdK
2edhu47vqEPFjGLci13klqg04hvjLKX3noSjt3VAqCQgYTiHShuTr3RHrZJgI/wm4A+NhR0eM5Y+
mobaDPikiD5xBMlhV5aOoESqoU3dHqNg2BAMm5puD00zsr1e0pnpaXiVdxjlr2TokU31LonNV3zD
sODddgg30ey2KtppSXpf5icBBOWOVC91z7YIPR7yqguh8ByEO+fvlgGiYsgT0tFbks3A+K9SZorT
AwXNftR2VVzvYloXGdecmu+nngDkCtbr9047F3zNGxOApesHbHDY1w35USzcWDUOh7NMnFEc3CLx
WZWHmO+j86XvVwXozWzWyua5RyTbVp0wAe6UVXaG1il6m6sJ6QGMhcLMHhVjWhwmVSd7sLRyIP4W
MvedScf065PpApaSD4LdjbhPOa3RE97DhtNPoKR45sKRn6/dxaTxFOjoTDttbD8bawwhZ+ICir7p
CfyoO/BGBnq1ed/qJbhl3flaFkvTboYVeFx5MXHw03FY34LfFEM/5S7JgHklNE+AG1MA1VPjJUEj
0TeBsOR/bAchB6XJN6/pb0mnJ18MSdWm7aVaA+smkyGLojDyMJIc7oF27+UFeYWRXtgX4njDii+9
Yh3GjulEWF6YvCCqKcQUgSm8o3hq4Se/SSFa2ILiM7sRqkLMzUfWLq37OJZNkfGkGRvJlUw6t4WW
tCC5/jWSu6C4fXqFjDmMgOGkf4kOge15QRWvAbWFGPJpx2schMR/NXm/dUxzOMTZRDIOt1TlOIRY
+Tf9/afCh5CnCNo2kOVJ+J4LYZNA45Ze7HFT8hELrqYmIFBZXJ1E8OFq0qHgO4zaPgqbewkwDw8P
JVrqq9qdcO41qql+Ws78q3+/AWq1sT0OVbljDJYKRsOg3LqhpC+ZzyNtVX51jv8OC6ndNxmDLzlx
Mj5Ft4ljr1QMvOmbPBOZtkvfRxYJbf8RnvoZRTuihybA3ZNsHCU/IsjCOpnunLAknaDSsJHsnpid
+khnGPdW997hBTy4EwQbtmnnTpVGLc3KEkQHuI2f8MiaKismJUzs/4huwR7Ii1BdKgqIZod9i8sO
g0jA0AC0OW56oTQmzJMaGztMCy1+Ew8Q/CGf1wIvOSVmZ4Tjg9zgILHXSjZv29DZFK1L70dvJemU
i7hs74c/paPoLOwRJAedDdrgUqJIMOOuB2S7wItvnRUkfR/nnoqeIy34SOLN8h1duGP1mFJhbU0+
QOJaddd1QfuU2f78T+vaX5yZXtQPw9xP6odemCqk51zmEqcXUNoum0huM0AteCyVFycZaFMMkZny
LnsGZIeZ8tV/7cxzE6TSxncZXX3UixahEN7gSwkPW/izYeOv8xziqQiJRbq6kYRuQA+QvEWO9ncj
iRuPAG3GRY3I9pD8RYR1al7jyrb5ElbeqjLQcG9BCClaMWTjssvH28XHwTmwUInije+xoVswuQxL
7raPOJpY4M7kZXln8LBIolH7B8ja3GSQxbD2Q177WWsehvpNLe4ERtZTOiRWSEZyBqr/tsfouFK4
13bVhkF2y6Pswc7rHiVd7gyJs6CksuqIsC4zI/+8ATMdLW+2pkjOs0FmhdHrRUvfsDZ0svdLifTC
swMlCSva1pWoSvb4335QqTsPDkV2KphLhJgg5T8U1yFO1ZwCEhq29S7XX7+smoXqb9clEfNiVRzX
tN8E6wfII4s0evl4PytqJ6/Twe231+w/ANzs4cV00YeAWxh/roLr4iEQKMmK5yo1Q1sNQP6g1hJ1
SqOFqol6QouXm2UfwsX9wlLofCIG4l3hDA3Cw7lrJAOnqKmdMLDddgcXRXkQvw1w9P95DRnvLNjK
jsK2hnybAgFAHfJ7cPVLep6wbWWTEHJFVo8uvpRXm6kQe0QZhrQmB49kzVgA4Khae/9iLNaKJDDA
10QwsSXVsqd8ZxRGZ2eWtjE6FKfEtXOlzaTW9E0H5tvlkMrXNhAStKoXvRr5q6ojb8hDx9kyee1m
R6i9rTbVLvPder5823mnOkLW4yzWz7TXEM2onckRsb4HkoA3qiWrqfo8nUP0M+WZLiPkChbwARCn
ysQxk7ku+tVSEtIiZhLWawqbNXo3sZzOQXJY4VXq5vIpKVm2XHcQNVbgvrB/Sf8GF5tnivUCumEV
fcsHOWa/FedA6TB3HGh5F6m3/YJWA/2VEx6QPh7gETwr4yB3oPyNBKKdqLfTfY9CJP9Z36TvRa3A
lr99rfhDx49OVciGqlr8YpIhzCWI1fgNdXi52Ol0aauQiZyMBy/o2sF3YQgsxUdiirCnBykB+HZI
bGXFbmGW/YFN63jWJ2fuF3HRZwIRpg0zUg2Xfqh4DDnGQknJUi1UvLnu2MRrY48FvH5kk3GOQv5j
2n0OEUV6dAa9IOvxb0flK8MSbIfTgcxDUfYF3zZ/xX9M+y5xqvcrLVfk0sCr6n6S8xJyQbFSpuFd
L+muc+BwTleDTOJuC/0nD0Og0eEWghjJfkF7jXmQqLKLCUJ0XE8ypRbCJAHOmjQ6R+lem/W1irlc
/wELdx1MCsNaGxh0VQQVLTg370PWtsKmeiaZo5LmEW49slHc3UjmoY38gmHwyfby7ouzBcIJjd/s
qfaJBICFwXZvk8IPk7mr0bWPPpOIn/Skjw7eLJXJbox0qqTr+FlXr7b/2Ccw7BRH1R82f64yybh7
kCWkxHpmWPHDQDe85VCvUuk6tGWIqELBQSIs0rCd9PpCfy4L/skGHdEGbDVaWEkqWbxHU2pRgvaU
QQisAmvFvW4LmUF3+D5Um57BxZk99XVXyhYJPKy5aDfgZOF1tD+qqnpAK2mZRNsjWCi2XUBMcF/3
Gk/RuZj29SiyviYvLb2yzuZC5Of0sK0Indn10fn2mW8LuN0uEpjpTYCIKXAB1aqLF68xs2W9Q3GX
yFhleWkAs1cnQ/xoYau7Q25vy53Md5Uf2iEOC6q59oasUTqQrfnGeZDyndlwqbZj+R3Raag+bUS6
xknqMoilRd9dPRt0SJuX78BcK1l2AkqcAv/ZJrpwZysqI/251OI5M0iwv7id7igGgIEUcRTmAZQA
YofxXVYQLwaCT0fX01yY7P2Bv2wRIvjGupINAI2J8+eVxw7JhzEu1Sebp1P+F/uPUTqG1ER4Q+sR
mS2lOpotZIraQZKLkhUav41pSjPo7/RuuFvGgZ6+n1CA28HGFKHqzKMmTekjPNBt4tg4bAqbythh
tpJoW8u0xu7E73OlOqR2rySZHUCdM6cNoxdwWBReqHP3KzTGIkGc9X/yxiLZYGGedRx/tHutTCrG
c+UYQxN95CXQ+GySu4eQ3hSMjnaCOgLCCKTwYeqDqDtYMpowVCe/RNjCUzVFHkGGD0OW1cCNtzWY
YxIEFsULu4CAdn62v79BpXRfFBIzBE4gNu98Wxughz8S8YbpNSFSgV5jYHOSvHwYR+F3l60L4VCK
Lbxa/koHCRf0YvAhVTAuPyxQVUZSY6iJvxFzm+8Jnusd+/vhhLFrOKsTtYn/GQwNN4+CYdwUUnXf
Rq0tkoKd1cTpbHAAp+KksXK99Wx2OfVLpXpC0ISQVHqb5YneOiQXG+UXp1iSNvJF7KFFdSb2D71H
oSNhQLltIjezegj+WlY9NTbJl96fpAb9o9pTfYHOpEjbb8lhJkAKVFF99pvTW9BbheH1J1EXsmTK
jWcp6TA885yKMmN/7phCrcKFm6r99FnuGMCnbbmltE4M7SFLcja5e/PRSM7yAN4MckMLs0AlgEfT
fmOu/e4ztS3/TlG3j0DutSkDKwfwzHUIbER5ZNfKizkto+boKZUK0+pUOn6uDTxRG798I/JCz+WS
6Q3sa24qoDIVn833cX0PuFfqIidfePeFbUxSaoRfK3+6IZ7IxRxF/wpI4ayjY4isqFlpkanFUkWu
IMGfRiRfNgJg/WZOlXxH2ILa+QXH2Bot6eyCa7bfxJg5hXXRdh+w9Gf2vL+pQd586ye6RYXLjEKA
Mt5xl8VwkZX5Qbppi7LTkUhLUR8TzWF5SXHmu5T9+KeYdzd5RBcd7M3IrO4Z1xww88GL6pFEhTpV
pxwUK6dqrsc3ANXl5mW8XgvBiVzrw4NlQktqh4KwZnaxBWqdFE0CyRTRfZuPpGAJNJ0db0RwkImH
nJCGCmYum2mvmrfhZqfBgj44erui6E7Mw6eK9CYkBj0yhc/3/wGF6/d13VtngESgEYG8vTCuFkvf
4q76ymkSwqBI4fgLZp9jvnFbkVgYZx8qeUbR7MswPYaBb9YBmFprVTAGhEz47zGpQJgocTGm3gaB
VoRrcfBHzOweq0658BRKQ1ktvzS3mLIP054lncgltkYw59pnhoM8YEqBXBT6gZN1YeKT3nGyAZ/x
JXvogvncw6x6zhNCJrc4hHznRb6NU2AilGaPfruUlseGGSoSShjmG61tBfiQ21BuuM68ogV2tYYn
2rpUXTrX3Yz8q8swBMw6t53s8SZ80B972Bqb9baYIf293CI7pvaHcyaCKTfHWsgoLLLt4skeAIrh
ojqXl1zzKP0IvT2xAgH1gHbjHNqAza28OkwJTdapw/11FMnaGVaRA5dIeSMYS1ww9cAJ4LmrQKMc
VVApbNAGQyI+mZ+l0WYmt22xeYSkr3H4H8zmO+wU56Qa/F8A0bZTvTSnOSgcQq4y8yiUS9JA9MdB
reQIPDm7xHlGHKbbQcQUIZp+cisgOsePbbaTyHd8x02+chnznyQBHlPXmEWtlZ14kH615sF5Huu+
EeWEfqmdBn6FP5hFcGaJ4FBeCk5aa+HzbmxTE7nYnvwwb561rRb37pYTrv128UdV8rFA8hK7cGr/
88W4GgmwizH2ocnt18HAi8sLZmfndcNJ/J2P0p9WhKtm++yLMgFlaeOZXQhk6kNxUvCCQwZIVjvh
hsIVt7DcgOGr7O0a75mRoxZxzjiuEzekN8wu+0+y2zlsBq5ak2fvS6cZY5S+s+6j73iCEdDq6Bwq
Fq2sixu5SsqbkSwS+Fvt4uZ4Lz/N5jXKvTAdzumIDSzy4Yt89Wsy2OWzztgHry4uU8GRT7xm20ca
VCrb844htI5E0C7mHzhC2Ei+prTD/xCMCVwu7rdQbkmhFJg9JZQFX7SFaKfxSvbP+dGQMr64A0Ef
m95/N8WglHyFShGLWwl1g97PgSRLZ4Xb1ILrA6ojAvQ3VTykXQpkup6N6iArEVlQh2dwDrjr3wNj
zU51g8yD715dCUcInEaomU6f0GQtU8+2F/8bk+IRpcQS7hNtBeLw7tIMqNNgSv4FYfURn7qK2EMh
pVTu+E2sN1TYg/c/W8qujxJvEsLzhQ/chpO3qbEdldnBqSI2aW0WM7oGJaRLdM81ig+VfTVp3Nzp
qBGGZIP6WXspkB9UOuMSDPvXz0QzpvVq8e/qEMUQorWq4XCaKZTZMmr/C0uVW2HaFT11UWLJFIS3
YDyveHt++V/nLqfYlo0efEMWyiXJfVnNbfymPyEfEILZSOpUkjtl4ihy+aD4Gt6TVkNnj0zaDI5F
70Xx4KaQq72RkCybK+FQSv+bdbud4LL2zWKQ5DjKLdkClaodrMWRF38G6Hi7CVxkhUm7+50o7K2d
4lAdSMyFgXbRja5FtJ959n9Wg1RfkYxVxx3aIucTRL5zXjtefuuhiZKGSOe3eQe2IufF0KY/d7h2
uOV0FqN67Hgue4Bphj0AyChGsdddVHwdahNcYstqpB2W3CXqdkuFwj5Tk7PasQU+ON70EnJ9MihJ
G6Tn6L9VxQiaeqX+7BQjL/mNm2r/e8tmLbnJ8XHr4mZSQF7irLpqgo+6Fm635FgP2KHsR1uhNIn/
EfpGE10o92eCaMLzeuiGEW4ZxrgQr0RX75Bwzbtu8xxqGl0DM+GcpvkJ3bi2ttYwp9jvEdzcgoTd
/l4TrOq2UBMuO4RVB9dZB6lLo/cz5UQOiycirn59uK65sCbxhdm3AzJmQdqXqFezEq5EW2ThV+zz
b1mjrN3CaQOnfiimJN7/cLPS1UDv6Bly+btvMUQm+gmV6WMUC5p/Cmp4ktDxN/XoSwyBRN8rDVmn
g+O7kdfRrK5Md6v9A+XJWUcwR2Ajrv8dBwH9NZtktS7gIm8YuqTgQYVhBQcjYw8DfbllsTIiyRJL
sB6FinA/sfWHrY1jfRXK0HO0UXJn1fQWbPz8j0P57mpHhVIfiNTJavLhjb6UCO9qFd9+ADVtQ+B+
ASEQcnjjY4xzaeTfe7A9IdpmXWlyLWmof1xb+cWRn67vc6osMvgXs9p26z7Rzl47a/eBqv18ggSZ
KUIEXkvh7y59NNoj3fp5/3NS0ok2TSwb951bN1S4Ui/JlFonvaqlJqvQvVSCfi/K0gq9ggZFamK5
TZCc+oqzY7SsSjUd9faHZXRZ7OQf/cLOqrYovNZgbPqJbvhmmEeuv3EPTDRqTU9hCV0Nz6gBscVF
kWE0qzDNqh4LdA/J94PzKiPt/cQ3FpcmhQbrHNUxVotarsGDqWDErEuKOjcuqI9qTkGdpE3FmMZA
5WIDZh741DrKUiuq2JlEvgFOymUg26qyh7qPxMC8nnM6FSo3+yTvRS474VkFCx0aqORNlbYHCpGO
CFcuq5XGASjU4Mf9JhyuYeXFK75/9JJOdUtrXx9OpQYnfRRkqLYsHF9aT45Bgo6QaLTA7p+wqqge
S300BSvCoOKCYDxoP2RCBmoyfG6fYVNBrilqTxs13OUaJTYMpQjTX0yBg5oNIGRvRnEv2yEZicdz
2EV0bsrjjM9R+wgz03xzpgkUp879hL+v/BCV7FAAuAr/o+9+W83kgXTHdBKGTL4hDnHwE8uIDAB/
vRo9yYsdVczdNZFfW4YoSZmn2VL976ANU0Q3o2ffdjqy8wJ4RdeDoi/0aCpez6nLy2kkhoKJEgWd
9MMugdzKZDlBOqQycrGzbJiZL2frIY/MTzlWkQwmzwVE06X3V7Ejay92CydjzMI4qK2Rtx2fzlmN
/WrWAPbeDu51SoEtEPC3j+2tNMP2d3dVIl0OhlrxIbKOey0pIMC5U1PXU6B7LrwpS4Hhv8UFMQDz
XYpjLmVWiWyJw7pLecTHPhNDXY3HwXUAXoNECwApbOI/ry3Oqd4S5FNko28JrIllm+3jrVZPSM4Z
SvJnzyYsCarJgo1aXpNAoIzSRoPgSUu+ykbvkLxYsRpZlgjsRaghYLmZuKv77vurF9fXxIKoIBj/
S0PcXUpH0pH1BFz+8JRbOf27p79rFFdXsKqKNH4Gl2WsUWWxlDLRvqS2v9k/KZ7k///iPGOp20lg
9+PnFM67Kjv3CM8Vy2b2cKlyao7vpCNZjhYu58iDlS8v36pNNS8iTzf+835HUWc5SAYRcWESCIjC
nQOKmuNN04+MCST4+l4uiw3QF7deTJBLF8bt0Fcj4s1I9euLq6DmGWaBZ2h1cUlD8mo0MXVOFEge
TnUnlH9ebfPKhH8o1esQ6iBQJI+RvRvKdSneYypPv1/NKs6ZZcuPljxDsBNwxvsqc/ml27hfKXOM
+X5/vTehDSdR7+B7ShOu8tpBAmjyG8aPuMR28sfHe7jqVUZto9R2LxJQR7y/yPKtu7ZReSQPN7r1
kf5CxW5Fa7JXKyGvem9/mC1bUNtTRQEbQxgrwFsA93MLkGg/uzzLYic1STMVdYz5KClv/YiH/lUW
qfNsckf51fpv/f9cT1q4wAaW6rqpnk8LaRx8tCKwONuAHzv5aCeJm9quUuNH7L/6wNLtKik8QvgW
/mUePAG03eALcYNva6Nzu0swo9CndcI1I2XWqi2HrAkue2agBo07k5ZsUC3NnQuX718gx0Hnn+zp
hqk+5hDppViIoW/ardOVecmcn4L+1Em9vPzvXgxMEoq0VPhMzhyhtEzL6xckONYvSrNj6tDTbxny
m11Cwz3T5xz5MdECkWquopLfCE4S1Bfe/W42D48ClVx7vWmOJznOoEc3YwfeuqozQLo8AcM18mKC
UZjYmUDvDLJs8D6Us96BRbZq0j+c9KtvBMbpf3wYT7xMfAizdy+jrK4WFJj1uBjxEJrNKB1F0RaZ
EA8Q8/4T9glW+NVMX1MWylUWQ35wgebIYhdM26I8gVBelTIwUHqTIN+Ae5fmCp3dwgepZgnt1HeW
idjmd2dG1x4WpUdk1l4PqoBlEFRtmVQdArLtR/TAuwXc9S5D09bbeR4gUn4DxCf/Z3+hmG0BAaDM
kWymuKbvb7S2Pyy8XVcPI+xcJjeblvz6u0zNrIV4L6e/qE00B+i3BTaHtMlxYkPwa8z26HoSdb1B
mcRiZ74LeHjUBoPR4LWCH/oyuQVhfpqSpZJLLOSnqDvqTB5JmWH6utIjon4yMZV4LGl6SLmn+OJj
qOg4IOOfbdHh3FDtX+PdGDK7/+c8/UVRiP3aSIaNB5p0QkHxcJ0HX0bROa7VbOBJCir09KHDwijF
DuJJ2ugYGJO3rfhyWQwEozbciEwbMfD9atO38z9CuSdUsoh2KGouNHOJazi4JsHkGGKf2AqFRu+V
6bbzdOnrxugPj/8dNnNfjhjZ47rtGilNLLwczfTIUULeoIa/FdgKT3ItXD+y8y0RTaB4ivYsbk1j
Jdly1lmobTjNsbWY9/ypsTGrnjj6iM8d4m3jFGDH4QEf7h+8h+8YUP3gU+g3CfeXVFYN3I8jneui
DM73Ms4sAbcuBW+ikft5qWcLu27fYVKyBKDmTNWjtcigxgJ8IT6p/5MoqnX0MHSULDCXV2kgTggo
oHDtiPICpnFju030HES/TjpxwxXmVn5cvIRNXpNhKi2LQbNf1qlSRWxQ487ZUbIaADOp1XT8DoQI
QhpTRk7mAoMZ9Jq1jGLm1fbNmKKA26rhGlCor4+mt1NXe0S8Nu2XfJ1OaMbGBy5Jo8y/nc7HGY4G
lB5NOojWVLCxCRRU2QsAMZolxMPncQnFOR8PStkYQOC4AHslQpB7a+Ql7wSf8FwpEzMdmCnzK7AM
DUkMj7oRpGVAiHs+ILrxKEaf1rDJJ0B7c+7SejisUw/7/6qmBKGbxAHz+E/E3VP2i55gZc1u/6Dy
eOOE4fzj7V3hR+CnPS6tx3olVww66yEdRq+hagaA8U6lYgN45tpfdJVRCdulAhWKsXumvXR0fJ/h
BU2rdKXkKAyhKgBnPg6Ju57Z1H1m36sRz2kT+ku+zZ7f3a6y6cTOY4VFE94OhLzms3+34MaJbu2+
LbGFWh/4xL/Jf0+ZD0C7fFe5oql2FnnUo5hOu/JAY6iGvLkP9IsUmx9qPea3ylBwO1tqZ3TdSMf0
Xah2qC4o25oVuh0MBeZN0+CYd4K60DRYb+OqOkYOMOU2H6VjG1VEPi28gwrK5WOUq0unN/T5zo9v
hQwhutREc/xCH3yPKdjVurRWmzg67f69FV/Va6R3uiAFZHxmBPOHHXVyVht1vKNRD4Jrq3YnupET
Va7pRMApb2q/UGWUktkcErrJXJr05DkO/2Ht+cm5R0JOaKZD0rGn/TqL7Eb9xzs4MG8EU0UUqXMV
CBTOrm12WxP9/Db0rCTyC0YFNPqR0jROX4F/8hFFH2mN67GRaqR7L8KqYqre0JxaWlDR0KbTjkr9
pfLoRFGoNommZ8CAIJLto2cmHBvKf51fmR7hXcfqRiaMsvJ8J1A0S+RIoRdbVFdLWlL9yTOhR4v/
zM8aYF/79nMkxfV0BDEIyyHx31m6WQfKwDxXHf6eMPLwYriaaRqRIozyY+fhWOcHidB3D7kvEmrb
D0Hk+Wgr/JRti+zCXtV8nrsGkhzGRnn/c45qOi6uc6Ag0syYDWAjtmSkAe8HXA6LjeYoYLAwwXIJ
0jYmkGiCFOiezC1M3vZtHgFBWpLFnXs9qwDwl0S5feLMdzxtfq5yyxdIvUbm0k/BATvwKkc6cDaA
7+F9Tr+5OohaMG2xycMA+MBjSMSIMkvvZOZzksNvcCmuNwjcLIIi0qXaO9xFolioqiVfcfDwUSwz
hyS3P/ixSOyFu0Bgvz2dXscK5rY/wMByCTjYwsca7AAnzDXU2BvR7JQYMiYIi6vYHo5YIX1TdFMB
kALNf1XRekKDPLs8kO6UjFEGawvuvVciOnCVIecL07oorst9OJDHhi5VahfmR6KRLE7IjHFUROd8
FHFmKbHSPpoi8TVqAszzkx/LPg/9ywOBjZZQV3TAmgsmw9lhERwJ+AcESHuaXzAeitTBN8eZ7/st
pgv0Hgo+U/OOQWKL9JWoghf7vYxrSFACj88Td8wDGiPLwVic7i0gepu9la3le1+jPQ4rfWHCUkGU
jfyO60ScePFOL0BvMMxgWickSvj+89uqZz2ByyQU7KZgNKCyrRPrIyw/K8NqdCilhB0aV1IU0LPB
wCWMrURuWfhTExFRKB4u4xpu46+5uTSvXUc8nxTxz8yInoK5aZuOtsHts9mnPsjdqzvH3B2kQS+C
n4/V24XgF2z35VvgPhym+ILWCUcFL2x0woUi3tiZt5V14KMPaNeKQgII3cLex+6UNEP2h0Er7Uzi
tOtZQj6467MOyyuhSryKHnf0wOsoJRFYVchm6sC/cWZdkh+EtUE89oLApYpleLtkNN9lHjxyj2XU
aUdUjTImZDiTgTLXUp1ffe5DKDS50r0MYRrBocpgkCX3FmrDoX0fZevJWY8i3kkhlkSD4Kbnj1lm
QrP5H4/N+HbhYVLyHOpW1gdwb0Rxav0oQOuURFDlp/1eCAXuJbqxp821d/3G21LnnGeIP1zpyEnk
m8geReRiO3lpzjG7Iav2e0tUbEqs4A/jqELuad13OG+p4pP4kiITPoJoY3h1ZfeQsPql8KJPVL4t
Y4dO5KOwCJAAnfWQAK0Qp3TuixMXMN/Kdb3YO7uoFbuMhgI7gb+oIh2Pqr9u6fQKNirAkrOi6PU/
VoxMIAQaQMQFi3M2zGZ3sgsAN+ResPuCtuPdXFsH1lGJ2mnYg6Y+3BS2nTT7IRFaebkbue+ZahG/
7pzRq1wKhuuapk6jvrTKth8TV0cJmhWpA8YtSr8Q6Vpu4RVi8bH7DQ5dvtOjmzd1dRU9sbcH6WRB
P1AiB3a9NtEW3cPPDMFyk84ZINVI83UMJzkJ7m/gCeAZp1XsWMitnmd/3yJNKja64OIkrEHqyR1F
DxRYd/B7kldekSGQgbBgGevLsUrhKquJXuxwIukyVsUIUTqdtEPnTS7i3aFSPBcfHFKpL0Yf83uU
v2TEB298+U+OU6ToXEvlD8vNGDUYaj45Btk+TaH8XAIyKgplV4Nfm35HKCuChQpS2qHQWasWi+Im
tMPRnDovCSGNfMqsIMgYhSibFwjH7GA9akPN4K7pero56Mh9BOVcMy44vrqvIs6QhbxKQtpQnwRY
IpYdeDotDMTB/Fd00rkrVkFW42XqOSBB/kVueRl+R0PZGFYX27h6TjcqV2Z3LqAuR6oW+ft5yLhZ
1dGzLzv21KgB02UVGBUP9TGazU82jlfzUKQjxSTAPJszOMtlWctlBNerpIbgLu/UOuxLG7eBkzsU
VD+GHFhTBg+qK56ktAYB/4GIQ/vum42E9+8f8NGhImNuyBGRPp3dzEnmKg0BQ1sJaSGWnaMFOYAm
5JxJtUjan+GiPlVakN+Y8/2oS37sL+Y1Xr5HFxUBeSfa8BMTZ0dd+TZiLmb+dOr41Ey5Vm80Ds24
bi9hZXvtu4RGKBrY5K7I7gT7XlXnJOY7C9o5f3T6Y6YB8ikyJeQNSgTI01etRaMeAR9qz0kjcu/O
IIaOhP6b/5Jlhx+N6O1ZU23BpFBT2KcfMTAgH839ysTyZJ1NEs7U8TQpZ7mVB2hjlUgkJPlt1Koz
KmOhmydikRwCxS/ciyncjOWFtshul0OhNvo0YuMqv9eFwYAR5zOEwsfzRNqsDaUGPje7whmqPJ2S
k0ZdDT6g+LXsNWSEmr9C3PVjOWc/umoetGlJzgbPrIPUngm0pxGNxdJnP0W+WtsB9GD8yb0lu/yc
TvLu6GfahlUYbmgKE8qXSAPs02lYlLdC6Hu8JDK/SnPzW3+fc5wEK6ZMYT6qbotA0+8t0c1Wskxr
UEgHO3xuPJGZsgV9RsiyeVOtrqsr3Tidi4iIbdH9vy+15fCuYRSA2DL8UrK1D/4KvlSw/PZvKB+j
kPlOcfpI7Kejth5l/mumb1D8RNB7ulIqV3w4PKfQtWlF+86NNajWy2L6l5LBoTvdq81RRoVLwma9
f6+BS7Yer/GjKFZ1V1ZZ2YEaGi4Jc2pQpQqRTLe0l1MJ/eJyJ5MdfZeGDZcNNKw/xq5q3E/AAw8/
PzNHkFQ85bxiNTX4WTjQcEjhW7rVT4tlvPfbQVTcamPYyBmSpVlfIUJzqgmXEg66Q48MgGSW/EaL
Lnf+MqGCBszNOvlFlCWbgUqAoTj4JQG+mEYv6DaEjtVvjbSkDb175Tlhi5bUtC7XIrUV67ut7nrP
+t2tB+6Tv9pAi4L+7VBn4mp7UqoD5wpoXZlFVTMrt5tmKhrCSPDfv3SrW+1j3Tuw6lanOM6w1aa4
iTL2PlhvPTou8U0PYk6IXB37BVLqAzGEwLDBmBOCni8sjRMn1Z77c7bJYdBNff5B7TWX74W8QcAT
Jo8kFo1JDEPGm7zwFWy7m+1BWHEFKs+W5UbXgXjrUZmNhWS16tsiQvO39ue0D94dSuTp9DYBeC+E
KxW51z/J9ASZBasF+30HpurDv81QPLrGy5/2XAiS9amdw2g94r/ELyP8sgNnoojvKdzH0YBA7Vhg
f7wFPA5qy9k/T+MUr/ka7s+4tP9GkgVbGt1/gu/lpq+o4LlA1ayC4LuBB2P1rXAcpcGfgMOiu8ni
dfsLZEcpBlvh36pIVBXJNZXKtuxaNLaK3Tjps1Uipk1opILoQ+n5tVHlNY3X20gOSRBSDqNWFMia
5ceWdW/u6jcLLSwx/IajXYM999GyDseS9H+iLf0sk66Es+IB6w2fzKZDO5T4zpwen+1OQC6jkQQO
99+HGbucQuOydl0UBxwxbic1eprZBPYI+/+yBhsntho4Tr1zbqXiNjgdBLCnC2I+i1/Hz3brnSnL
dT1Qjo4exO+bm4TSlkeCYIZnA7Bob7B53G0jlOIRGzZLX7MQhiAFvEkYlbw3C7kK0obvn7QgBAEF
HIwpu1qv45stesa+4sUEAcMnap9bSGrKW40Hj3FyNYgQNawuBzpUA2ewrPBGlAPURvfdm2+8wssR
zWGHPuf+rUkXJWWuvPgzJ74ySbZxu/EXe96LNpZL3ifhHdg3j7KlX3PDGwQDLe5woB1yMizdCfGi
M5LPYgKguCWKlM4TRH4mWn/gV4xSPiyYgs2okoTRe781v+T13Bi7hrr/z45kmENCiTn27auZRg7Q
z7S4/W2PNmtLDS/fI70IlSHB5AoHdv8KOOib3WvQhd28HdDgSyA6yjQ4dKplOvMsPeNBXpw8jtKH
H6IE0myjmAOfm2kaz5pLzJwi9OAexop2lFzKbk/4CMcy3FSm094wa1r+bbovtHc72u1Mt2ppmo7O
ioAAf238oQERkxE89z6iOV04Ltq68KTOY5/kR9gm3V6CiXX3YEgh/jEXKf6AUG+7n9SdSQ7YaNR4
DBYRvqSd0GKa29OvnDSnSmI+6bJJ1U++efH/44D5f7+tc1K8oIzs4uzYuHiSjhc+DmBlDxuC+Wf+
sUBDmEgVncuXkH1H8ELIJnfpVcBPFO0R9j6kUXhVXBS+Xwogt2YfJljQitj6tvbDng4SAcoBxcpe
YPzaLianeJHo1/tfulNt1rsAGTTv0dQx9njWYqLNhzswx411S3Rl4HSkfKhGt+85DrpJkYprdq8X
K4igLkNnsT7DGFbdHQ4SlD0OsLAivkyVrhHpKVbprAIEFk/vE+ZR09c2nIqpnCWQADHRy8WCy9HN
RgOvHnL1KhcpSIcTiSx2ssX4KR/duAo/5kqK18TkYzrj3WfVXQeL0Jmf8asl93oAnYTXiJoIxVnB
IOceZPmekLCi2ti15v2MenzAtxb6i5H/bUN+D7wXkpx+Clz9lX93ga9X5Xpkpdu/LVaPd8PJQbuF
0uSzltb9vnJ/iMKb7AAYHodI3PGZgCizCuFs55gyZShctaWeOoUlGvY0e1hqzyCcUeJx8l/JE/Hb
zAkaE3fzevZvD8G/VDYqTSK/QVDtUXqiNlUnipJn42UHL80D6WXbzJvGfvaQ/fwO6aUG6y+sz7UN
hbjPvHSLFSE/TlqWnc76Zg1CmNRgc4SJCP2z4XoTTNveo0ls2zLeNjKEt9TPBwRGUy1Nfswh7M+f
3/vYnJWVi7ESO9KJQ2MB3FrMRvR5aIvs39toAEcgs6KLMLvkdgTyYZwHNvr/1NpfQNvs6bavDV2P
PCmykhQXnCzJ8hSE2FHkwOrTVSpzym1SNR8neKm+VNrx4vTUDVLZspT7nkfSAozw2jL3AO64/cNl
yzmXbOj0eTwc8LY5XdWu5nJel9yvr1dUwj9ceyPYJJ3LRWueCXOx+FrfQxT4ja9hZJ0ibWKIvyCN
+XW2EEXuB8QjovYYGjmFQQUwJVmpWacrt5V1OuieSMQrAak6AY6QIs1ubOPXbbPaxtv9viat6FO2
C0Tpo0Vqyj1aU1RPxIOFZ+ePlyz+7KFMiaZwVzLWau1k8Tpg7VENhslQJWCtxOoEW3/0XpijiVkd
eGzTEQPqnk0lwkozNp7e5+LNxo73yPM1sChqh+IAeUlhRz88j2eYFmALTZU0Z2hlO8TlVO/1Pb6f
KesFXPN4aQO4GjykxCIr6t7HGzKzeg3PVxL0LerdrOkd5uPd8Vdurf+Ezbv0K32dGlfy4ca+6rVl
Tm2qhEoWAF4U39unPBshSY1thXPcRBMMdIWBa/5vPtlnb9k6zYVE6nHk6BzlCdUJSzxnE5jBGAOt
gX8S4wRoMmKmBMTJRMAzNsF/OTCXTMfkBSpn1KjFIIbWmCVUrHIHswCeg3c5jQlUJhLdKUGzNRGQ
HIxlxK1Lg5LZs0HAJcSEizBp8QYMyXIAMm4VW8FpmgKR938WfcpeUNB3bWLjxGciy5NWKRvZ+Cn+
QskJfz8A0+7jOP4YiPZxu9Ao6oXqBwa5z9LVAr7I0o6I2HXUEVchGRxiwiLS/WQSZ0TEM2ksn10Y
QTJ9awc/k/OwlHQyPJwalF53tV9hHCBpQmDK4TSlWMyVdT8PMXCLymx2+l9ZpUJ4+1GkLZfLZpF5
7hKXnwVky1Utq0Uu7rY1iIPHuu2jPd/sr3zqfnLInCXNZ7WhRxck1u4WrmIOysYPLbM8PUarCbqM
e00Phc9Zdwigq3K+Bq34jEvDNYfcx/G6jfo/01ikVaFtjupj+1+SekKH0MmhKMiKCJDoXSozA/P8
V3GkedamcgwpQYIf2SxsMFHr3C40DLDAl45+Pcw6C3H4ZMDA6N5lBTzYk9ri8d3pmwenc9UOokKM
HQkoW3/dFMCr9o6FquauwrquBI+RhPHlIQIQ1XOwoxuIdJJy1iXHLlEjaGG9A8aGeQcG6ZRIgZxO
DzsV04TZMhnZNMxZooDIbniNR8lRF4EnLNlXg0Gf/G3ASKidzZ500Imt8tLKU50HsUTNY3T3+E2T
WgYlljQrXYjBHljv2VFAgu/WNDiw3ADb74LmDgu67/UjKXfD57bj37h5g1vxSLhGx8Xnx89ZHSTW
W8XRRnJeOlXfTAbiVgsLR+aud7ycMywm5uTlR4cgESTTaHiyi2EG7TVku389C5I5DNvvQDLg+2kn
f/9HSHkpRBq4hYs6Qr2TlEedzvyCuV+2frL+D6VBBxmpqVbKPBV/gGOvbc4RFb3nEonlJW26XO1s
i2MpQBE+shnXSbHu5O0/gwWDQUelNWiHsgArllBMPPiSJfX2MwwXLh+lf0Txor/amNekpRVIPbDH
+JbgtUMBegmEPJfe7eLSSCZYBHg5ZtsuuYf1hFmQLvDah8+QXAmrQEDkwJIAJ18KDV+d9xOYjppU
T9wtuIg5tD9O1/W9OL1EmL2F/JI8G2QIDQUEEIL9WGRpq6FFKzRFr669HFJuXyWwgUGsgp+m7vQB
bnZs69mohkPRG+kdRD6JaDDPe0aJf3mYC8uJvOlxMa5VslQmG1fd2wVfP2gjfPF8Cvf+tT2y4vJW
VVa5Alg7Ntjof4zb7v2AgrHYVhP4Y7clHoId+t1p2MSBICFz6aGCmhRAgEMdx//xUdd3FGRprIHD
3Mi87K4e/uXsmGIUZaR7bCW4HYoyI6zpEYtnLL2ua5nPhAzyEdlTMnQuOeVEWtj2W1KVDy0mokYC
k52wXD/LciGgarR/vehowXRFqPyXf7/zNDITUdquIEmEiXdCxka9mUCogf2tv0OPDaRXlMDdjLFx
wJYi/nPCjzXbYkr3KfmgV3tbHGk+V8YiPT2DazA5QFG/jFikW5utNAHGSHDgrOuQd0JCtSLIqKjp
t7amvbaNNC8MIvYck2R7zHoW7VigjknIdfbmYb2JAq1VsH9+P0ccaWxzUAaZuSPZmbQmWcfI1FHv
KdapTIxWYTsdYtBOADlin2P8X5qMPv0UJ+s38Iouf2U+BF+2v497h0hrVGtkMB/BGUrIv9ZWD6uU
YvuY85oUMFjxdgQESTMz+vf7LRFTgw2IRy6dpJCGd4iVyXEBJiZC2/ovOEwQ7av9Nu9FYhAFKabl
/GzX9IlucDmnCJV6qwZcpIwbUMqaGOQOuDr7SnVKPSUdTWHc1+I1WODXfC8lz02+hxpQHIayZ4j6
HWrKw+/1fGsjwQeG9b42P/X9XwM9/JUSIgcAW+PlPAw+WBHbkryDhiNvMgMXsyxrsYluAHtNLSxg
JSbYtmQ2UhqavydFB1ZDlBXitmCCNUd7K/jaJOO06BgcL0yVZBVCAv+ean45jv8zwQHCZQzTcjPc
2fP22Yz/3Meq+onGNVLNQWCRvGrzQd8+7PmSOEaNQloqm/TjO3rEWZcpVNQmdniofaPEBXrIDxxC
/mQOUhv+536pBUhCz2m3FNbQKTSYl9Vn05nboilneCucIYFf9TJjQjmo5vWg2GxewhHgZXNjaeDA
pFEGgPUKW99W3wUCpguxdiycJuW7HI9l189kfsjAZ/pJ4PQYwL0x5h1A2zdUIQD8aSOL5iGkDTo5
Ih8PKx+bff3dKU85P4oEk8aJrM7/P9xsYL/oFPmKokl6qKb63EIWyrWUQmfl5seH802sD/kaDnsf
KSBNlY9kQvS/K73OZMqlED0domUzKYhKfWtou4g28iXWmPjrmz9oRdYwlNgwcili2TG7jkJz3Ue0
icUWjE2pqfT18CRMGyihU7yg7W3pZ0Y+cW1x4+hYX5eff9DSzNKRUPKG4YO5QXR8pM+lasUJnU0h
q/H94/+7DT/sV6wDzzIxyzhqiHQvZ2GMEnK3rB8w+nhI0ONn2Gil4hIcoiPWLRgufJir/3kpC9mR
XzuCcSLkiFsYQe4yR4JdAWvgRsUJnusfqfA1Gp9z9GJLzZy7ZJG/39+FF4de+whLCtoUfskkC4KI
dvgaaXzF4jfkwjfVIckSEGYacSIYgYPi0N/j/FBtoUejFWijroVUk2a+81KX8HGquTI8Ap/skdgB
1X5pim4o5AAjUjEddqjryTFxX+oJs263uq+PrcH+3V6huWBHOnUNL6Mr+XPLTlXVW9nqp+rogcKs
o83I7OpQniN5UudZfAVWRr4MuL9rPZop40cEY43vyP/uX5bpdAce23v4/LcMTQPxw0qhJYNPZZL/
3hHZSkQKWzjIymcTXsMpgIDRxL3UbMPfkBV4FGFo9xHVkfYHkN2CfYqGbA7TB3DVHjcLXEqvN+uY
JAJgPLb4op/0si2B6TgCWSsdvagYUZ3050AmbyTIHuZNYmLzKXHyY8RJoIaI7p1VsiWUH7hag/I6
Kx7wATs2mmKH9bfd1mXLYpZq4uUfHnhwSbcXI58I+lz9/XHha35kiv+/tFGyoKjF9aNi42nDL/tA
kdYHyT3X/TzE2dkXbaSC2hszWJfunjHVSe0lUIozwim8/K0QVorJZt5rIgIkvFFuVNlL7IhJ9CiR
SweD3QEj09cDL/3198Bym7JvVqIHXCH3RSZ6jILlNMuu2ZtzesgczK1149aagCqCAjSFxblULuWI
AEV7OpS1M+u9Vl9nuOBXhAydqEotpWi6ntIMuRwEQVe7NWsFnyYa8jE3l7y0iMrbh1FCg5xzt3iK
OqNyJVRu8964pLXPutH+t/OKvbX5tqeuSXbbgF4oukNQoVoeE2AMPqPqoZFcc3mspXEyERKolaG+
+YvD50muo93Ke5OeXPNZ1ooKAPtAh3L3R1pext5NpUoBIb6Q9kQG5PSBCxQVRcwKMiJgxneHJTbs
6tBneshfMtpuQUcgVO9lsyYgMDsz61jYz7aYdmCDDOOfOJfDFDUFq87BGIje/TgJH4607tUcscy/
bJAJlKWcwJVAbgIQ+sJCYS/hfCUhJQapVm2wQxPjotCeepydCP2jIFb0fVxbWrXNFk2XlpJClSBK
Gzm7Hrwk3r/bp3Q3qER29c4dMmVIm8cyMM5aSfVfF5VrnobebCe2OsDzllrRQL3drVRtGAGSsOsw
qce2+FuS6J2UYeRKaD1i2E+l72F6Xx2OW1/pZEC1SeaL1BhOsRlruTIKwjvPn3jrbA59yg4L0r9Y
/9e9YXp1j15EZHbiv+k1Zab/E15Vk8m6i7q3JTr/82q8CQz/aQSSOjuoc/DxqnWs/SFoAYCjxOqB
iQqmjeWaMg36t5rZCkLXpvMm4yl/n25pIfpULzV+YQh1jNOOy657yekHQlfeLtqcl00C/2qyJTk7
ht+P9Gs2Og5muI1zhyh1VrBnAMiIEv+Pggxf0ZeoCPP5S7RDmi2nuqxAnQd7sYdeldIjTPAS2IJr
bDS5sQuNerMeXL1yDv2ZJ2UY6OEcIKQEheOVaKRxZ4PeHX1tTx7xevBibndHkiNPlp1Alwjp00Qe
+/rz5m4j6nFcCq+E/06xGS9tlATRFHoPi+k7XPb46mBWrxh+LTTrLk7Hjfj+6/h5SnRCPYjzx20N
yj9+y2p6fPZRd90PeMjAdHnuNW50hj/6lzMPrkSX9vXP0A2lw/1R6dLIQE0N1VE6WlmYVeVSZITG
gUjw3iAm+ywDddLhhQJX6yyXVH8PxW9mmFWCWwi3Z9a9WkPcJ4VWOoZ9Hfmh8qHL5odNpqu6FXHG
rbWY5CIR91m9uKxqzOAwrgOni8QXDwPu6fCY2BOfTQYSLYqzVhlbcUzjrUUN1koPjEqFNVZXvToe
ZV7lvLlWH7QXlvrB7OHKk8u+66jT3Ak6AWtOHLodY97nWlm9Zd4Do8sNThJp0lSML+aT65Kvcrqe
6svZocmoAJCbWD/hwI0ao/sQ7Po91V9KJmH4I/x0AzrJvkv89IylK1Ah2fUsJZPFKWiZo0GCvWRR
z4k7GpbLH8XX1EncYD2GdSxRoM/OMJ3KHAFVUN/Cc2vYaPfUzxFn6XdKYj1Loc3E19VaDlT0byiK
aTrI1fU7G2G4mxW2ViaGSNYkyyIiVUwivxJdd0QUgU+FhBHGeoKUlj7a1/ew2aXybiY5EvqSJ8dl
OQs3+5XAIAlDiYGqd3Iz5AQS1s1AZzxXbPH7aUs870YvblKN0fMtho/P0CAyCGSAiz0/SbFg5BAH
20rMTKt1xA5ycGZx7ennG9eqsOVtFQDIvKC6TbdmQNd69gI9sGNyDZAKXgqDkUhie2f7BqrlKhuU
lSWYSmqfklJPHyozEnLXOuW7Q2WPFEeOTjVxq3+5MXK5lky540hgNwaZ9rkT9pyh0PbnRvXtWgfJ
f+fVxANMUyM5ysgQDrlIFNRSxQOkp9NMmwXqkd5PrHskV738NuA+o1Ft9UFt3vOG/FmPD+zqSPS3
YfgKj+5Azd8YpZHKwSo6tF7jhf46h0dny2/+11E4A/toGNZuE5YFkyvaTb61Nyx4HOjjyYjiB1qK
xStQSupLsgjO9mTIRCWqxYM94CBdLDLkl42HWQEVZw5iLuQW+yeP8Mih3BbayQpKqnsNEFWEf0KG
O1ow1qyEZpg2v/r10pUAnKpWl3JLi3tvPc9MHtk+UvLpTWYq+MHJU6tFYOOEzWqNRLJ9fiRNXL4B
nlRFxJ33HiSip8ZeeVuyo18t4nMidMxI5kgKrQqPUicDzpIMokFubwxSt3rpSXoa1YUso3v+XlU5
wh71os6/nX+crCOZfanlvVnxu9KqSbs7xJqpcXjUGxCNFRQhyWuFKFdbBfsAvL3PzedMCPvUXAPy
P5BlpN3XRKRkOKaqO6mSwSzCrImtfiC+EtKfmRpzmpr+W253NvjNp4ei1QKRivpxF+QfN7Zq3fGI
r4ggIC7d0QHECGIou0yK00kxQmQNGrSqKO91+y3r320DWb11kzPRUmOVtE+4KVXEPzV/2LrUvCau
TzAsxNi1vHc8Oalq4uNJbVyQnju96i/SJ4x14CBc5TpbAifI03qpOn+iyxusLc6AglSy0rnOaXqE
i7MVYIv9SBlQS5HbXT5uDknyaIXtAuw9LfHWlbw0QUySo1UbNWE1FsvrOxeWeU/SP7PM/8UbuZv/
L3mgKeMCYd1yUg2SdXSPMp4Oy4F2IDd73ZKXYIfxJIED0AsvxRRZy6OaoXRVqDCuD4gd27sjUyMI
OHPL8ZldCuOl0iN+20/w+0gUYm2rv0cjJivHhHUvk3GTtEoa0iNN1QsWEmwzHuc+9lpjXZrIzgio
4g2+DmcYs/Ok4Xo2jSTAUrj649OhkfjRIrw2e0mQa20jfpWB11hkJ3njT/d8SnrFgdsvpoltDqGt
nbRsIOkvDrXbEuciQAptCVXoLeePzLhYxylg6SRlaRomtvJ6i3MgUWINeJo6MFOoPxPoAxLvuyLQ
ecFvExF14E1NQzRnVoaL7i236d0r7XV5w7dEdj5rlPnlUDRbvWKg0ehHnms2HBfUw8qsjNz1P/lM
52SUP+oS1b8lR4/t6Gbx58H+HXNxgK5sY8s4+UVXkbrcdOl8WFY22HXQcsbTAN+GJw+WWOXI5D9j
23L492zU2g7kxtmYH3ezaQElTeXCRpCL5vlQrWlNW6Q4qPVa5BOjq5A6JKs5GTh03ThhsrFjshpV
GggeiWr9m8uDbWgJgCagxtGBndV5axnvDbCGHDSeBGbrX7UsDgMh7u6K6AiYbBUR9ZBrlEjmtB0O
afWo1TyQVEjgKA5fEsC7m0U83R399CAmeJH18S0wrYIQewm3XxwRdXoaeBnuh7WVSn/xuk1q0Fnn
nnX88Wnp0KndKa0OfBSrAgmqEUt6ZTiGf4fv1kQGpl5lC4XuBUjYZ+5XTwe8bbS/chfvhZ4hSrqU
NglyQXBYjIaEfnT7Oy52/x20fkqYBQyWhNMjWAf63IuYptZ+CObnuUlrkdQNuxMUIyxWSnrxl6ho
D2rwtuqIb0XIZl8F13lbFDv+iGhn7z45givLZTVjCfcHFVODQZX6qgYZCWRKoGO0ncricIoUHall
+FJubygTOT1qTVSMAQmB59h7tp1Hb3c8oYScYQtgp+Wdb+59gL0Rh7L5s/w+YVVsw915UT/cC8OP
NzmQ8SgzYVL9Rzj6UnMxr2RTBZmM9hPUJ+/qXa0SC5D8alLCP7UhDVIrVyaLRiOQ7bVYMKoBRpxA
pNiinlpJ9/ScuTyAMnY/VORt1giyL3aHsLkAtp9cFkWXveb31jHlMZq1A9cpVgKsD++wJWN1Cwdz
OBgmgXlf9SdoY0T6emLM2M+bBYVgME01lylvmEKnZN6c//+j3wKnJAOITyJ+OHHaIMDgu9XUdCtT
AzHDYTdCVxoDZimzjWR32BE8oksf+sgZ8JvADO8QI8pgVz1ejz2CVx76aJiWm5bUJffT7zPmMUYb
nvH21s573DtrYShAEA9gdfjzc7rB0sIhKojXygguru22n8KpmnRTXOiKTyAi8eX+kmnOgVDxvQg1
veF2PAcbdLeBQ4V+78hG/stKcVboS1XQVjrLduAD5P0eQ/ERM4V8EVJDWGYWhsfj1bTpxTe49k2I
qtEs40NXPJ9/jlT9ainx/TtZxLbFvAljdZiD0p1Feb6b0w6O8/VnpHhun/N4FkWvWiDFDtktyDAq
Py8dPCiU28FSZg4gGApxtTySc6B2gkaG3IT9DJikh29RhPCOwGbl6EZqTTalm13LPpbLg35QO1y5
OK/b502BNuBSHHDwYBn70mPrvzMyk9QCPCo4Dbwkdp6p7IUfC85qC9IHSAOu1be5fsHalPI5S5pa
aWjpnjUuSs9hYPBbqov/U4YR82jW4hfAy+0x4N1airgvM2LrfYkmOJjCkgyFcjkqQvG70h+CQ0Kz
TpHZXhorwKuW6dxF6PAlTEZaT/ODXB2e6jLP1BT03dJbl1pz2HTjDdhzdva1gVLILjxFEaHmxh85
x/2icgum38c0idhFdsMtiNaSy1E7n/MIV5jKRwGMfhDzsgl4FyNp0gqo5RQmnJtn2IfvR7JnyGzX
OKb2GbBsPhbb6Ac3J12AncmxywBUapoP9UxEikEIWB5rD8wVthHId91vyA58ke+r4vaWti9diyTp
PLkjurcCOHb4rJN5UIHQ5K3V02IhU3Z+OxhpQA0GT7FWBTId4BI4EQ3IPVSpP0bk+hJYtG0CSAOo
A8JV2V4+cgTPeRvkzA+8s5As4ihiYckCnXGUwcEMPJXxau3rmy/QwB48XAT0/zGVjphOKbWAD0ty
A+Dg8l2j81uzBUQubk22lMwno8yItEJG0rR0ZYXqDefz5rwk2KWqQKyZ5XKsg40nRJv+LgZMrc/h
4Bk/6ZJf06iuxkYHHCzYHmMM4dlnk30M6PKbsoK03fEFNT36G1eOltn4UPrwC/DzwwHEHB1VBTw/
J0RfoNZ1rOQG2+nPbl17Y/C2nCHhdr5TNyY62XjhiTT4fF0qgJso5wW+W6O+0GrYDs2b5R6sEhw4
1kcnTo6Sqm0Ki4Ds8MMt53w6qCUfLkFIvLXPTdilkNwOgDWdBVUWE79Lfr2j6VrZuGWdGWNkeCLQ
ua3inV8MaF27tFW2RjYxR8udKLILxsrczVdAfYd5rx6ST7YukP8aMsnZdBSm04f3XifL4AOJDKFS
WJfVkkDq3cFJILuE0A3u8CDJVKGPylz0epMXWx6kZj/xkD5oZsKPTwXMMX5PDzBqAmHOAKgdq0y9
T7+Hreh7Oph8mC338m4R/01TYwd662+CdMTMUqAXbm6yGkkIKu3NwcyrtdDCpWK/cUoBxJRBcl0c
AQfNysrTNNuFnDf5t8IE0A1ahYDzj9S7eET7XQgLhyhmvDs8gUvOH/Kuvrc/eHk/+gXxBGRG01FH
mVzETqkcA/KOfhNs8DK8vYUegxZMoRLaimE2FkZzd7JUFBMOe3K9sqyzbL1pQJZcBSYu2vGUJbZ3
rpsemGYRvovuZ363SEyr3F1z24A35sMJsbZx4v43MMOlsqs2dN3uMB9DizkLstw6CxEoolx4mPUO
BhgPcvCSj4X5KapCPnVC2V3OzCcm0AvGGWhnBS0bMhkrSLle6dMilLnD+NV5qmx+LJ5tg8FJlDhd
P8wKvnqtXXV7i4c8AY2xG7MUjn46y5r+W8kfq5f+98v1tRikI1za5wT3QXoxzOm4q6juP3Uinz1y
sTDhLt3Hvpn/W1n7wx3D6V3eZZsKErjLINMH24NlNrIAPrXSOPP28y8G5ESN8svRDV3bJrwFN7To
2Y5XKc8bjEV253lfqXCEkf7L7A0+wNHBGDu36Kzi/cyUnyu3JEmbiL124na1Da0xN0IUenUG6EB6
ggcJMnaIFI2kEaaVzX0KJn3Ag5J3XLnvEzg6cUeVeUwDRIdTUd8TjygROHxcTpyOHGp/rUdQ7pe7
gLh9bqIHgSBDMxocYGpssaEFqnqqmYkCD0PNfY8P1sEPZWHtt8W4ADK2e867+pNx7KQAD6Lwdasp
Mqw2wWjfgaTsvF5GJIctZBHYc9ApKhT1DSjxssDBBz7lIs4qR2wRteRsJlNIM7w+hxjl4Vev73ys
5tuJqketagSesW+LMbQLuOn8dJw0I3FMUZD2biAYQrwrqsbQfCvRicxM0OBvsX9n8PNf3Z5xpqu6
WgzQ9XogQAB7LWJB2IDZiVnCIAy0fX3DKdahuWtDapN7R8yONW7KnA1K9S2XquvMVS+VV37RKSbB
YhBh7erEOQ9SKU8Q3BdJrNUu1hjb5ae4UieVaJLs9iJ8fyGpowk0k2yNewN2rCUVSPsfyuLTQ8xH
AcYI+3f1tvktKJ83VvSvpbIubswaYa5gvjEutpARW6opehgJTS/QlcKYvSZ7fmp7v0C2T/TCrcUv
B+zlHu0Qiik7u0VK15QXjs5QzYbqqS/0gyqQzs2Q2n8YetKKmqvAmfxpKr+rTyIzgfABcGAOwrSi
zY46h7hDiSwS1PJz1oj9uS+s9HNEc/MUyQ1clZ5TY0MLwGmgh/vq83938STtpeUWkUzSBwEGwMXV
yi8+Qb5VuQCMfdMOrYxPrA+bQjVvTgwKsQnnEGl74ybHFJ5O6sRj6YH6PowvvL4bVDAOGCDzRL+t
eQjwLQSEANLxhAoyZB/a0pcWHb/HnrLy9xM+LvjB/UbwBPRCr4Iby/rM4AAqCbfyv9XAxsUdiRRq
W1MdDe5hAa6qSbYPxYT9YLGw0q/3wmCv37EfAiFIkuYwuVmBqHkM+ZmPWjST/wWon1unZDAFNSz4
jeG4FfzpH95+1Y3cT8XiJI9p145DZJQ9p6wbNjANXZCbUTAIuvQWrm6NKR7poO4gXb5SR0GculSe
TgGB5eCxqK0HFYxx6j5RKWt2pwdxuiKz3E/81Tq1AKYBlYM2NJUPf/ag//xjvEwvGp1yybtDMQmB
1F7JF85w9aacAm7e3laqhd5V+Kv/1nK2d7ysj0T2C4BMQnQKwHj98m/amd6Tsdd6usE0zqu2uebt
/PL4AMo1lRD2VsCviTXpL3pIdXKi0bp1/i2fAIxNsRESZoMnnIOuvQyncloeshKeB5pk+/+6+uYL
BWk2E3v7AzhaCnWEz61Ce7U5CW9bxiuuGxYdpvRWGt0ugsoSy0jq+g37wkPUCOQw0DJ/A4jXKkQb
1ysRQIbMtADV4iom7wGSaT8EC8IvXAZOfE6c/w+2Ne91xSBnaUVoD2ikYw45mVr0kxSTwnWrFMBw
AJrebKqeyrtusOBFQ2q+3NcW3uP/8DWz0ZMB1RHYX0rtoyOtvFuzH8z2mMSnqOUaZHwMqnHOtPd0
HhOmsKsTDuxT9m4ESKdNcGJzO3ND9D73AnO0STGzW0NASG1L4BLjaRm9cGrHItqLm6p8GLckoIzo
429fRDzG1hWSzXB7ZWUhJa8DzDDVX9L1lNiXS+IuE8r6dIy+4ejw3SXzTlGFpPPEgcF5H8jpGGCD
GnAi3ggYUO0LY29/MAPQLXDd1bKcafAqGaJ9DWxyeaAh0DBZkIsarvZvw5AHqX6xKOpvqqOzIb1P
xheEzwPezZB7jzeYptEEzbZxqOA3dxJQ8dZr1CvKGCpmlfyrVto2nbhR0R4DCZYn1q/Q9VzO7uY7
P3agtdoEuwX9nVTX7ubl2coe7zOgjMaFptI27rKgXIZOENTMqgLC3mKvsQkQJ7XnqyCYX9pWiz2L
y1FgBq/kIgsP8k97yT9riHsySxViU/0DSmTU9cZKcx2DXVJpqjvs1RUsu0ZM9UPDuUSHBnWPAy7a
mVFkU5rC2DUJhgk1VOb2TtsrNdWLapJ7FxF1N1fTlSwxvwI8ehS6SIVrfeFBYGI02FPeXzsTt+TU
pEG1RUMxCWJgAKOi3LNLh2YC7bBWX4VTqIxRBOYEAU1/G4pO1gzKsyl+EE+Unr295MCz8hZ0uEPC
SKYib6OP45R13/IawzRZ6eMyIsKWsXsdu37pZ22ZpnnUHJQdAyGmH3bwjojDlRhTinmh8OS5aQjk
jJLvUTYla48Iqty9/nmETEE3tx59ZPRR/WGjJDcIn0mkbHdeXSSuV9u/x4/C0LTU26jPl8KjrhCt
0/Oo1HyPullX710s6eIHIUJyB8y1nWgU9phnfexg+dF2roCfvY5jlyYFccyOHc1DMofkrFQig0lq
9muGRZhqWIrCTZp/m3ZoZbmDusZx+fnFRpQJvUy8iGD0WbiHHu7eXoATGFaghIlrcQicj4FiPxF9
9+Ink4tj95buGEgrUrkkj6MiGP3eZ8sa7WWmWnwwjwXJ0cc1BQirE7v8EfpkB/KV9f06fF+JDa2l
y6ukZthL7z5YdnxAqCabbtElHE2aT58mAdzEKWrvwzx6Ni5ByfNk/Fzz+chRzSKVXB9SspsslX5S
/Tc9PB6hLAsAd4QessZgYKjZ5PSwIGMTxmf8RdYXMK+SR+j9oxGWuQpdUi4vSXf1/dMGi3kIYNIL
tVjkMp+holqa53nA+7tCtY3HW2DepJ/g8wOPIOV4hCxDur/AkrHHQIr5mdWgkLQc5ppoVkGjXY0D
fFxs1TS13jIcd3cW9qxwm/Uk+KH76aQyxmeWCn63uaMj/oXthFiLQyUFC/UlgjaTeA3nnK+l/kmN
Z/cMkF4Hpzx/KjPZv/bR8sr39H1vvKtdjgCjvqHZBwe42Nr5YSRsCFbXQ/73sfk2s6cYYgGqmVv9
kKqJycwKUL7uxUyelcRkYxL5ZLmL+NLhTdH9CbR9WO3wTbvZ0MRFz6v2M2uzdb/jeD2IR0MlOtLn
JmP5U9ExX0nKhI/SQxrB/mWrBtUV9NRVwMsNA9NcrfJad1OKZdnYHrwOMmVWZnUmd3g76oOIvxNh
yzF+kbLOY4NhDzlyOaqlRK5puNSlq9Pyt+4PZkXjLH8PRqcx5uYbBzag83MfMql9TX5vsStc4WP8
nuLML/LXaqSSyDHcILM2W2XA7tsDme/siDOQyUmSfhIaL3Szbu0Ch5J14skIkG7/aqmaKXgsFL8b
VWJLIwPAHj7fa9HW8/JidmAwdNC50UsEnrNKUnfXzeYEGGFU0eI0OTwC9Ru+UrZBZnZ0wDpDI44D
AeNNB72f1wuV7cqW5KdYPikpLqQbeHagDaJc6oMhCqnVBbrpj7pgA8Ir1c27ErQL1Kn6uT3LG1Z9
1StLOOcngvbozY1bNws27tcTNKGlWv+6YVdSNqiz+F7/dA/3pMsTcsT5Q+93riFmeEasxQ3ehRin
tplGJMZ+Ke9l03YJOM2NFFkGl/yth60rwjAOi4Y6Pyrgy186MC2MT7CVZEXwTmcPIikp+h+9mzNO
kMMztR0V8W67P4UIXj8Bb/yKfO5HFM/5U5QEhWPxZwzx6ZlIwHBuhqMl10fvq6JuI4Jzd2lIk2C7
IiAifUPa4TpTnE0m4/rUNGv5auKPbx01qsiky//kNKAzbfnXQUoB6SCiPMAhAqs8aa3wvattwtPG
DhF3DmNPnPA0x5I3eVxVYXckhwLw7MaZ6v4VUIKgFfyHGr8IYF5bUQjap+1AHC7W7/CUwMFvzDkB
Vv1smQYSkfijzIqI307I6nMwMQGM40Z09olTAQLa9GsnIuwYBsOzXSfIpgowU8/j1LYW1862ZNvV
eeE82ygwewEb5Xrzz7PC+44RdVOGjzzf19xIJIK5mHyHouMafbOiwrGiuUmWuxRjH0PsSSwNSM+o
USXFp1r3orT3LA8c9TCYC5jpwTFUHFacLDc9jAcQsyxcyKOGQ4rpfm6+h+wNuv1XhLdE6gV64B6X
6Nl0QUHHH6iBsx0sl+0UfmurfPUbIfsIXLEU5WbqYztOmX8LsaAG9gizjDfN52j6X+ClfkZu99ck
2P0O09INfZtcx888H1GjNHaysjB7R+bAI0sfQWDRMO4whnUlFimEWbCT01uO8bGMcQvCniSXj07L
wBJwQlphnb+HT8Nc/IxFh0IZ4WQWsxv0TgidnJQnAUHQLEctozoSVQWUysYDXCJuEQUOGjruFbtl
XuEOklwyBHd09vqbOEc4pvqD5CWeu4DKAyEXgfTjn85EBp2vTi9B8JQgmvfC1xV73pCHA2PFZBgN
RlMnksYOeLs60dqf4j5mVhZ0BIquysOjdUlVaXJ59tXqf0Yif4KULzN78t7JGlDFuzUbJkAC1cc4
jcxeUT73ZzaA+JpCIWOciHevbWuw/uvFI9jHUNsRQNG0zuJAYf3Iccu9z1ZJbjRxODLhIGBY/MqJ
bMMmbPU81KKS/mlLyZLr6qGDoVpLkHGcAuZw5LXE4fsMvmnotX4Sr02ByA2dqX1gNLKet74xTiJF
GLLo8+36a8WXTtlnO0oxG8CquD7AUjiE625514Tj3xlmVlaksz0C1yu9bvyFTczcNdy7VYw7vUud
p7arTWBDqPwwT26YF/LnA7aGFWcHSrOoX/91B9hm/VWb/QypOCN7cWjZS0yUufuJWve6wfVIDhdA
0LsCpiCDP4LncHDARqC/utkhEosVYllALv+t13WbWpmzmSki11l8s5G+8q2FUvC2//4LCyoM3fv3
d+r4UiHfJaXDpHxAK33GYv1YWkYFz2kFVmskKBxItpOZwAlUoMmGTwmvFcpzmDTxX2xM+C9Kg55t
ceVLlwXUsyxAkykjSDuc+vl+/te9M/WOhjjR8J/EYcq2IaFz/wi0qd0BQSw15hVotmnfEofE6k6+
o6Tm/wItA34kgjX1JsalY/IIC9GzPcNUVHTprJsJIU01HX4GwurZh6i0YmviV5V34Xlfri5HIrkG
HhtTMvDI6jLwDnl5bblvvU/V+kx7C3fNcS4OVueuhrlB+F/ebrHsOSXYyeKnhyl640xtRtIaBIwf
uFKH2gd2hM8P79CRee8LMZFr4JyqzTUECI2uul/8G0s/MLXJXaMQwTMN6HLO9nSnCIQNbcs0GSOj
Xj3YD3cihtSUgMpHgU0NPXjg+G1gxu12vhCp+Ba05mT7/B1o2Fa0ghfXfOvJWgNB2qhmiVTtRRai
iyOR0YSaxh5CwbgZh7zjNLuENQ1INQJ0kpwy7m2Kv98FNL35flIFJwPOdWl1UXW3TMM61lh+gSqU
f+sjQ3EEbQPVvYNm1BIdGb+utPb70HApkA/E548TrUvwTLyoBoAJDHFWWNkSjXUk/rWVaafN7fRV
l7OIGvfbXcBh9cXSvzwk2OLrMeA9kjIjuIMKrHME7bYG/oLAoM41HfCZw6QOvSc0Dyy5bu7WIciA
8Zfa/0wkrvgMfr4fylAfZvWEsnRF0gq3mBfbuUFYVqbUn3iKsNRJFPLmeT4cK6/YmC9cHrUyfJEp
XRlafwhkpnj+5PzOXt2jUnl7g5VfYBQ4i3ajwSop+Cjgvcli8fgzEx/BPI5ABdHfIeRNMWUDqGS5
4UzhJu48uzLU5+6zFKK1l955Ao7wIj5IyY1+oPGT5teRxPWCedWN+ZkxBOtzydpoNyKCBrRaU96o
Mz2o0v6nqzsJ6JnxU9nHspGNSdN1OUjZcFH7o2Sn4D0OhznZVNGUdPopaRWtwcX40XpinkH8gqjV
JLLyKzIG0mrQjrXbaBHItdvRMob9lv8HSNZTIsxJRXQ0ONYgASQFGBffAMqDWEbmk075/Y6sW9dJ
zX+sIyoHQhxFD4AGWfeWxg5sp028DhylzfZ/W+5yLgeRJ89ux+ftwHhRWR/Eij3IOnldpnXqea+j
TuPnGLzG/0mQubvaLJ6gGqJ3sNZwgphQiWjTxQ/PLkJLrz1NrZ/6BIzsKhM88BuEHVFOTdQTxfX2
TMFxF01nhhRG/0fmHi47vNw1BbvoR3qocP8Mz++LjOIRZCWDBr/m9VdKHUyMbmeunh379zzGkDpJ
WtgIFdxTvZSOhmGo0euZ1acuFGvh1eWxyvVyFXZbUvH80QgpSlwel5XNSNOVIYmiatG7yL0HiXSf
IYpX4c5ENbj/WYYfLnziyaMGFfUIST6Ix1fmmfOb1bk/VoR8Z+yDZXEt5VG5YVWJbYn9fFQuLKbm
ZOgbyNyKDuVJi8sZ8ZPD3lJIn8u58+tGZHYO+zW8+vUymVg1o4bqs/m2d3sXv/r0ZKTnyHRgtsYG
dHWALR1wdfDnoyIgOyl9GzFnvcanqw6ltyY+sjrlYGUvN9WdJL4buMD5QDdQ3LIELmYopPlS1ZIf
rH5s5lGiUWyjuFZEoZ+YD+O8Lbrc7q7p8ZM+znDDcvyqRrqKVeMT/F0NSIxHtgsmTIiDxGslbkZE
NjcBapgKZ8hNmtJm5tCBZrUpnESk0DxCh+sErToBvO77nXWSBlNCCLqYx/e3z7yYkSBFo6nxoZB1
WMPt4hPHhEBH3fDhiODH4Q2De6YYRH+uiGrdxvGz5CrOghP1H2s6GLxYuaawIDzBrt4GCtgqHteB
BdFCCNqKC4UgGqXIJMbeJfz4PPKnQXdnSa82Dxc5c85iq4mPM05Rl9VAV6TldkW8IDsxacKoCkxb
2S3ZycYylRzc/pqv/oIED7iOHhCwmmNPVct9VSBj9H4IBMKBWg4tW+w189vGljLZnNVVr9a/KdVQ
j1RhUJlpLtyX+890fGbXJjn95c4UGG09F+LZYK9gRjFur0QRuZdNpeqNgqNkHPQqJggzd/t9FdD5
/C+P59MRACJZhE8o6uRdPdng+oeOQ89AlhHVSow8kkvmqzZuxDp7VIa0Y0fOW9N3J5R9LOY2uNo9
+kkd+cBCXbbY6cjFoERnxBU+6sAW+1QMsF4QYz8ZbW7yUixELrt0AaBZ1OS6cFdbRLM7wkiwSreF
5VtVbY8szIT72vZez9gYlA2a2TMYH7BYvb3N4AQLRhb0x7cglNfENDTyFAnMwn3oMs+vTxOu12LV
uGWxRhWt0R3sTpmRY0TRFIiASRJt8VEKQPYMyhKE9M2WOLt3YoyLV/EE+vRZRMBNfqGRt+kHRPhf
zBbZRoynBfNHxbut5tBxUsAV0qnZN2BNDbb11oyntJgFPwOnUlGWAnNR4PYnTudXQp7UswLbSxDw
e52if3pgiZ5vGqMtv7ZyzUwu4Qv3rsOqYSv1w6f3StEQJNlDaiQFCJdAOY33GSSwImRdTd14+OMv
FppuqAzPjpIDFeBUBWyH9Kyu4Uszc3kuKpSwKjpgpA0ADwPD1h1xAF7NqByHwUl36OatiLarN0LX
9YCKxZ88obp1YD5B+SDOMFKmG8Du9QcDCZJwkba+IyCHujjFy602gR9n9sIp68fSH2EtnVsqZ0zE
4OYMg2kG2JKIg5xsdPU3NM9qf7ZjBMvIySzMnXTKgQjgKEr5uJ+/m61O0klBwFGhDQ0Yab69BLUT
I+r6/95sYLZHPmkvLfrDnq8V5i1qzxOmEBy2L/xGP2glcm7OCwhEHxhZplFDeWOdrUmQVa5CPhqu
iU3GCtmCRcNuBnQgM7yOZTWZUa50C7UZNeJChItyJFfv4b13StyCka6Hci4sDJVClt1m8Hga4bvR
P+udQm/bdlbg23JLuLUzTJ2YNaLs6nh8oFu/aAuux0ND4UGL0tDjA4lOrSYEKbeJkxHA3yS9COza
bgHf79x0xbKElr9vOg10aXFDljEpw0Q/YSeLaDUR24APKXVvw22HOtDtU+oH72SOs0VoNhQLYYfU
LnaHMTmXGrWpR60AhhFfXp1WtQ1Gzuv4+k2oxH0mxr5xf/VuDiP2vUE4VKQC+7gojwT6kocxjAeg
Dmu3gWxwuVYzfD02zZeKpD+TJK/JZkTkoVx8bucan9ZHkK3g95gOBDdR7fprBV1Z43/jLxpdbEov
r+sgXeVKdlP0UKP6nlSCf7z3/myFVmC6PbFyxAhjchlyKq7XtetAdlPv3C3nJF5nis0ZIJQ+XZVA
CTPO/iE0MsqfG5QX4tdL6yeMo1E1N1ZX5VLYASj+GJ6/n4Ch4V0EIkijvcV+p81bftjACPFU+JMy
ea82O5aUf92Q0yTZqe7nBXiapUsmlQS+PHLCMpf5yUO69HVHrwTQwUejDztOU9VQVNJ1FRDAu/z2
ywHT5DSEYFk4fdGfXKww+lBLzsJ8KdPPus2TNXk9Z4EpRjg2uDlWFbsRlOjq2iodY7sZALV74Tz1
w3LhPJDVFZwH8oOmKM98BZpeCgpA67aecHU5xVY+80mClFUb7w9TOcATVhTOmY3qgaG6UeP7yn6m
faWlZ9X7ai3/2CWunJ2Ue69lw8CUfJFPhFdOC02bPS3a3tatg+RhWNqK0XtSDlGMTPCyTGdKKYNg
dlx0CniB0aPWfXZN+prC5ShPM/LBpUayran/wWvKf5peMc/ss6xFRjwjluomxjdIFRiauv3mt+IS
3cOCQt8vA77Hr4i4HLflD04jfmShZDzmfGODx4A6tqTFQpKAzVvc40uskWNmyztoW0MvvkOaVCJ+
a6/Ws6zome5LRUoRYC7JxbXSMkwJkxeCHhU00rH4Pp9pOD9sWi2e2nhgJdXWB8qGVxV+hdx3qwAZ
BZDbIQFde19oTg592comAeFZLGKfIcCkawtCEDDSnyxPthweGTD/va3s1yHiREf9lGpS/t/2pwwz
/NBnHiLW3uJz4kuJM0gad6myxw1G5vruojj2TRYI0ZTK19rZVy36onRQlGcsmuuZA53CbggaqijG
PStgz5SDeJ/IpdmhzMdhtt92VnpfRkt04wA/SiazaeqHOTh7E+ESsO9SEA74hdzaEAPG22guXTKU
18RKnBe4pCX/52jUVIFvbZa9aSJ9+mmHBLONLkhc8ohp5Q+li5djALu3TUe7ZwpaXLzKX/PzLbqS
fbmji1X+G2qVG+KE5J5mCG6A1rAsiLsvbVmkvTs7r0kyLzdVLOP1PmX+SiQk2t5BqBc+g2hXQGCX
cpTxpAZ9uhyc2dG9czMDM2usMKw4e5qxYlRoJJPwukFReWhMQH89kEIjxKkse8yj4Sk0oJUtWHAR
/YEuMEmOagrIYSoefI+3D1er3irOJuPu2VHZgwMwkhBFvKS1z6M9vKPPNF6ACaE6D9eZ0P/GtkuY
im3MgGYLItC/EquBItKtkpfVDw9KQ3Zh2lEzzWA7pXD/6NjgKqJ+U1tI/RxfeutzPBcC2Fx9oA/9
ETmkWmRuH6YBVJZRSN8ibF4DM5Caz3t7k3LKxCQLAnsREeKTfLltZteovkeQ/A7oejGaGDj2Qykp
KXu2+Cjn5+7P1bGZOrxd8vHM5LR7DoN48/AiawvMtopKRBdjNTy3euSxbdtOf2oFEmM4VdDGL+Lu
Jffl/wxSGiGKTYkS34oOA1c+U25W1JZftl2cgOoXCd/tYuhum0RPCobdIpqHrpxQ+fu72lNYTFSQ
hs4Ypgk+HSyE/WIGUv6pHWJ9GionkPJsjmizrTu/ZUVDWB6tz6SxSCN4up120F50uhWL2wLqL61j
LRyvxAVbv4HBJh3PTN2ckXVelDOIOkUtECxtJlIRR/0eVL9S1dsLxnVbQeGc7e7GuJq5uL97ssqr
IN3maGtEfsH66vdpVRE1beyDFgFQ8kYSdwvLaTLUTsf2xU8HBYGUVU5cZ4MlPchiRG02ccal77Um
1ONRvC6AzyiXd8HdsnW1lH4eOKu69s4dyqAqgqbc0UylVHKLH51DYiV/0RBV+gDLqUiHIqMvoceT
aZMM31JekZpm0McXlMzsMFTXhwXrrhYnvkW7538fjgIqVf+Z6233h3N2aytOdbJM0pjukWIRNFqp
4Z4UeipytxriMpy9xFjRLNVU1rqB72ZO3GDruyFKlfp6QfHRX/eYraG7yyjmbeQIaTVZTW+MKjp/
EtJYPJlH4wysfLFAz4eGrMOeJVW0rketUlW07TUREnQP6EHZnUkWja5t/oaRuIpJOrkrpVxiE2A9
UyUVpaK0pyCRJtPKdzJYVFhYFjQqq7cgGLCMj8tOKqVnYjFHx88xM3h9SMIUpN2GuRGSUGOQM+A1
NKhc2Aw4RGVbkv1XpSLWaXDIL/d+X+nP85Swv++QB76HytLsNrZxSr0+B4vQlNT6iBH/b1tPpGiB
wAltumtWyntUN+/wo98A1e4pOgs5E/9CYEtOkhd9gFRQMgiNSYcL/wkh65WAIieyZVwACPfhYjE8
RqfWl9KCRj186rgOLzIq7x9O+bLaEzjvLyRdni8ln5KVEUhSXsoO+EuIOktaw6V+PMeAmar/LKwW
0l0ZHc0mpKtaTueU66ZCLMLCr6lpdkWN+QKCRfLv39R1WIDTwN0CR0uOzfjxs0sUAoWqorBmdpcU
qR1U98X56rGq3p1P2Y2o3XqiP6cTPwKHq4oLVnmfoiOEtQdmcHiey918jQqLjA3VwYrXzi7+b2QH
ij/kKXDLFDkkDkVa0OxYXIeij0TMmBsN1lYHMZuHHLUPbKp+eogfhD6H2L3SUTGicKy0iWeI6A8G
rUN7LneX5KIcQQ4uzhMMMgCRj91gMVrYlpehm9bFOGZMhEqcpcmyxDNOxv1zg/+wvfMXL6GNrfnU
XqJotTafZ4am6nAgbodxOsG5z68AeJfbQmxWk7GxxLC9761FOywsvwFdXYS2kODtpuKLsrotN+zf
SexaCxSgD+A3W/iakPblGOmELm8LBvYCZlXTuDBk7gWtFQPrvnjQig3kIy1081o6mf92M+jEQfE7
xnAUtyacewpyeOCFZGvLtpYaxJvVumJjkWVTpK/epC6hrAJvnQNH5pfl8bauh0i0KnbmFPW3fLq9
UVERV20aTuerIRciQxIB2iX1pyljxddnw7i8KZT7woU6zdb3DxKn7OqLX/GwliHuRf10MjGhFaZX
xootLFfUB6RS7VVryedk1Xy680pJkJSetHIZGe5Xb+6bLYpydMhwG0UDKJ4D+WAlZndaNwYU9BWS
XRCcA684QyiCt6YjyN8oYS06SIswTjgM5KdSq+ClaoTAvdCypuLls1Nd64fTit4hgYvqUOz4WjBt
0akUf2OJUoMl6ftuYyHNQec8jyBBFmU4Xo/AgE6j3cxYqWfHZY64ebH2lS0HlKuzObf3Nov94Nou
z9M+Z/RjB+UdV+GJ7Zdan4YndQyEvwLyztXyU0aU3iIxAdrpFaQ/jHza/ZRmdcRCvBeZibSLHiK4
WJs9GD0BHT/TlhV2Za3hElPVT2rzp+SKUW7V10uGYxNlRw7uKvVFI8WVS0G8MbPyWSaaibzSyYQ8
lc3r0jZ0z6X5oFi6dKp7pEIEK8vlMfKVsRRCn1J1whuiThV0ZGjs8tcDxwX/QbDCvqs09j1EANVj
MuUJX3DgLmrPTGZi8zKhMjceQStdbgpkG0qsrIpgoH1dKXvyYPdRZlHbP9xJ+sz1LeaBm/lVmsRP
WxD99fup0/tVbPTGui20utB0obNvSOBgKi/a+Yhbbkpj3O0i91pYnueVzQPpnieg5k47wmtrwbqh
6EVFqQv1FXZJgRfA5hpQ6XYt/60xoBamRgwPeKhbbpAVXwNZV8YL+mkNH7WuRWr3+ssDtjPFlY1T
f7IHHAGcdqH+rhd6AEkh4eYrqWwqNDdCHm0NvDd2zYrooUX7WxZUOtuZm0U+0em2mMNFiC3WpUzC
3oE1bRuMofSVBlLVTWb2BSWuQ5qiuvezv5HoIn13V8NhbtsM6lek5S+fkAN4DrFGcpfffqkMiUrz
gZXBDUQBZLRvQpZaegVxMFngwa3qdNk9lxw+Ik4K8dBOSCKpEm0aT7at+zkNibfjNLqY2rCFwzG/
kzd+a9wkbfhitY5zsXxHNcgN/q1aFtkRnk4K+5wi4D9+qbDeJ1WOJ/kAp8AQDfp2GY6TkEttmpnl
xFQTGH2u6M8sIsokpIaXvkgmjsdyfMbCm0oUFjOF0zYLrgJn3QEHaYElEyr/MRJx7Ex+3VGgbuSH
YMWS10HXUjWLrLGDqO+p3Pxg0M565ua/oGMqbfVrrSHylB1OgD/8KFhImOYHr6wuzq9x8yfozEFH
HaTFm1YlLOAtjhU1YtJutKiRVL0Q0XudUvh/qQ0NlMpxvDUt6YoJl7uHBaFV9euwQRstBk+NWFsI
AaCYvQqvezdVCpLnebElEzwcCfyIYOqXDrKfcw3mfSPdaHm1jiEbzlAo2JqO5a5NTDZIiwImjKKa
JxGkcDmm61rb1q8/g6NrPG3RI/NFhQbpCzYt5istGKlnAoMYSIwjdud/unLpVMsOkceSvtSYK6VB
Q6BTvDgNHqMAp8wGOlqknRUPVjvBZtjP1KswbK2bVNN+FzZIR2B3am3I2fX92soLMO7boC7dQVxs
sIsumpEWjRIXBZlKn6kWay2PHVca9hHehplR12LzjqR2Ha3+llHD7W4c2HaMuVGuQtkfe6jRJn3Z
Hcj4vZaZRvs/u3I20ODE7hGWx+gPQdXXMltc24iTN2LJsWW8umSZGSpTIhWeHG/p4rnrrqDqW1kY
tVp2ygbiKlVu6KPcWmCM6y6cLA6LiMdxhjtR0twTamTmDpyvYSmN1queCTUqJkfFYHtoQXPYjngg
ObhW0Djyz+T8QPbJhTJiL8bTnIW+cvwpiowVpcnBD8QjpfjAaYeRAegzNJ3P5/iqahX4OPO4hAkX
OT68zgDM20naKOAjn559wlI/TM/B5RFEzZJWZgyfU67vW/Ji8FSgsUzh5kxouCexpRevmdXG4ZtE
JxRnJoOXZyiPLXQSiNVF6MN//7XXJ+NsweYAPZT+T3ReBxkjACRHTNsgrE3MIL4rplhbAcP+jBcb
IubEC/zzIWlYvi3zcOtuNos2kvmIKi+K32Zm8PHQM5gbImt0Ut4vosMw2XfhSfBXGlZS2sIL70sX
RCTtdQEAkHwv/D7zPzEFz4NjYax9rgRpxOq9ZCeokeC5ZoqNf2+uSGcGIdWbtr8wFbEglCteYe+P
Hg5Xmp7NFQiwOpRwtbaQYG52VG4j5tXWzZ0srPzBexl6XEkrTYacGwpPBjV0TSM2zRW6Gz/s/JNm
ClJN8bYzfMSHr7dRdFavrqM25KnMHb2WhxUy4kyoU/7UZwCfQUXdFbi3AlMekbtw2zM9b+cE2xss
8AbZkV5FKqt5hKCMIbQu4vKMpBdbNxHDWLhqCFfNuV4g0a/n22Kk/hDOLEh2rHGO6CumVpgQWSg2
f49Sw53MDhms23HIIxq6IB9p6D6RP6eyj04UgaMvH/8IdX2SQEhoyhdokuLA0dPlkbyXkoxoFVdV
5z0rwmmssNkjuFs03LCYx8OIEutOWXKb1fKrKiUQbZzV81wo8a+F1tG38g+zxtNi7x6Yp8ogFgIl
X95/A1bF3sT+kbwqwsHkYX2/E85PzwxSP+nJQLDbqGRH8r9HdyhcuNraEE+XxxgwaYtnbS9JjkpR
qDyG7RktHdD57AkjfPAIDoyJHgfidDz6nG8RR+IamYAves6dqYSTvRle8d/j+yAS9C7lVw8dp4W4
booJxkjdnCe6cQM38+GVGubzMF7y2CUF/+PddH653KiP/IllxY6oZmQvUiHaz+8Q92hgRdZ/1tkg
DsyR4W9iDnB94QkhQUaoYI8SdpQHWWEE46bgBb2XRGzNI9M27ubYx5H3Nhpiy7cKuvuTLt6vII+Y
1wh+RSnhWLZZ0ejpmKRyTSYWbbgNdoYwri0LD+n8s+6qHN0cSGJKbEUpl2yN8uPAETPmg5BqBVfg
J+EvdOWq7AAQc2Vq11gXrs+7gxVy3GlZi1yPlmczzzhAJ4AlBl89f4h9Evtu8gBALRh6RLluULDT
V2mmEGW3rQq9Y5qem7mreumVj2xj0t0prjoLlwDYzkhKy/LAPlgEZIHhccTgC84ThdtL3d+7Q9bL
GgQmMbX9lDEhg6BGz7nFLU4ZVEQmOFxoFvymakArY3X34y66efIWR/sY9Oga/AAxfIy2wFg2r4hX
KwFnSl2gO85c4BkZHwA2n2gX/Is+1TBX2RdAAX3rtrUJDp5jiPPfPJGgTZzXFNWm2SaQHzhkq0fv
CjoVCeF8Of9qjaChAejp6elL9HEzXdubh/5Myv1pkSetPBw0WKu0/J0q+9Edm4LbGihbVXsiqPQD
txZ5+X3vXqYxkSsI7cEgStKbpF6+2kcNHOQQ+fsY4/L0grWpvZ28juxC5SaqaB/m3WEBUVdSpdyc
Z+Tr8oNS9LXNfm943HsCC5Oi0nMozWSfiXWPIIorLexu1ArRyGSTsBnLNkn8X/gUjnLaePr7qgRg
fC4wmRnfxe5nIHTs3popAujEQtZvKM5l65mhBsKsD4FNBQJOA6ojTk0KZe7zzGWYFuNf3etvFBgK
rKpFC/pnO+qIghPc5Pk5Wo6b47phvXqrLVbC33iUOCsuqPvzURchdmMh6g8r71yE4jLjn5emJyLT
h92T8aknHmldpm+eAa+fOZALWRBqbM9upEGgNkGV1XVKol1jcfNn8AElzfHoS83nNkaRnzkG4Xu0
SCeDFy+Foq04+K8OcJc0Ws1L0KJCB66ePPNPu+tVG+E4jzIHApHNolSzG8JNrmynGiUlGKFNGnZY
imqCFgSV5omxCC8fSILFR7wveolQMEEShezvELSPcTb7X6EcEP60TZ7kMrlNeXA7pWg/6j5xtrX1
Ie8dTZ/XSAzdAbFv4WS7kEOC8+u3Axr99C/u6j7N40PLRPAcDwj7bDDcxjdwxQsMJMq9sP6OUug1
TZZSJwgatqO9HLEJ8XWYi4cASUjW82TgQcwhOd3DNYNHJ0OgGWx2rM49sHE9836Yd3TqWy58n1fJ
2BfI1rSGLHGtvZhj6PlM+cZKR0z8y2Q9gZgYvmH+ExljvjgD/Ux+JQTzY54UzoCQf4uCruC/ElnK
JECJG3RNDyXRY8dnyodx3qYgU+M+nQ5xWwqg9jX4M5/bMaJz2FYK4YlHkUtw5eMCzBcbE8TJUo1K
qbER1Svzt4pQKIGZe+7RvHStruH4f2F2hTzfRjFJVvfjypqZN2jbJhRP0+mGDMQXkcx8kkQIkUez
ELMTu7ltB2kmq19LK9rw/TmyiE/jIB1yxkm4ioYpI3l2ryy896Ix7JuQ/brQ88AQc0szTCpCuzau
juH5L+I1jcp/XidMa8HqH0lX0bH9sKAaEj3519bUkyiGnP2xZkt5ImyB5uJvEPXr6r+BrwMFWETE
fnvrOmiuMcmzh/ZVwuYDr5pGR8wlKpQNMLLMkqHEiF3bfMxKqE/+hIN9m7WT/S8BJDM3ZEXII/pD
H+r9H+3HRHeWItoi/+/YJs2icmSG3dozVk5TMw6F54PI16ptsG8YcQgmh/Zyr1F2wAU42tyU7GLl
FCc3Zsl8MQuCCb91kHp3OTyTP/cjOMY0kiIsD9nC+lh0nAkdYhc75AN7EODI6CSER1Dmo8Bl1OA4
e+yfJXprf1GXnLo99U0N8Qaf237m0x04ZaW8Xc5UxAKPYhJT9xe983Q34DAl0hFEDdFLG8c6rBey
ZuSUZ4B9/D2gJMhBMQncvRWEXBmGSxT9lD7Y2MYCx2DW/AvWhDi4kaw8sHYvmX+G6MhzHMdgVoxy
YLGRdG5mkO0YbQLQQcA4oo+mZrwObCdsXGWG+IvAXBHHfNX7Xsw+VM75MUgqeXfcJruCQRFGwut7
Gnil9dSY3/flSPlmjJbRJ/K3ZvJ1FFrPywnPrN1gY1SSBpp+E5w3yt9Vurutf4VmNONTk6AFuarB
ZWAtmbjM68F9fPhIejHjv7Ok4ihUFD5kBCdV8vGd5D+ib3EBcy87eulT9Qk7loTBWy+hdeQ/8eaq
hTvMX75OtgVbptMzrUdFK2KZ4LJtzZ9K0oUD+isqMh5HCjgxMgSfs0eAfvaHEO4fiH8hnaofhNii
JJdpTShh9DgA8NzmCGC1tCv5AJtmL+HhTxSuTFIPNVpeMAVcuvtd4ncQozU74BRKmXUY8h6paFbg
9ysh8XHOX8iMrXznYI8MpqFMgEZ70Vn7XKiLXSnCb9omtFXpdwBr4Mx7RPt1aVDyhJOsCcphfRid
M8If6TYKhYScFuRRtk/mJnd5yvbj0rln699J/duDyF0lUxuhbGZPndiIKX4hZZco0K/JJZnZAiwA
JyBatlo1zF83NEoQpZt7SDggJ9OyAAnSnDAWO2JqMEmjJ5fD/XDeinDfLuxEeGLOL4vzQVYNVvk0
1CP6vJtSmbaP99s0tZxYTM8RA+HyusS3xkXns/PJNSM6uR9VnDZPpcqM+JpUr4mTM1S6MYx398yv
59BItaTrTsn2Ab+2LzZKSvpuXVAy5rXd7e2V7d2IE2C+eU/K2vVuxOGHzVgxGHPzbltNPiDen1py
KOW9EbbCE/eu2sWtVS+l1LojF1JHNXCtKVLG6MqIejfKmRNKPM8bcvvwlMPa13oBBGaPIPevUXPy
zIEOsl2VqphmyBBxAEqk5z4h4qBoyrhICAKa9rhsDt60wEVgJNK0H2huDJvZUqEjem2ieXZx3gz5
gcjuNePIf9l4vV2mMyQwnI07P7StK6s7S4mL6N+rFBI+jf/zuTXvCHiJ0d711+n5+zf0m8yMS26N
03RJpKKy4inaIMmORp3WdEWdwrGKheARmUo2nojD7m6T8DpXcQn8KLYiiiRPs+H2GKAz95BLIf01
kCTWwFBZj0fIWbjnEqClOOQhUvZmFzVew6wChIo/nsacM8RRdo4S/19PQj4Ktf5b0rQFuPk8mc7H
88NHpj3/s9knQK8BymbcccByRaRUt4F2tZZ4IrWPfD9MxEGHQUCVSUQkPIiMFw8tiEVKhaVxgJLH
IyoHpOGfkzqWTZYHSXWCxKlfm5yb80QaMthPe25xy5IORtlGfu0yCwHtGiDpo+dGzRDDPA6MNQVv
MP7h/kIvOdlHbrg7KXvo/P5M3khzExcukWLYZRdlwRGPQT2OIGWLBVMBJTxuxwkm364guesdPO61
HIgvVJz3uXPLAzPpXP+/U/H3dr8bijiNTI5HgvmHz8Wp3FvBk5J6e71fx2hTBqkdh/VNM18TqKqy
QaO2wUn7eV1g2THt5mj+VJt12Wmm96/R4jY80+i9GA7qfQ+rgyJAvC9oi2WD0F3uflyKoIxXiSXV
AGVFsqy1HODhOgmf6FH1kGRa1es3b6mzDhjJ1r2ys+Icpq6ZkNnWDduIOrfuQDt3PXBW+2alSsut
oY78m/h4ojHDgbnUHMvAeh+JeYr/ZX4OqOdv7LgYtUF2K12oSwXR7UuygFhoeWqQYigvNaU7sW2b
3p93EUWzT/jkSRXhTHlv7WsaCZb5FNCBUlF2cSzEX4AUesG5YmU4NyLaF4ih6o8Z01sNwTwjmWC/
/IyW3RCaL5Dooa4/nP1cQVyswlV/HZTeGaJ1WpwWm0MCMP0piybgldFUTlyGgSD87gY8OjU5+T35
ddCxZYTUJ++Ye5q+ypeY4OoNWnWEvmksNb6it0sErBUXwg1BwD7FjEoDfxQuD6XkwFXfv6AprZ1H
e32EF9IOqEH4vqeS0Mkog1Y47iHSkAebNQUWGPqdc7PyVzSOBBIFZb5eSEXGLU9rDn6P0ca7Qp7z
335rn26agIAB7m0dqr/eVQMpAAuwVWGzGSkHP17EXIu/CFEjKIXQ8e92EEQstgVP2mY8uwXQDf9E
Hv/9oHjXg/BrTUnA5yqLv0zB1gfBumM6WcRo9UFO211pcE98Zt6uLkPHZi86u7tGk3M0lXbja/us
OKGbuWuAAHBE07TrrsheUIN9S4kljTsCdksohZnNa20FP0kiDHXgU269t4cSA4oGi+AuqH0tT75a
pu94Q3UpVI9lScKCq0EBIU4Sbsh7FezGwSvJ+F1pnYKIFz3SWR4ithRu3ULMdGZIOvuxdxsor0zJ
9Ur4Hx3H65TyujoXpiNdrNCxvw7+ggF9TJy72AcrYBrclER7WJ/7Unvcw7WBsAEXcANe8R44kd7d
IexuJ21U6Dbe881cf74EkELk3mazsUazswpqDg2FXYqfFjAc6WrW+aVg5VvGqyoTo0nBadX4gkQI
HaWZYfnp+GngncyIR9CoXf4N4nXgfV4ZG6VX120aYtTsxLU0py9cg9rdsIprHSkRNeR8kA1zH6LR
7lef0EnusK+FxDg2bialMOAwgxJC3nOYf/acqQS9AwH41TmYVxBHmGog6s7nk1iRHm2p8NesuP2Z
61mQf+7CrmJmxwFyQm51LM2p7LPfIBxcDap3lm7K7Co32Bt9qCryiWUl15o5DedjDpAjGiHWhvwI
0BQv6TMOHNedLZ//vB2saDFHQhx3juUwWTi33fbfOmeJMQ8qmc9E9s8BhpVUmY0BeVV8NZcxmSEl
rmp/rJgLK2Ex09viROo5IvFfNdJ06y47owIB31r7cJjZ5CgYoNY93aJ5KN5ztnIkeoRfp06cHaPa
wGDEJ+ZOhGoWC/zDnPvyyHDs7a1o8522pSW05HoW4w6dydMyQJq0tCPepnqQVxde6OZ9EE48qtpy
an+d2Jl97Q7inC3YZBH+XEYNWhZBCFjl0Oxs5X9iiOyreTAogKQDz5mdVpZ5+sWqirOQUneC90X/
tGzgUfsITZs/XreTWQ/om+d7eUu3WIZLlLlb/BWpuJ+7rARAlFFHD0q6hn84tT4M0ujVW85GF2D0
pb/NANiCMzTg1mml2lPeYMsVtH2d8ONLWg0MC3eSdqy3SR28nzV6q29uFz7+TnGbhdBodg/fIWRU
f7bpXcxeA8UwMtjaAvkO2vbArA4QjtNF5zkoRmANheDHMy3p3p6gq+R+5BAM3AT65W2+jXSL9/6N
bVa3JMIQfsL6Zwp5g21tPXaIlyX9DUeAR7uukv/3ZZDjo8kDHWm6DKFnO9hwEDhiICPwC5vGFBJ9
oF+3cGJWYVbny8/BOcsoXwUKo/gyWV+FkTy4lAK6hHurhaAgMZXVBTBkGWfUT7XlJn5evxruq1hu
+VTPGBq/mPnTajRz+DCCcbjrYDupgD1BhmgSjZm+TvGQ30QyfR/VRPtWZ8SDf8ivC74iJEDxgPyz
3RYcEpTWH9GmE039XsJXeelDvDKSWKFeZLIbEKlUE2Ur30olF/9Y53bgeLXjHWR4NDuZHJDi0fJF
CNzfNYADqLLqTmqkh/YgGImN9Aku6dRxsjiC/r7rBeLACLZ4SjnHTmMf7d6Lt+SqJoTzUAMfucGy
GOQKuLiTm0Rg307jcCcn8OglNFerWd8mF5E2jKh8OcKsP7jiwDcezX0omzlIzjeFyeyfEtALpGZ5
6ON6HY4+Xii0tS6wy+WhGL5OPEHls+cWzwav8R8mM6C+BRNHDBgzqxu3vpquOx9WqB+c/lxaqv68
fgZmWm6sf2nfP/tYufIBkq0au4z/JvUa+SHahMvCyJw/znUeOD+4RlT9nk6A+4wj/ffypQdwD5Ul
NB00t6p07mEkAFMbov7JiLyPjkCQu9JQhg+m0J8p35M0PMjGXo3GzB3jI8Ig8MX5bgZTyffSYNO1
nuljnrO5C3wWRXtDEArKSCk1L2dJD16k4yTsTmHwu+LOiA9H2M+60gbMTUKulCh/B99d/S9PJb5H
ZE+93hFF3yRLRd5gN2iVvTHLr0tSnfHrBWVZ53/n8WF203Hb4/nxPpFBiuZR7rd1oIYCS3TksAPC
aQ6/cTL3WiVeL7DGnZwEjkugamIW/MlTQCkgTUBcyu3xoyk94N2WxoSq1BCK+F2OSJvajQ8C44VE
fG//Mc4O1NfUnnTQX/Qj0Kk6svlAdu47/Xyboi6kt8qZrJ94gY222LspSABGEkVseNkN73L9lnKw
zfU5/wPjEnS32fJicq2bm5hBdfa4Wh1si/RdcbW6xb3FR+yAqjqo7J4LwqPbSP0DFTGM2VVJhv3Q
7iRiKY9TnisYJXo7K/d44I3j5i2GO+wqFpXkroIFp1dxJ8sxOmy21qUiou1mrzmnJrqMmimW7nug
sdFrA/jlQjjydB48hqI5zpomSYno+dycNP3ew3MlDI4pw0B6+NQrShPPlhYQnt76vt7Fl/43GP7z
owfaQ5Lm5EcpIUC4FPYTmE2CpXRiMa1RryLPRvbnxjbR/JOW5NHlAuFDanlZHdr3wX2Q5OGD0PAg
HJiLvecdJ+/cVSsAZL3Yi2egy1FxUCa0kVOVeZ6dmsQSpztm+7FurVZNGIQfZIA8cOm9xLYSZpRP
gGBXqgBRh1Q56a+mnzCTw+QYpIbS7fjqOR7rLbErib6pCwXTgFV/7HFOCdaHOcAjirGflp4PMfea
VTkAiLNAYvCSOgWDCPnJGUsErF0+Q38T2icWQHpqhnKEUslIu8OzH4zexbBgO6Rwf8RCmGRw2Z+J
DbGGnIuLvC1tgirX0N5m3sPOxNt+FcZkBkfHCSPbH9NLxxoD8VXcM9AEC8EOMwzSAk1jWeJkw/qG
tjbqT5pfbuj464hhcKsTpS2RlkAmoqvmVmwb0XZ6/Fpv5ew+9WeQSi9lDcw0bjZB5yT2ujrcG+DN
8qmCa5ZV9Ci0Q6SPp4G9AZNb/zC3VsdRflxuAkiA+ZUtj7qQPABuE66Mgecq24I4krrcBNtyBale
ByISB07dCl9S4N/hl3jYZxbD6kV+9ijn96UiDJK0wJtwsNsXt325W+imsFRaQhHHS2SqMoNJg/S8
AfwHBm8dpayIHujqOnwYO6z4t9bfKFOU37iZ26pfOEQ7OJwkhf2N6KKqdQ7+3jWLG+ELtSxtx4m1
qSkMQSVLdnW5JTOVevCCOKSf57CnFfn9a0G5O6B5DUFf9RRlelGpG6cXtt55W0TFCiK6ru+fsZxx
/NgFw6PfjySPDdRFPIK+rjp18EApR71a6RBJa6ErOHEvnfIYpWoO02M+thN4cS9CinaoBlPXwPzP
MAAnAI8TuQ/CZ/aMfC0s80Crae/chbG/ILQkrpJDrxA71s3Lpwzf74ctYs45mGwJF7KNgDLvjbFQ
SzCKvTS4A/StMVzY8InDugXWuMPQMJKvjgv7IyktUVzanxmu28stJGMEnruY/P+qkFWw3y9AskFU
Ob9U3hnrxRC0kMjijlRmZN9IYx7g1Zh4//9/CBAL2TxKCSLYh1Bfjx4APcnumoUZ733wlgwyG2cJ
YdhK4ScVz/n2tEYhbmFOy0XzU0Ntb2n2bQvfFokwFPgWAENI/8OgzefBK8cAV93UuuTXgFHmlnJQ
wKZwwNNgQXhI7hU8Z7jOKO1Vol0kro9ZtQm1UMfuCx90s982mV8AF3p1kHHGu5ldRq6/1JMN5yAQ
+AlpmITHLpn4LKJiH5mccmv+21iamp6641m9jef4+IUFG7V2YGB56gyb+MiXcPuujDI5fvPdFrRQ
ncEwIsNPnlR2/C2l0lwLoSxRsOsCRXryiv5z6EYjjJS9j4YZtk1rlkolr9RMOZbuceBaLmwwJcuX
r/JyoCY8m+Z0UaOp0J36oYt7q3vacPqpxbCRPSSAeI7oNzXEB7UZOQ4h+gLJ96k4uX2jJbvI5RI/
xPJo+roQXfnmIPSZEIUIZqdnMTuHcMBsGX+7UFuzAWyVo2UCHdLmphqoEeG/Wiz3NoM/3nuQ6JnO
kQagn8ITCFKh3FJQLgGLxlCp3EJsWcBtNelXFFlaLmFKbZaLHizhYNVUAP48TfuuJk+tyxZ+0hlI
6rmwWpTm9cVhRezd39whLzHOuBPx/Ay74dRepu3t8nTXhf7Y9GWuJjnZ5nUdtYoyOlQsPmf70gAe
CEnx3c2j+FeGKdBlJhaL0mGzPKrx4mLBkjIO5BIdv/pggHUL13H5rWKNSxvMLDMGRVjRrgclUm3X
rSieenUXcmZ3m0WMaJs5AEub8X77APDa/ctDeIy2F3NUZ1vL4vkldEhqFk6f/LdKHEsPd88gKn5t
YApfR3L5Iz1ZleR7iJp8IC01lFaxDHGt+2VOvGtzKw1TuzIwdpQGubdFw0tEFihL8Oyns14CPYVV
zAX23UL7RQZPgz1aBTqoYO2vs6apcTel+r3AsTXoLQAFujvtZYqVrbMPtFn+YOoynrZlgI6YSoMo
x34y6UkvaTsAXs3Ub3mkqZkI4KfR5zA23Pw3z0VzXKUBEyvY403E66X9U24IeAhzck1hbLNPbDD7
QP0gFhWGCDxeSs/Hr95gJ4Fh5tInzLLAdBet55fryrTmvrB6lDgoqkJ7wL6Igaa4tNsARoTkitEE
6m9hf+f9QBEIVWv0PSbztATyylbkP44Serh8IfKfIGxhB1Lt1xdowvt0YnZmkFr+HT13v0x5qFCd
Kse81cudnrOo19oVEQuoajbSO55XIZU10dIkJvJqn7rI6xjSg2ggHp2DFVJh7k9tLcq5k3JEDVJN
AuSzLb8ORZbp4Cmyvr+oy8mZMAIgmB/KtzzdJTi/Sryb7xGzUjKFKczLczwfETX+lA4dHp3WAzrJ
L2Z19It0f7S1XgziSIGKwQgCxTKGRVAaS+Mv+l6Tno148eudKk68rlWLeOnIxa9tCUXhE72ZJP6M
qF2cAuUgCzI2weU/E7j7cr+AApSJLi3yb5FnOwLm5jVuQHfUqCFMuOO3P3KMrg52dJyXyZyHSHe6
beL2Lsxvvu2ZRbcvxulPHUhvw7VNkG18NPdWFzk3+c/f3NY7uS2f4bLUQpV6CQLm37hxJWo8mSDr
AkQICZbRlUmYj4LzN2HxAk1yWvwKTLugDfETDTTo/ZoprcXYl7JVa8d94rNfrBTJzn1Zkt6D3UvH
Vqkni1DjmUu54gnX9iEC2p8/Phie33K3HFtVuz8nHtL8C9YTHSzOScepWr6cJK3UU0/DEdnOfkq2
Df/FtomKkrUyFyavmdBHY0KlycyJHqMlCH6F/DaeiqNM4sDE2vSOH6EDODi1E49o/JNSR34Qnh6q
lACL3uKOsCeed1h5URvGq/he6ot54JvAVO8v88JEVHVIeKFEANj7aUpy/A3FftFh0TR6Enf6uini
SSX/lJNHEEP9xT9E+ixgQroR8BFYpTa5FuuZdESHJP9CfRLkiOo9RrWzS9n2LjWbU1aBLMCi8gkg
UpsgZACR3FI6/jfrqVzWcm6I/ZwafeQGSUMCGNQE5js1cvdTDNQYL9bQ0WFXhg60oK1QB/e9KDAY
cNiAiOtojeUlK/blljBoWS+dOgqsqsOm/elRAgH8iUKQJX/qv2FW/pgsuQVPcqjTYkU5MBvf2Zde
A3bEONZOwBSbEPNP3y2K9zxnlZKl9+3Xxow0EQcBBtLxFoxmrx9lZuD1J1HHF5fOsBFDwnWdIjUP
C07CcSlU78WjaxorTtiHO/EMtQJJ5nC1vH0k/HDRfvbMb2Kolm1IE0g4Vm9BQvvE5+MnpLYPokoL
/qNYhwNNZEeJ9Yj+Cg5i8HaUKB/6njSrO1HAyCvoAnxO99OyRXfDJpHR/GDkPUfOSw/I1+g6CX2t
jragWSRQUxvPM6xvG9qq37DuCpyEe//oKpGFx2MNyThspmDDyM8OiUXbKpZAasi/2IEilmDZnNWn
lHbwVONF/VcuvUTgxOdhLasdrikzg1ahhkcGKhY0m7Dd7YbvhmcoCiSK87hktx69TNIvrJtNQn5F
HiL4PpL6KoEVfVuDGI0XjsHq1QZrAl1pU8o7tYI8dmbaq6zaLPsABUikHcGwBRLUfQVR8FHrQOeX
93rU7+Aix/z+D3FBr8XtraeqhNPehIR5imfTSYedQ7l4136YzXaEgABvL5/7nVngiNvL11oklnyG
udw+kD2NG1BuCs33klphZUKZ7HIEY5aQw73e8aGEZg9SpyzA5AbJKxPJzKMrBewPw9TqflXY396s
dB3TboSnYd4r/GZm8JWDvF0SSzZNl+EAfOz6ene168x8arqCNwdNvHuSw/HwykY9RsYI9aFyEOZ3
wWXdRzHxEC/MfH434v2MMkvtpCAP3fR6vhWKLFs0h6i/pDJQRTjjErcTH3jGYB/LpjLx9WXa52DT
c4Mre+PkrYgP/KOCYqJ8fcjETgM338+o9rpwVwG+tS0hD+M1dbDyxrMhAZ4ep9zWLuTPDBVHj4We
UZA3LlW4kWkFj6p1e9mILKd2FjG4MvzLF+G36ww2521yVZzCAK6+yamm3bGYHdoMvWjnWjMwL5xp
2zn2ityK+HCt7qPSQC43sZe9WNW8PakuBrFohJmfJJ1c9l0WG+2YICKAfqjnPJdjWl5WO+/RoqxL
dh1+1NzPgM4iMwt8xGpgQsfpaDpnAT7ltmKiC1kcOxGBj8zuGaaez0yk6V9aKqtQW7VoLpkrf38L
l26IwPAcOvyyVvQNPQ6vy8HlCBX0zp/TZVR8f0uiZCr69Y1i1pLEf+WEN8avdvvzpp/XGp8vK88G
vMB9fGrAAvLzS/Vt8cu0nQatOBPzTyh3dd5nPZ5jN1YI00ZHFlUr1ZQJ5H9MN54pPCjezvRF5Wlt
wd57vpX19ve2adVCq/k+i2az6l8lio9+HI0c1VK3NfrQjaF1EK+JiSLjaECLPRIPQOhR0pStA/5U
TuCNLHBAtALvW6Blt8MUAXDPJjF2uKuvOlfB5lv+gf1htrNmnU8s9vSRF7qJOBstZ2E1EHtvBjAe
3wuI7qxDymor5Mtwv1w97NMy6HQUv1UwHzuL0jZr/0d3KgYFI7NEIsSbb0JHPKzYQlnoHJauCg6J
I4JYxtrAvhOAgzxOKk1TSCt3k80N7zEXGVeOIR0uRgD8zmC76UKSfnhqMkK5/PdJ2nEBxlt4ddhT
Pp//exJbkBnG8kLZTHxm46rfPhDmPN2TjhUxipRfTYDsbEvfiULWy0+nJb3nmXaPDs1TCfLkSiCY
K11ym9TsHIJ4oJgXfvhAi3U92jdxdZnrdYm13sUMqFIPWezGOWrpySt1MDXX3xZ6KFPW+sJViwLi
Zso1aBk1qdkKR8kTWds+TH9rrob1bOWBjZNpv8yXSYyU0B2kXoX7K2XrSVQsj9cGoO4eAi87VPXy
6PkXD5OPhc6APAP6Sy89wO5abl3RY4bO9PCajgZ/uZLKuSxbVjdZzwDIsiNdiIEKl+rwbS9Mp/7n
krRVJ0uVqG/0byxXBHHJkb31gIu9+LLWghLQlgLWbgEbZK0zut2SE82e8sCCjivLmiveJjMa3+Nm
CQXE+M0RHMNujD0hLO92Kr54czHlV7qiJ4YKNbApy5+oI9NPA5je4Hy2zA7rXea5Mm7uQiJ1zN+5
aUa2yPv1DYFWGq+MA2XseraH5emp8arc2tC7orLeFwAo7bONlPbN0fX/9jNlHM3DyqboAS100/wc
xxXc+egiXBJs9koeTyp1SZwwpKiaKLtQ7jPqphDR3cZ4+VK1WygNEFIVkEZRLMbAnM4bnnu+8odo
ddD92flJbuWcJ4WRtwq9dLnHTFtpiqFThQtJUKDTHUhPvE08YUUDIQvWP8pSPQO1L4SJUfBUbfr7
1NqawLjR7ORPt5eTvoYrgcves+n/9OVwqRXkaN5yLUegsrwSiJV6J2cDs29lXIH98R+MQvGl284P
w0SdHDniqLLgT95IHBUJot5C4Mro9Hq36kGdFa4MWMcfg9iJ9fstYyGJAP53FcGl8g76VlW7zOkY
Ksxt6RIulMVBDknSNHRbeRdJnqQGcWEWYk1x4r0529VnRA3a8NrQdY1rpFL5YlfZJVImDKKdMQ9C
j+lw0WwrBsfTpF3Y6eewcI37d7LSc47NmbPcMjL09R9cf3sutGyx8TtDFwKfS1x1JwMvM0XSvdT9
NoDSfMDMxvhiY0N3k8T5UrPxZ2LQSs+hUxCg1XQoug152Yb5QrCl3Cr7ManalGXMaX3RcKRTJnI8
pgzyKrl3eLdUOhG7lPrY4fRGniJSSCDnkX1LkUu3fMu+I9atl2ehdA8L+qTqepyMqjWIdlgY8f7b
x4QJwmc+cexG8g0bGWLRDPtBR0PBOf3x8NRpNIMyI8GsOhUydF0hZ0GKmaioHi8kDnIdWSe614na
tmkQdR8rNFBGgsMNLDHeQDhD0ADlkB6YDhd0nrY7gkINQmMzqpqKbtx4mZW/rzRjSDphV/+6Kdix
YGGj0NEc/Flvs7xjnfMJ3nkCPO5XI2V6t1th0G7nTexrBTIsSL07iAh/BMhbX01bGn/ncy4+/BWq
+RYXVIbhefesBoYWFnTsel/uwfBFznXM08OIUiKNt9Sjg79XQXrjh+yTa7rb8BI9nb+7b1mdT6oQ
m3RlhG0BGyQ25TSvZPZql8Ctxs2U3sLcEO0hpSUAVWkg4taGMfASAn/mcWLGARmlpoWUK5x5PO9D
GpX1QF9Mr8H1W6OGfkSOoMK0BQLZbzbmXW8oh2dtsSuQ7xiW1gPvXJEx7L438N3rM1LeStmlp6aP
LQinOlHlq2H4pzrMq12/+Wns1BHuGH9egQ1uAYJpSXUtfx28CDDnmTUuECeAh8yBBnXTYWMy12df
/E1tHZGi28ogWHGSbNAGfd6IS+0vpRoeNTazYqE6WiNHgMk3rFM5NzbTSjg659ngU+WrUaSVQlYr
5hZQCTPmuV515s2kQnc+cEoMM204yMf5i9qgnnCQofzsz9L1jkg3JqJauIbKv4ro87yx+TN636NT
FE762ul24POwndpvAY0IggCTzQuxaTtZpdqc1lt0tTOY7bwTSZAoooynm7A9lRtWDHc1AZG5OCHn
Du9ooNO9TmTtp2axIGuF2SwsgtxFaIo6DlQ0qcBDrpuq5wRIeigmk1uYlT/Vq1JuxZg8SRZYIcZJ
LuQElkr9OnpHx5h5sL1oYM/pVwKP9Wb8H2wKu66U/Uy3+3S6oqK4IEUuKbSZkChM2moO4Y64Tc2f
X23sbSZENNpgpxABAj9gu5iI3ZqUA1mwGC2weadbgKHX3pKUOIFKvC3DQ0FUoUHl8ItjasePW2ib
Gjv7o+MA1mkIdjrWoVJafbdIx8drs/LujZp19hFjSCelEXVrarbwZNS0h4mS5yBPNOJsTQNcEQDo
USfO6J1/NcYw4dpld7rNYz1XngLU+LG5t+6MjvKldCzF6WufMzlsPcnN844zEA9pVqx1IwZ5FvtQ
2L+q9qUjVB4700iiEtqJJJhmkBItGNCP7dc5KSPTbFPQCSpkfDyPCzamXEsFzwltcfsySpbqe42+
PN7DGtqcN0mUswF9gAee3T1yfse2FRf3mR5xTE8JeUNWfpYiXpXXZFDAz/O3vW0YbvMd129fV2qm
nMji9CwHQ8GdBpN1QACr2HX0L5lLT8rAzMN/Z5DHO9oe8G9shJc7f2gdGsMcvpVTAXyraYn/5YqT
+j8HNeOaeq3cZDyu8tMY0Tj/q5Sq01C3PfOblHnwGgy6DHSTBE190/KrHGRH8ac9WS5RjokoG/a9
k+03egDWS2JDGlYD8JJM1hLViswJVjWNog8pae/JtyQV1Sa1N+H/oB/pW+XrUP2fY0IwCs32iJzU
0R0DZdtNNlCKWxfHZJ2FCuqpcuLZASb5f8ZDVTi3T0CHbt21Vd+z3MSU9QZkmOl0Ly5A6PkotSUE
RF0BwpgXVN8LbrwK5IEwyDBre610a1J3q1t8irVr5OnC+GPh+YoMt+NGNw5WA0q6Bkz5dQekZtXt
EYmh6R/hjl2YRbEAe743tYqRAdMOyVGSLHDuuC32p0+p9CJJf5AhlT3qofqGjmstlKN5zqjRy+jV
8DifknoCqLd1NdZBs3kmJxztZ23832BntTfQhE7rZaKBugzMkR0JMw79KjUgOMJkCGfP4ErHlKK+
8jJziIL8cFyJzhDw1zdEo4YO/hx2lEO/5Hw0ZTreK+ne8bQFjkHb9elzQCpWJWmtgoYtccXCj1BP
em4/2uaxW2IK59l7XiI4omBhF+qMBlDhcfcl0soJxdt0XhEseqRlsjHMnNJgZeKHOBKOUGJuUbj5
K1TCUMCDfwFhTYowbFy3+qwcG0rxvRNDmgaBHG1g9iJqgQzWrJ4ML/+5bWkcEaNYfdcgWhLTg2RQ
n3NWjx0/PkSbVBuW5ii//Wy/QO86FxUfmZhKYu9wmm5lY2JNbCuvIqg1pyO5jT2UZG63ruC9UweI
Kh5bpAi4usJtGFdw0j8YYgBKxoKg3AhlUZaoaF/I0PCmGjJi2m+LONK16o6Yzrqf400CAN+5Ol0r
nuzjTsBjqVzAaOrlRtX23vbw4uiIq+/LoVPIu5TIVYYZ30MvcOvVCggvvGAs72cpjRCBngu99EV5
mX4EZKNJpdQJtucqhPCraZV6xgEbzXb66S2aAij/j6hSUvTpuk/OvmB3rEBJftOumk3XUcVI+7Uz
YufKN1GD9RRyvrkGDwYenQEtNDSo3UGcnzp9tkrID5wT6qQuymbBFIcljtZan3eNrZj5v08dNyAo
gyepxyn7ipbe22RHp8oknm2ZbYOFhrv9miSO8BJyuftjO4IHLcnSjXPf7XKAylPYftJ+bC786E9e
PEvMRKF3u7d1CDKxl/9/Vuw4jCGnyKydLuuj5LCja2zqqXnQkKH33/6KC8W+Xrf2TTEXubiC1bxr
Ltu7e8+xmGq94DKKFYLYyng5ac97RLjQM0OF2YgXsLwbPqrUy/k/qcxFslg9r91ju6zMeAWUJIPe
pv3Dmm17+niiEqFdknwJeGgRFaEyWRrKg+mp9XAn00Pcs18OJ9zOtWxuOptnYX9mQr73IP56d/I3
gXRqbtbg12LUy2AaCYTUdUfxIDUZGnJW0qGQx+4bh2ZCHetNsSiALbTRWyye5mC1+iutI94sFiZl
FLTG+FzyQ87k2l3JAX85pIfhNnZuO/wojWlPl7MyBKxQtrTeVNcZtdFd2CeacRPMZHApC8Tumi3c
Q24lNmJaZRnhNrZTX7tf4qfL8nEOce3zVRnum/aXqGJVyoqmOdy0dnuafORFGli9w+7+hIwnqNnZ
wnlEvEE4hAv36Haf8inhU6lIgmoSp91mTfQ5i68p2GNS3PTNk0ltj3SAHadWVvO2y0xxbd+kvPxn
1lryDDg7DccP3OZzsJqpfPARMcLQGiU10Lcli037Aj5Z8t6GOzxL+pgp5/fsBi2q4Q4yZ8kAHOUk
JmKLylFwHXM+xp4R8mSNV6YN67diiE+oyRCNwR+yaZ5j6ugKSiWoS3mgEjkGj2o5jIJtDYquu9EG
7BBhLKmg/msODkEPZXeQhGiUcxCdv/qT9t/m6I6BOApYjsJ3nvUvaANsVo4JkZYPFqX5nOpkqhvZ
QC6gS/eEEpgtJRbDJdYDJnuNSEL8SZt5baWkjFTgxRAq2jqgZYv5f2V99EVzTvxD219Gc4hJcdKQ
ZTlf/DsGwFX1I/GByjDpDQkfbYB6Yzfq/Dw7brgC2nhFtsubMKzTqM5aaIbo9QZjYS7DdezfqvYu
qNHjfFVc74S3OYy4RVdfWiMM23idVDRu26J0z/V2NzwPlKvAXjyuB1khlCzQtT7WlKQijZdq2p1W
TlrBJcvs1jl7sfEMJWnnAjy9GNHcsJIDshbhnBmTWbchHU5Q6rCsYyE7eY/SaHwHFDQS8R3L8gyd
kI7TBeJO3x/KmEbb9LT1Ht5Q/5B5eC8cbvvneuLsK8y3XYXjfu0lNrKxZPZUpYCjf74tXoef1pA4
hgp8Ef/Jhvu8uBm7ldhTRhQnMLK5OnakNgwH6nA0D0YT/3fU+F6VOfi3tcU3WoenhsR9ldMsOVNT
CIPS36LV6KxmdCiWI8ONwt7bGubgReUTP/E9g5ZW9yynDrRCSf2aViMhlY9hla3fxPwjQ4sDcu0V
WJ37tjnwIBVJuokDaTwUBpCtxlzqhVzc6o1T/Zs3pYw2rq9h3eTfKfGjNLGG538NieWri5iblu+X
+T7jB0jBjsrlM3DlTbWxQ/HCiukPfsdgc8+mLOYPeKmJYypTIYpdWzeYDCMuCIUUqYqbod/+2i5p
73i7tyOtzbDPKVzpw8i2DcRNi0BlJBHzPJewPqY1oBcUnja8FCOzKWjWWxujD1gyqee0WsBwjtWx
9OVjwqp6bHnXYgawImgvva+werrpccySF/79X18wScGSRVIMQ/87rJ+HNj392VU6xtONSgOpXWgz
eTDotzSGQ0jitYOrFR+D0gmWEP4xfGMDxH47mqPlZF2HZ3idiQCmnO6AEVmEiRWa69N+6vSknhpy
q7dMI9vkCyE7hGOsPEsfZ/Pz8vieLI1pMc0404/m1kCFlGyMIHMUiW5Ip+WT1EtfFrbEUZtTriAs
TmU39nmkkh1+3fzynDPOSM/qQNQQV7mCM+mmn/QSt+tVJ5/taEUVHuJ8cVjLwmzMq2BXAjQQwzJ4
xten1GR5644yeqsHxxmhYrLt9Rttta3RTB4CqVZiaCd6djOncWgsBMJ+dowC/xMKI4froVsNDZxB
KuOoxYwEfqde97ISlhkZbbYUEYkHyy+JK94gDzKqiefYQvFm01HjXLgPePVq5EHZyQfJ1cvM4xbv
6hlZM/GhaoVidC3W5KKWB5Ax0PKKAOWd86DNFiSz4QpN8HhWkovadMGOlarHGgFiRu1Xe9GWxWM1
nHKtNhVXcxA9dj97+ENkH/sMFdvuCooZHsoyl+zHtGsiFPOsTqePL82gUTkgViJbj3ITNG5DzdGV
6RJrutBkhu40ACohRCtwOqMMG9/6oCHgAGmHoDhqo6i2LMc26dlcxD8NdtWrf7h3Z0t2HsrwQdDl
ODr4SBPxigGdyRqfw04aPbCGO/v/YSkQwmY6Lq00i93dMKVwCsguTuT+PUUY1Cvq3i7KlPoeD19y
CZuMN27c2Bd+LMm+zW+koZgn3Vu05GDFtJDTBmERmZXA0yzogzP21mhj+qO1jj6qbMc3WychWElA
ASjOiPo6Fu7ttaYw3tDOQagKjwEx2Nn0j68cynYjyxM1X6j300q4axk0YgXXu2kUb6i4W0y8F91s
uSjShO28oWOBNHaC666OKC1sBcq2EY3BgFd0c74aFiduUU1fl0krFGrcko8EGb6PBiVYn+30bJco
i6i/d1lce8xwayz1XsDjgk+ZMNGhQGs/+6NGsmaibSW1zi3wx2drwLBjcAHbEzfYFrhPplIB0lKi
QOt1mV7DHI0Iq/aN8oeLpy65/lgvnfb15s+bjlxOVfczwFaQ36NKtKvxBFtvszQsAWNN2UyJMqO4
R9YO8RixrEZM0bU8a1J7O05RuTVG3QMQaDJY108sEuSKp5u4PcUz+VYRzs34jYR5648v7tdUxZXz
GTRiRakw4OAzMVIVzXx81sB09mR0+5uaKEVKDg7DRHeSoCWSccCt1OpwH2WS3loDepeblx8T6n5l
ojHUrJz6YbliPDQ31wMlgJJOFV5gN5ZHw6jQ07mGVFNF1+5RBbOHdGfyfyCmKC8V9Fepn+hf5VCn
ltjlx8nVLkFqXB8NtiWx86YqQlP5UpRuAoZTgBPYrJxI9030Lhx3TdHmSKCEqLsIIufymZU/xD1B
08otqRxCdN73F7lkxK1dLKsXxE4qL5KJr+7OdpuwohbLH/2kX9twjV6LtGv9Rr23m9mAt5Ur8hTo
C8OqRczUq+7rDtGYJz+p/ig9PTB26pt3bMVeQvzQP1zbbgI9Q8rrPJVvuWLeLR7S0coh9MCuBGc8
jTyc0/HrB2GdCCaOETLBsXDlnWabR3TtacBE4Si9s55o6d/Td/8L++QdHbTY7ZbffhHdvH8GMGBY
/YMOftE6yp4xpYAlz7doITfKf1twYBSPBX/YVqsgovgEriOFi+B948Omfj1Y3c8T8u2jH0+GnDpo
tIh1q7RlYRqOA+5Am/qXDq9Sg2LJ5W5NfqeSz+KQvKlBpGMUF6RbHIxa9sofbExjF7p5nmXe/Ewq
J78pfy8mSN4+702Sl/PmfkbNIQ7zivK5FEsJ2MVkFOe4foNh7hrMNpluyzpgkXpb3p2HDTbMwsDz
hfqTCTZOZo+LBuoZQYUkUnRcQOm+0JyAVGkMIM9JnaigRff1X6hW2EyijooJl5gzfZHeNOL7hBaQ
LQp4vul5neLIZYAUf05bgV2/R/uUnjvT2Sm5aBYFjQYcgHJfDa+8to7CAUNkaIsbhkGy4vz8lI4L
EAwZDGu4WnMy+tnCQ4EdvoYbwCt3nT1prZVPp8ZdAtbPMuDjZtQN7bYMJMcMRrHpizEDVd0dEQPh
wm7F5vWTu0HFlFNSAfqgiZaA0N8jRsesvkMPL8SwmekwRPI+tHw9YLAY0t9hFqh4kXNPZ9F15maQ
AYgvYNHbWPX9Ewl3IpkfE7RFfnMKnLtHd5+0OdLNWlZViaAKFrESX89k5x3tsHUMBAwq8YAaOKLJ
7fC9S6GCx5EA/+ECyHB0twQvN6h0HiD7uwY0eBohcro74ARiELo2aRwQ44XC9xCHsY3ylnC2M/qf
NGG0S7DWvmrDwVJD2jzMrK1MzdlkfmqG5O7CyIHlg3+R3vttfKczbM6BQKggmoIP8oHLXHrVNoMd
G8ZoIsXrIGa6SKQ6/hleIVHRUOeAF9oFg5c2rqNgoIQQ9iuqbMwhBFBN3El8sf6U3soZTx2OwBlJ
lGTzlta9j30bX49ndO1CvcEH5vSG2yuekZXwNMF5Y8HTgzPjHgVGf/knrus3xJt+addKB9s56VKf
QpPRsNnQcK/yGzV5HFR8SU+Bu0eJ1GC5BC+c7ibc5YbAGZy12PRvoR/l9hSAs5K0AYaNozEti79b
EcEU5ouJNyQIiHJqdC9QzlgpERxi+d8JVFu+to+wf9fbkL++ojxchlRU8DJ5eEuH08iVPvpkeVVt
DjkBc9sHEinrz5BEapX2PoCdeSaUI3DLcU/C8jgSin/1k2GOdtGxMweEAi+2fpzIPZ7PJiqEo2js
HcNPu7S/FD7Am8Dv9cERryz/Qry5t3zdme7limkzQ5K/tzC8jba1YZFpueecHEnXba07CszLzqGL
FX74J3Uh1YLgHZeIkwGWBLKcT2PSQM2inV6Xv2H9xztC1ymEktS3vwIM3mxeWka4WTbg9D1ArVQA
uiLhqpTY4wTL1fVkXLQFqKDHuy0X3+qLYh+nFPNcms+JKhKh86n3ZtFK6OqZebrBfvHfD2iZVfY1
Q2FVnjhwMh/v4l/5qNSdD7tAlDlFXoWOXHjNiQttIB4RQFLg+yrJhGvaTHc1PD2mk55epXfTHdFU
nGS6psUyrFmmIoyq3+A3rdxAt5sJtoc895dw9i0OY9n/YVWQq77BE1Jcwvg8NXVpu1C5f8r2C5os
snJJDaIvUZD4UXg0UrauARd0x+Tu6bHm1HRAP+5v06Hwbsu8vX1q7a9Pa/popKSAU+1l3+Dx+QCN
+g98eATw5JSQE6nMsAzCevpz4qnNToGy7fX4fJDtZGbvDh89lWQ4PxH01fSwz8y9gdXDJGiwZo04
R4JdVsZo4zrimpqKTPtYdTro0Dj6kpu1B5eniPHYr8/u4PctT7AskJGSL/5mBvPwr9Tfr2nhTWHH
OACdxUi0IyQcdaQzEqaXGyiYNAlbGbFjQw9eMZVHmvSgIOZVMmni9vCNs4dpW7vqkGbJUI3+2Cak
gegbCbbe7EWCtBNZyhPmUC/CG730UIX9TlD9/WmLvYd0L7dtQ4K13vboVtHMB7ANetNNk52rOy58
aeGYR+AbucT9zP+tpazNY7IL5fA9tu2qIy5h7uuol+RzpZq1ZpE+EZDS1pxuehz4F0TYRxr3IMlj
Soo128mirju6BBLYO3JVvplwY6Gs6JaukIeSGnKnUFP6hvllvT1kLPR1mZ1N6e7JCPRjpK1z52+d
cyzHMVjDxfhGXGsbO7d5DvV2EVmfKThp3+whGx0Fhxalrn9SsxWejmWefyVCM1qUrjbYGM3E5Cvw
HaeXh5i3kwZ41YVYCfCQvCNmAsoFdQscNjSJNKaNX3Y2FmdI/rAdNCC7qIEQkJjfBpR1y7i2//Xu
Eu+wngialNbmntSWB8vK3H/Z4CKxKOWgMmNtc8helCB1EptgNg6kN/cikIyJ+i1rOaIqDDLvHu7U
eWWNJYQN9/jMk8F84uAbVYiZF+59tgnruuQMy9gGQju5mQ7+t9dpCuVnsaXV2FfxfRrJB0fl2Rlh
+iHfMYS+o+f4KBcrKdXGenY/EhJO0snBTHfN7diaakQhHuHbqFLfT3mtvHjCo/AVceyhzrnyl6HA
jcrFHYAMTqzxqbWCalmn5r8leh94jAxBrrwgbXiqlhf4J8cdZiYM9RoznujxH0M6OOKh0PPeqEO6
ExEJaLVR6xDF6+qVEYlUZM4P8+KCSoI6jvRoHRW+lGNMo5R4QOMnY9GeHzrzx/f3rMRIXtyoX9NW
d8BGrBn0csNhKIoLkz6qkcl8bhxCb9IYILUNkZryg40U+VNTi7Qb3Nxu+PSLWV64fCkI3AS2ze2C
VNrqF8fe4c0NNl+qGxaJYDc/cW+MuS0k1LrBvUt6Hq/C3v5QXPJO5N6Su0yOCF6XpRBRKOo2Y3xL
YQhO8244sX/3kow6Xfa8UjscT5K/PKKJWVnCHbkGQXvj5IoEghyT2kM9S7RZq92/gODsdBqAPoEr
iVw251kSMc/7p0EusfmFSUo3c9tyf1qyBZurFMuJNs2VrH3QPftJpRRFZD901aaUzQ2cPU65jbPl
HaWzRSZPqQESvbMpP5JGMPAPg9eaZd5kqt6B+usfyjvqduPWinUxjPUQGHg+Yjjf/LJyEZiHVj8M
3STqW8Scwk1dT//POxgyN2iwmZ0p9S1GNlU76OR3bF9ZIwnmelNs2IhlYp4/HELGA9vrzAOSjVXo
dehBat8590sPKZdyhHFBRZ6CksJzwdIxoCH0/q7ZY+DNaVI+Gh385lk82GisNhVtdelFx6NH54NV
nX9qlqEUtic97zbxNdaLKAiIfYP5eJ3qNRfqtGG8Hq9dPO1d53MZflFS2pFLQ+M2HBd9U1pMi/8m
CFOFbqxa6VwvagMj5al7+/pAT/cuRtX1YIzKpfPSlDuwdNAFZM/oNYRSRFoeyNYWjwVe/KZg8wmK
44Y2Q0XCXZf9iXNI/iugPeXpXkLOeW5s35cKhhPfQlLC0buQtE0+tYpImPBdRM4r7G0zvKySFn+I
UaYkJ5qUFbzIhKdOBZ9wHyKg9JT1Sye+JxqV82fO4gM07ItKtcaUXsNUJvmRLH5mTVSDbV+1dcXz
KZPx1wNlou1/70rfx6Y22QX5UrmsHgdy7NMbICPSCA9YSfLxfCCbZP+TP5yTxnrBdlsFwqEdnnIb
YgOw8oTlk2VEKeV1WsU2FnIVBvcJUMNVLdv3Wq+FPgphqK/iCY5eHkdlZuaOcMQ39PCfYdhiYPDz
U5eUaiiRrksWi3FWkFKWGTChNi4mVrJl+2AjD3zBbUgBnsFPLs6+q3HUccDVNd7meud4Zq2+fJN3
aO3DVHJj88AUxPn66oCOS96RQyXrEzxXGjCO2uRMrW06bis4llW7zue1dalzAApDVZ30wKOM4QQG
S7Q/ZUx5IOoTpZYfEzvSUQaMRtXeWZ99mR6MsYxFykO1vMPwL0fzSBBvWrGsLu/fdcaRDjF4o6K3
evoNBjds5TZJ9ydT70sCfZU2amNyIrPINO34n5LZ8YmDjzcf/jcT9UUAKUksLMfeHyWEXEKIXLhv
fiz8Ra7taxPoyDZ0mqQBsq7mZ2IIuoFuz3DA6dTDe2L0ReU/6jkgwRhbHOvxgjrwwGdrTL0bZEbj
e7GTrlAzSd0z6JU9xwkB4MLK1qU2UeA5I4mHWQfLS7mXxUyYSbsLR1AAwXKtkrQMJcgVvBoDD4TZ
vUAeyjfZTtWpF+ZS4WqQSCgIvavpw/To4fzYh/SwVhKWY/aPo1pGG7FRA3wVrx//VNwzz6Ju+JBL
0Nb67kwcCC/hjI7imxOnJiF+phCPDVrN7mTfR9C+ZBUyUDjC6G1a1DWtFKPTCuynaR8eE7KQ93Qc
v5B/v7sSsXF5iJG+XxcXIlxCRbDNTSny1El80b0xvmtVGLnx+Pfvp1bTkw5M8MpQIpW4/0ZlQIKE
Zf5WqNBXH9QvZzPe9z9Vyje2TQsZ2hYYODPPe9PiK0Tvxq8fGEVaAVEnBJzUDtTPRNzZ2/cR7yL3
lm7pSQ9EtKfA1W1HNi/gehxV3cK9BlmWNEXsyW/A/pSQjBTGR8zf/muP/JeGeShU83XRvnKFpSLd
hO1yy0DDVauIrWnIkidKrJO6FRqxEIi5k70pTqNTttc5M+5yZUBoFVFTueTTiwdFivWJf+MO664q
WiYe6iHyAChN2wlOMQ1So4nfD9ik70ldXHgQdk+okRl0fkb6K9RsPvRunKhgDdyA8oAct6ZVprQQ
5WqfQd9ApPvBWV7guLGxl+kYj8Cj4Q0FSJuI0rasHNXH86IK1nNFcf0OSPYr8a2RCic+ujoZlyLF
sq7UWOwThDJQy6buhqUklqWKf/Ml4xoxR6Lxta/9JbprPRzPnskFZFgpucVBGHnAt5w3RRCdHhxU
0P2ClBJ8gOaSiVHFjTBC5QlZobsOs6jmCur3gO+i3FY52BVzn8UWe3KdedrCYynL3TiIe5jwHne3
WnqJEYByo9Hf59yPvHuPSwzdXE3+navxqB4dWFDTmnQXuqxfpnUsNwBy2NZHPVYbPQ0uzDaPu9H8
APO44laSBiEjGtJaN/e+UtCsCbyKK6RCFWL0vUixQcbdbxqSUCJBl5CbVMjNUonr67NBLNqbFsKA
RPDiuQKGJ8/o+UHazhFqj1+rj84wN2FLdkRDzb1d8e0tK94Tzx0XAirGDuiObTb9Gu/Xz8awq4OI
vmFXWeFpxE9HFHTLWqG2KtpIdTRHbVqGtcQEf2J/wJkJRfdNzSdZH4EDDRcm+Hfo2gp5EZrdCzdY
rtePcuu/aHVdOVzYulqYzztZj4thTIBZEhB6TSg69kkApDTwHEcpmpjz0sMvqw6p5LXcpqvAyPhI
zfTr5/LX2+TgvRkpPAe5FRG77S9DYtRr5QDljaWGd8tqRJftnPLzXmt2yihmocrXxhFOpVIOPhOb
iptZ5bLrQdTW7X1SYma5J9fXt0jd7Wlr74mzJlQ1MQFjwCZZamDzI9RWT+Ypuu9pjp5THWi6oQQo
rlCi2ZSlUCiD9DqmUrEY1mu7XCfHSAp1hVrexfp1i9IArXSCn9PkerlEe/cO6tHFnEwVrtkMy/Ft
H8qZ3CFt9TyN2YaLKv6NiBxTklcrf5X2yv4sM75Nn9YOVBfIoaxc7k6ZThEMtjn6OcoIBb6k/vuY
P57xWWTk/iuAr6AU+LQmGTcJmBRTxRW7yvizZf4UYV33dWLxtr8I+YQjT9SUcf1HE6QqHVu1/N0w
qnT/ClpoyLjeyT0CsYKn5DGkbXT9caPZ3w9CcSB9WrLKMZSGVxq4uYaIunnRP/LvAsmBfY804/F8
82BZ7kLlrcK+JQ0O1WHdPYwVNiYIYo/13TO34rq4CJdEFHrvr8OO/G/5gahgKNw7vTGA9gRqRQ7x
YcxP6+JGdmwKkAN8hAqzghrTdYCu/gGlwq3uv8UgAzM0RFHBXL2vUqhdVWGbA/WduLOJjQn4E5Zi
dBRNpdaGAsk97RLr1CvPAucQc9mZ2xaW7T0kgEHaH2I/jDlolbdWkMmuAZR7qaJgK0GWPxBdezWW
4u5KwBx4/ROINA4ZX68uRz8IwU8/X/V9ShHtIDCevpRSyt1p3Kh4OZk+DjxOv4mLHxVHMVTACULl
hk55BT52D0/JPRrCow9o03duKqDoc3aXcKmOxAAcGk2SMie0GeEnUmLftP7yf3Vol0ZDk6qyIMkE
sHuCyzfVNJiuI4HiHOCHzHlJYdth+3ZGrVca48FgWmmSsuJ1anHwCCTigZA7YuIVJ1X/NxFu6YXl
ym8bFPRZ3yyywLYgqOsgAlG6BQwfMjdoTtf1PbEs2me8LHaYWv6AhroxNV/yTL9bFqAJaCxhP1ha
ZeZt4xissm2K2lHHWLJAbBh0LiMpr9B4ri3SgNwxTGo3BLHKvN94afJT46YaqJWCTR4fySOdjF0s
msEM6yp5Veavx8JtlrlW75DqPxAhZssdN29CewG5CSQpuSvv5fyjoCclFgJpzX+DLxG2lBtmIkxp
affTzCP3YXonhksq4HmCkdomqSXv/sLmKmjHrxtAkKnY2kXZpiirRU0AJYtgK2b9J6XcVky8vsXS
QQIxpjCA/UOlRjvTkXqRVjjwHz3EFBDHZd8k2NZmyxHQkf43y6DJi28nHhf78o711803YrGl7mkt
+HAXAbKp9KsaShl0jVjmGYjnRADS8BOu2E7+QSEWkwuhdgAqfwNRUSR9Pz9qge0Kz/lRVrFPKPBz
o0+psZXU68v8TnKC+WIEth8w2fAjuN4u8b0yWXMyjRC6Kylwjq/886d7apVb+PDFcjsuHUQQ8X2b
xHT7xXq2GCwpNw7IBNI2RKf91JGXu4+6EvaE6eonCg5jSfLCfycnaNWCGQXWZUR0nnvr+ItfFwFQ
uTqFCF4FvnNEzg9v24ME9LX3GGtk2mZGuff38wDzOhu0wearwG3Cxpi+kDxfrIqC1oq6cdSf9Cxr
uOz3f2SAeCyPXRWcvyZm9pY1w5+iZzI4E7tE0dBRBtFpRBTbzkVcePawh3DdDsplqvn90R6n19wq
7uhhcNOUUZ9+eiJVQlDzzifX0A9Bti3X8+I5MsnSAK+CeV1OS09w5UuvMJx2uwDk/0GjULZPtLIa
K8D9lD3HBpE95gnDd8TZrMiosoHw4z1E6kd5jjomwIY6YOlB8xNR8TuV1ZH2JXM7Ncche/PYaVTN
Bj8Nc1C5wEMKLpbC+kDdzrz7Wft9HU0KSzlTZC9SPt5YWMMgp4oDCd7Uneyn5GZLhUyN7VTCtEYB
cQ+k1aRFQ8lQeyemJ2kmEqJvLl333o2dKzptGBMOCbA2NPq2Ay5UGxh3MER075lKQKqFNQaNs6gn
Wsz8ODVv7mvtqITyuCADPifR0fsYBF4FXyaBFMJZrG7ygLEHvr/FUPZmbGW1uSzJaQms+++0rJ/w
tAmR5pZFgxoZTUqoABXiB9bUhSs6IOXxNkugHZ/34fqWl8KRN2CaaTMvR0XEp+hs+amx7DYH+0rE
vlDDCCXsYmaoNOk0HiBD4BSwq7WGJ7fckRWciZSzeEYToUfgdxVNQUOp4Pj5v4PA3Ks2qY1aY6Rc
9Y/bUrCHYp1pxCWohd9r48rYXlmtN0LCo45/X+nqUe4PSL33b4kHU9Jjowfd5A8vIinmv5xwTaxl
31d3rv0EY8lktSdCln3Q0C1iYD9Hctlc/sbFeJcprhVh+HTuyOgS7Plb6/AfMRsZ08UEZG3kHgSs
YenPKmIndR/xBweIQ2PI0MN4OdiOtIdR/SjEdlCqcBgOTAbQSDj440ZGKXqzDAZk2/1IrmAL41tT
xhS+HXoDzOQFULNDJpAA7lwPx3KMos0V/8QKCVRwGuHHaLgC1awd4h6CKM+y2yitvAqoY+F/BoU0
6++hlrSaBhd3aB2Gvys4Tv50TNg4T83V34UuR6zJDdKL/ZWYASzmdonMR4oIqojACHAtt1l/WCeY
jPZ72keRh0bRmxKvRV2qYrAwVxIr80m2UFV4SxEIHBAyoeEH2yMAIKd0n8SqE+PYMaij8OcUfAzv
iBG+vCWFXAjyvK14CAuXCuG+VhNJ+GetsWHJll8qHF1ptTeGtRcXY0/hGz1jNZX8FS9g4SJiQksD
XJ5lVTqPbO9wEH293zb6ggICpQamOY0k5Hu8zk437BwcdMlSvLysjXdgycXcTwMh7TAttpjHt2Bs
AmRUrshopCw5qR65EG24qz8+TH8mBlwhi+ked9Egk/u33dhfrqg29+htvTlUz+2lGj+WAo58Z1gW
7GRMa7KXDulKII7D1UMpQXRleD301Grn+uWqNsEdpN8KL/jhVHMuLIAwPQEbPyoTdjBgNhut/py8
0KwC8W5oYWO0+ReaRRD1bIpb+9F2Qorm29ljcLImDgNOD4lrWcDo8D5AYJv7FEhtDYFWFafyI4Ud
VQxL6DFJbGhLzMvjf17Hhlwk2pv/3Ybtfui4bWT9ZDrSjebW476cJ04tCPB5arv7mDYPbmgzvV4i
MWPESs1PjkrxTI9lpf3o05Dck2IdAAvL9VLBSn62mr9txSU5gHqyW3M8hCgdBYeoyJ7XqKkqF8uG
RWkMkcAMJOzErr6jg5ixV3F2I8OH9wVa9PcptBGPU6gkhj+RZ0RZtBqFBFu0ejVRQP8gs+DlPGmU
Yz+7o/KljP1TWm25OXjvi0/vRXwzzt7yMDacVu+ywXUtDocleSU7GnX/56oB3A5IZa/M4ANCD6dJ
Kiz879M9NyQKm5OB31nme3v7bbJ/UXnQtlJ+xfaqyo6Q/VfTsprcgVIsfmD5ZgMJ5d/BncG0qIU6
mUfCeB7mCvB30xWWQRYTX5SQP2OUlYddH0VamejLv7sz7YGrePLBVBFDiPgem4Cpo06aBiiBOM8u
Xy45gMCzvzKQoEmp6P17rfpoymq8qGBcS+H/Rl1XTmEnMTgO+5SN0b7x9SReltZAhIAagGQLVPVp
bJgjJoQHf7MfLWIVC5MX+u3SaqWHVcC5buGZPiCkzwGknySqa6SqnFr1si+DDfYuXxUvrg0CyIv1
8gIn2m7yG1HRCpAZ89Wactvb87MwuTfPZWfYUVzU1bPcYPzdvcu68/xyLCP4QOuZARBZ8IhKEZvv
zeOSi4WC+jC2gjYdQONg9HjZAVy3Xf0yFzeEW+xhsSD3YBEVfGsiqP2TWu0EtvaGK4Q5/c9tLXWG
cpXENC6D+enaTJd72dPpTPpRJyfTRAL1fLU7CTHBvg7s7VRp+xcrflqenBeQOPDLnrG2d0mtsvHp
9HNz666Mb8lcE1HIYvqa8VgW/f/1CNFuA4JuAAxvMksKyOgCKb+u2NmneBCoOLF2AH0S1E6vSzw8
MHNZJ6hDII7rR2y6L93Uf3Ntc0/dDMQPEcGvF9b9SEcB/HgGBaAyCamaFHFt5ugzDsG3Skvy9/UN
84Sbz83zDXzJyad5r3xaVTVNXGSAnrEsyr6CGbj+P+Y00vJx74mP8Q9fP3hqllcNtFEFo6evKy4M
bfD9ovd61pbfnO4wUtZCIgCeZ4x4Qf0Qi6A7oe+7IObCkv62wjLyckBlgB7ypEBYYvIUb/qxs8OJ
dzRt22YKDarjot6vKmxdc+0c52mpdQkfKCqTAZIzgo42XQq5vN6Ed/9Voy0NLBZ0kjTS2kdSq/vB
Hq+GWr1Z59PqlyzoQ+nMD+u5Lng4BvxnRzZnvzlZO/JAy52N1DSQ+hPKftNzYmUR0Hxq/XELEWtq
fHlbAiT1CArF2wiKBXVel6fLrQ41Ln842Xv/od9Th3uWwiRsneg+aNoPuOyTukiNF0lzya2aPyRx
/uUe1XMh98FaTmPcBlxfn/9jp9xSS4CeXeh9930QJmTeBaI6EHajnXYnfX1GLT64nlClmHGOB+0r
4Ajec+cdM2A+8uJQwF40T7M+g9+GlsD458hRNLjkUh2aR1GIxS9VnxjGsqH9xpfiU0Bsa1IM7o+Z
1dJNp1XbBdSye75g3hmDkic+NkjpJ4xgiQNAcZyjQlCHaivUkcVSmdt6RHei6lo/S7dDm6AlwSoQ
UAUbM11+PU+YnJ9DPj3T8bxiqMMja5BwZpQ8SjJnRfs5S0t4LLvJ/UehZxDrhNZl/OYir5wLY3R7
nfQn5yCZQfIbIGhDg47qjBQkf50RmJipOmBNLcn9yD8UxVOw+jYzFMt+liWkBkAP2LzugvTP9F+I
4Zm9t1nncolAui9PM9NK7XXk4L8BnurZCcdljwb133whTIHC4Wk/hKs7c8P8GC3DRCZELZO4SjLz
qhn5nNqHt6xJh8GjR5XaD+MfD/OEEUSSUwLJImDyEJTVns4YVDN0QPANBZ9rvQbgbm/Kaw/5+Dmc
Lolb7FCKKkevQYsPI9Rn/7UcCJ2LJCY1sXZMA6WBwuqwv66atnxj09u0mItGduSnvwNUgcBhdoyU
SMYL7hkj98ssMoq69IvXlICwyrIL2u/zk3RwAHTCObzZ1C6IGfbmI1ABr+92YmGRr1dHT1QQh90J
R47PUUWxXo35L6ETPhXwfLqX1QxqANOVD+uonvmk2N7kw/tGZmuQfbCI2+wNmKPdWSDWceacsaf7
P5pL8QsmcY3ib1sRz57o/5JmIuwryk3Gf01YPs3JbaNQ7w16XLWvLrASQ4zb/nj40YavCvS0XvHk
jBCk7ZfMOR0YSYvbjYWGHpUYhydEmgsbEtrOKgiZfthqnSeW1jk1hhZmD8hZin9xks3elCHeFOoG
tAWeqtj0BJLYBQRxyf1xvRRIY8xAjhPRkCPmjIFiK4eSrLEpMhOIlyPdPdAT41p27mxs0/HPWyzR
u6gxXCa6f73ryN4CuKEDgUrcHc1yHMBymIc8N/oPeN03lUGVRJwUougstbt9aY+uthPHrvGpbrp3
aLyWEvOIzd5NjoZ7hrNiIcsTdFsr/gvvQfTe/dhNHI0YuS3eKhAGvBSVZ/T9jjiBKzCGOijwDRRV
Xyjt2SKrnFEja+quA6KU7c672mRSrIgC1t+P7uXrfSWTIy3l6jMS4SAS1d2ZbgL7XXIOM2NhhJVr
phchyQwNDmVWVmdaLrKj8diV1QZ3MIGN3KxU94vuCI9NojzTYDXtb8mgmPbxVrnZNh8Qp6sqe1lY
R8ReZ8699S6nGlJEo67k39yrsVg+Us8iCn5FrBWCfOHJmeb0lyPYj/zVTNX/hGqvwxcHBD8LaWHq
ZBqczyDiBsAk1wOlTXsAQ/lqJeNpt1hiavugfDq9K/M9EiPCUs66N3J0fLJaetOKHdwfWnRyYO6s
jl8S0xY4igZcLyetSlyrxgjhOIqQ8FXRV80NxK1yPfQVP6ReDQa2tWSZL8TfZ2xceFB70HzlH4d5
4PhxTZ/eh84D8z6WTL0lQr2o/q3zAPhfiKWizU/zy+lKeOYnlXPeh3P11Sdy8tif3u4KDET/KOrU
I7TJ3BED901lP9opVwPBm1Y/t3TRA167Ja7HKVOLUG8UZ3OQ8ZoP78lREePT0wbe91OV+oT1psJz
BXXVo1Mw2PaPLeU5M/lmTDYuWiSxByfs8AMspL2LPEpXhzIiGh9+ayauzUg9VMKwXEVNZEbp+yeo
NSWXNkB5H266oBQrSjFcjCXg4Oit7mOL863EJLhazil26Adzk7tE5Mon7Pqt1gHe9niNPzrz+No7
ceqjLSzIHUXJTqAIIZpApyXuO/q/J4zFENtZTKvJY5z34hOCvgHtldke+7lgX4p5tKSc87AqKhOC
LH8iPYzXD5kMoVuYpPfQBPPNcespw6GoMzrMStPGe7VWZjJie6SyXZtYZNt/XNt09EFqIZf+F3ez
I/1abYdxK2zS1DK0+8LAWhd9ZtkqxbqJz7BU+j6DTIxLxnzsHIinJmdDqojRbtFE+81Iz2R71ZVA
UubQqzBKtgXrSaVdnAptpcp8JkAUNzRCJYVdJ9bKep2zNZF1wbcXdBrbethYuNC2Tiy4U3HoMBw/
DX1qrKO6BjTk78BlFriSZFlsqrOEOqB+kelqgT4Ui185khpsnVvIW0OmdQgo2R3R82A0wMREf+xf
Rqiy3M9L+wB5Ij8y5JQAYNQUh66KcvWPGg0RXBLIECnCAfe5qybJ9BHpcBXzppncIvOjwuByg7DW
mnPawz3DLE3zfVprEahR3mlD0na9b70QSpSqPTfK0NKKiSS/wonY6qKn2jPfZpkTFYjHuWM9E2/R
+KS7DYk7kVl9Cfpjp2FS7TTlGNc7AWqxBzrsFnrHPnNOp/vE+yuMT+z+bjrCG131IHzXDpp8eDbH
ER1NuWDqs14JXBoMYeMtNN5z4TLVaDktSvmkv/2imWucOsdSJBGyzBHXPSYrPViVkE60hgl1tRrD
PBWi02QWDZDBeEbFiXpkgNS8fuJk1+1x7tENXk/RSB8j/5sZQs6rYSEBXhYPy8JQtWhgqmaRHxQ0
lvxFZdIwHloVLC78/G9ZtLOmPRImAnbd2GYdycAYqvUSi8NLVwt0MxRqVn90LFxvej8VgFPMWjaN
sfQk106dvrxIY5+qIWfZbQngWoQ9YDukee2QqNh/+SOkIJdj+nJ5mHaoN6ZgRC1CUkq7XetlCXv3
gqVTTWXnKXRVG56bWIBgeOasJntOJpV29uouGFmcQY/8XbRcX7n+Ob7emhhaNyTZbF+S7mjFuu2c
OGRaJ3peCA8xhpfUTsJC/bK7kyejEz8Ws9mnOnv/1X/nfQORbICuVs1kKY54DNT1JjRFw1ObZdV9
MouFPMZrSu7rJgEzq0GU4jtSxv19nPf/9BGUVIS2OzSd9lHddNpH9Oh/xRwZfFwf9xW5svKyTkmm
CEcv6vdUSRyTFXyFzSmBCd0CoQHAe/ZwzHlT8ioVFfXpG6s+vAkj8b//V3MTDg4WRQYo2LKVhDtP
GrxVDdt7kMeDxbm+Zf+ikWfx2VmwlgC042MLOo0entevfpTC58YpYgaLEvLsu20TP4jJ0iGFrgkJ
/y4GmKFcfO2Df8f7bcX4unAgIAlSibWHRzbngNZaPvscsXIe9S0wq+8KAbn/Z1Ex4oKB7DKMVKDo
68j1KMC1K1XH68NDbHZ/v/WVIarbaH572qfAeD/kj904L83/uULieszKVjEaOJdJ/174aoQaoSTn
b2W/w1Km5TyneNCglxAo4Y8sJBvi/235ZQWYa7SZzCvE4xn2gpN6eS9l7iZhTSSjV4sB9Hj4/ck+
Xj5uw5MEIXYaL8/GzQs+qFnBdZFD8qVyiQ5wj+RyAIEjAae9OZdcrNYB+gdx2sQTsgkHU8CeXNCx
jEKpqiHtbs8314YUzqpm240ar0zdSHE06SdU+WLRz6v03ldhvQ3q6+abFtrksOgzGaXjJNP2qTWS
eoirHtmT7JKU2j+VObeDJX/4w6AP9QxOG3M2+GNqkl4XD3J25Ksp+tynKwVIcbbX+k3sLqw5+k8i
j7YQGw9AjDngWwicmYh+MQTWuJD6AcTQc3F5/5h++YyWNzgukldCI0y+AsSglxoy4T0ZqcPIz2e8
5vNyfn4YoTfBFSWIh97X1jcAmHyLXX1u3SIuiLPC24w8lt7ikhydzilQfOS+Z9/xt0NPSE1ERRIy
3dcCu/Z92l/TDZ0juMKCh2rhiG4ZDp5kh2uBIzD27Bg2vUbMuxf42hZgdNhTg4cTjUvbAk6/1lBO
prV8J/xB+2TQCPnahOAs4gKQmF0oFBSiOyfdhpP8JEWOiL2mgQ5O3qnlkPNETYEoFd5c4fQnE6Ex
hMZ5b7LYxu2Fso62bAEM00LFKzLk9eqxsXIp1w+SYfYpTPDo3rn7GIV2gjRoZ74eEsHN76XtKh/M
ks11NdKAQgMEW6eexf54khypkTovNp9okAPAqeGwnCL3ZvFo5CToI9rNXiP+ofDrMpd5lOOAtHYJ
nkTFfJGu5Bmq4Bk9dLPePRTvvPcQX/PAzZCFmcycKzCgPgfjSioUjyWiwnRBuuxQ6VcdYdk2Ta75
3NIjjNPuidzHts86GnSS/Pgt/SAHYffh1HM6wntHIhc4zDJjzv+7u7t6yQeCwsqPX3ZtoZmRCsFJ
K/M8Wik0hWpHxLqiGWHUBVPtQxhfu8/qruVBmc2RjMFgWmUQ5ZvRufGizGw0XeeMc2EQJjvWDA9w
hQ77x5uciRa65SbNfpSvQ6J9beWZ/ZUpE1FGoQ4yPf1kdu/KOG0P/DkjuzfTtuGAPyPJS3IuqQcP
RSMg25RvFzxx7GdLuLVYh+XFRN/E0+NITe4Bnz5XVli7dO+i6YmpDxnzvK/PfzHg4rrtFVZA1aaH
myR7myvolvxlg1FYdXwP2YSYS5Sh3QrdYJb94Pn7EoPH61uAE/fuy6lQPNl0nEqg9hMNWmEPZ+OQ
bpsOTcHGJDjPvQATS8fGmE9uyfVUjLwyyo66QH/Nll24/wdf1pSs83DZ597eGkWvRO96LwaetTgQ
3xGzhyuTSlUXjd0BO5BSP8HcfEEDI6fPomv+9IW+uM/OUCl2uBF8FjO5JP+lT0wqa/kNERPhHsRO
kvcT1IJ8b7ZEBBeDUO5nb0XgC3OFgtrjEJ9lqoKiOmhiKp+0pJLKqkazs7HBRtK+eEQWK1MHQEH3
3qb+sFszADjHTup/q0uaQy7kQOWpwDU7kbaXK+5h6avxK1P9DWn3utWuYEWOutVEreGNK7MUzlmA
YImyuNkssfP3cN7VprCt4tc30ObEWeM56BNp5LiiH3e/rZ1kFoNtGtmIxdI54mhPYYHjAYDrz9AS
CNhQ+RfPpaSXEk7A8HzSlkkO0GZLvi3wDlVX/kflzrub3UdscVY4dZ5pNo+Yh9jI2JUZ2wBGojcz
mNvNnjykDk1ySlUEYfglxett1Ie9+C4d7VLsHzN/+tWKrWd+nc+MSwBlo8pe0xg+/dhjCG7MlD9g
RS0eiyWd8sUJX+8ON4ZioCtbODBASZjwJ5XD+9ncjqQOZFcJFbd0xN2Rjb0kX6gzakfTpt54Dn78
4g6Z7pv4mwz4l84IuZWDIKe9LJbY2HHKX3AJpY8BTpVabIy3ocGZ6161t4gEUjm1urQzMHgBAb4T
wFTvbHEt++RKIAKIG6sWQbi85HuVMPnC4zbZnYhLkL6QPfGzx+9rkSEpyOwkohWtiUWw5HzozDDp
5p2iqwpRRj6KaygrMUkUyUq11L0nKQkUPF/pBupbuDR/4lrTUFLR9wadZyuQoLiu+9zF/U8V5ol+
mU2tMumCgURAES9gEDAKQ6LlDgfYpZY42ldRhapUTG+xocwqL6AnayNeedZyflqpTYnlBs0n4DCU
WICa/o6wXriwsH0MvrTQ4deoE2qc0I2LmFKs7L/+LqCK1gy7XesGpsFSlu/kZTlM9EhKZoCNUWY8
wUvmy1t++0sNTrMR+2Ly5SBvcB7xPAwexVzveSGW+A/jolNDQ3Y5jBnseYGz0FqMciXzyj8MAA8S
jvOqsjzed9uXo/EyKnQhAzJiT3cuWunpI1HBGFwTBOH9cScfJ02uEeT7TiQY8QDiHirP/T6BU5Uu
bs3rQqxrTH493LbpXGV0gC9/tLRBqtC3EG/zXifg1Yo3MsgNeYr9MRWmHUZop81ta4F/Q74f3gL2
VI3aeowDonOHGUqriUJWehZyohc6Xr93Dx3IdNcFXfcD0ImrSzev8ooVSLBAG//pnJ4jFai7hbaH
s3SGO8BAxsDEWkf1T55nS3C2PMNxRz1FKCAFYROp6Qg3OWm8rGl9IrYdTvvyDGy/jeB+9wtPrDBI
kLRiPRKUNjDVi2l/6q+8lX6bUw15mj4FRdHyyI5C9ot1c1BFxd1sxnQIvNmHpSFBZHB4WXOEaDlm
N61ykXAbn+j1iqcoiIWOCIoIeMuLBounQICsB+HB8JnU3Ex3l4lF0Yw9aof2odiFDvoLVcaNe5BE
i/PxwCRwsm0vPNjxKtBK2ARsGVG/ZW7RscO2Wk6fYW+PYWIJZn6XT9R6jz3io0jtd0jFWPqh9oBx
s5cMummrwYHJofCPYEp4UuSQKbTPIyw2WNbHIFLXpdR4C+usnzkYNko0ro1RxC8NNHy0Sp6xyWfp
NOUrtpCXiXieQLbvpt8xMLLPAzIMg26B6+vhRq1zPoqudt5Yb/GhW5N26tXvGVzHLfJUiiSyKFyx
UlVvQ1dBwboW7gG/Ap+fTJ/sV6CmRNK0hjRejRzB9LGyC+CurnSIlzi29ZoJpZdIb8detWIaNMA2
I4YCo4uEucv36v0ngR0ETTvYNK7aLkofqjCHyZlAvOZbvtkzXHhbtCJdZxz6h+yX5zPLHPS37a81
4u33IUCJnbSOD06ImujZGOQ3O2QAoqCH7B9QrgS1ra7NFFQyYkPszymz5ibpwX5vHKOf8fvlzWQx
Clja3zUJBarHMNkxoo7QmvsguZO81pdw8Ik0GO+qF8bSuTzmkte9FBYIoAvqEE0zI2J+JbfANlYU
amRudkVOUSEhYJj4RZo7LcY8hdIGq7t9zUXkk5Ov7NOyE8QHEsRUObMb0MjOZxXeGrbwsJHFP5rO
lWhL3hQfhktwSZ5Nu/ixHaPkCRlVCIzZwRXOO3biz7FVedWXqkGAZMPIosC80X4LlKldXNB+4OrK
qnK+vzhqCXOHdyPjtI/hMHQs6OS0NawewL4LCEvprJyKfkFb68VgUPuXANGxUfuyHUxtpzym7sbg
U5zFNxT67olZQS67DZFFc0tb7dBfrelnKnXFG2scwxv4I754GlxsRx8rtM5Ki1x4CBHCCBeZms8i
oZHRKfxwSOz7oZxN+GPtZScg7PMcYb+5Tnw8E02nHutTIE/nTUNVSaemO5TTW0wvdXVfOaq64zls
3xwrhpABIJMY4MPxKPn0tJO1q+Zhq4F+D0SYQuAPZOlG+0kQn3tLq7f1/PjKi/AwnHaFCN7goek4
kA0+PHyAbxp+rfJz6Y8T2H+gjFcRxSdXTm+NgUabftjbCxgRYcfA8dFVLsRTT1wN3LdbGObYMbR7
2kz1rGorHZpJvoaigCZpqrVb/sLLZLryKlihm5TNK4CKzrAQL4uZwlVWCwYXqzPJs3HK6Qljmclv
1dQsJJfyCNxLnp3XdrQsPMy5xdVOp+NeXg9CrDtSvLaPyBtWQWhr42XITkZYTziiuc0pnps9SOGF
78BP+EmjI2OVm/UInVXV0wpFlsM3zudQOeI6SubVlEBG/uZIwfUq+V3+SmPpdAzvszym8omxfzbz
LX2CeuNW+uDLiSHeh5tGJBXWtOEjvYrOR/yrhPwK9LBejPnpaQIRkSKPUaXsaoHhsPMHb7a2XAiD
vEk7/dfCtTdhKHmo0L00jE26MaeWUAbSWSRz2lJU42QLbdagtJcZY5DZkdEegTYxiQbzqNhi5Br5
pi/EwWu9nVpKM7NC2LPZYBnYGXIqUWhGJEOLiNmt1Soy0Q2trk/lgkoj6/4SFPxXGStswGV3s3vj
Xnu8ux3MzKNSfvCUjSVtqDx3VPKhLP5bBHcbOjYf4bIaPBV16k03ZQzLsm30azSUHp7C9aOsMiwl
aOLU8zMqupGK8sTj5Cb8O7hO1Kg8sQRB0/7K0Jis7ncRIdTQtSROwy1SB4NhYkDJ/PlYYpCz7/Z7
pfC9KGq2dqNpdX8ExvKNv4101lvfp3yRj+So3w9PS5qiUFqA6vIZgkBg81zUPiiwyidbBKorgf6w
rXTXSk0m8kmXU/d0lF9UHjUYWxAfT32utouJaAaqw2jybRJPUawT9SGOUv8zIPs9pVAM1CkwGBUF
00S8C/CBnY2uASrII1tnSMv+Lnk4He0lGIzycPHKW+YZ2XmVQJzMG6srdspGjQAHgr0eDVhMnxf8
YifGEcM2a2A0EzhYBFLhh8RlQ3gafOvMYafjx6U0t9Nyv2b5Mx5bvhN7ILTGRQjGO9t5lm153UI8
ocDXWbOWGYZ9wuhBe8DAArVdVyu0TA4Mufd1lUgDyzWYEDtiRw/LWqcO6A0rYVPQcRLIj4i0tlyx
tfg0WPjTZv/1dZVSHY5m3SE+MJ/BqYqfbgcTKlT6FXCo4kkPkRvj8qRM+oYuWdsxpi41Kkopm/7s
tncjCGWh7CNvAQL0cgNTYAKVWi9QCPhS5cuq2FjpHzWYqT9lcTYXsQs7f/0KUkzHIsLVFEJLjN+j
Xz+vaMpojJA6K52+Y+njI9fiJTObY2PDFmNCzmbv4uMkvujsUzlCWgEdFIvN/T/Qe+DncJqU9CWB
UTaBNxCqyIsOND5oCXcYDoIQTglMnkOojOerMZ+j/6fUeCGUWo1dgI4q6CfaOJh8ZTKQVFJm5DfU
iqEGwfh87ZVrR1LRPdPa5a1+KzEPhY0djF/FRkuWfsCyHRHF2MIlHIctiigqcjKYXMzBAQq3YL+G
Tm8CRDsDHYktIaewD8Gig+PlK2qXvYciBAvr/5yeQoNmfk+rUPx+J6vRqKSs5I2DuV159wcdbDWH
sfjxpuxlH367YRE8WPZLdDOBl5vzYNdJg14SKocNtO4d0ANtF2bFZ+ITpAfcFSxDGVTmaKtdJVXB
EqihsXGl4HgPLt60JAupUQXLeDarozw/DZUje8KLHrIa1hHao+5vrzVU0jOIyfQQ1YXIOCRu84GL
8IolyJk4BGNwRwXqwY4Bi1VVuSHvy2xJLMbSKmPG1e9VlUxO79gQCPu5PHnClswkGYipdy+gt762
HmI546MiWegmeitZM7he1RBwPPTuBGqIVDJDF0NAdj2Pm4kUC/zzyBgdmn8FwCaDuZ/yIuyAmPUJ
+5iBVRpBS8449NW8gqtwZUH3gROyHO5Z9g9TsLzGfR43Eey3QpLIaehuQPNoBfNaku0me1axVKu7
LyrJ+M2fzCvR6qRqxdW3z/OFrhvFoBBkvf/HRZYF64JM5vzWtTEMOu4+LXWq3TwCcP8u2wPZc6nh
zn5qmv5XsfbzHcP7yJJggoBcNt+Oiy+m/wBlMAQhmokxPq4trr5cou5fAb1SbR15c8EkB55l3ZvD
O7cWojCpWxm9MKMLfOkmnfrmqVxtu570eek+Lbm1GQQafjt3+eHu+qu9/7Y7Z3HC1utmfLJ7rxmn
71WguLYvuikRX4UvjDO7Rg+WIEFzkLIvsKfBBqSIgwwbR1nWvilBwsby3Jhc/glxZuu7KKYsQ0a1
OqU94IhKYbZAjLkR55qlaj0b8g1GHtR9hUpjpysUHcfPX3NmthVmVd7N7dZjFj55w/sMETaW9vBP
98NCMcFfqtdUM494HtYJdcjyi1PKTzCYTzWhH78uwTTh+LYF1Kw5QFG/0blJC/1SxrHhk+ylQ4ia
NKUFDhB7gG4ECAthBxKlQmSXwtzDo9XDgbfcb114X88OuE0/VHD2YVP1T7XmAJCDVI8Q1dWeRoeX
8nDlDsQ2hVyPBlUdbPrAn/D7NjrBBejFQdBrhG/+D3YiDegVunmuQDxwyjz6YEbjsT+B+4RH+jDZ
0L0ge3lArF/eI6k8Ug1xDPK2WRYyq0Dw19HdUFmYGv249Ei5T7U4S+Yx3rVYM7/BOygXT1CfPmki
ZlwZFYXUsMoQalSkpStBvlPKqJ47Pu6BzkhZgldnEw7akW5lcNWduRM4/deDzY6rqRsYRT6qfBhT
5/kfcoFWSy2Tpr4I+dWRUkQ1LQa0R+WyQ0FGIRJJfMnFE+XzU3OiofRX2KI3iVbLMbw0BKBKvgKP
T0bi3mHLppBkyqsu0vv05IajkPU5NJS72BaZHMw2jwODI5K4JuYkGqd/3tDrq1/r1sQjD4AMozdB
Zmp5KD/TkuqgwGFJdkXjz6ZY4orSqxVPj4hFSQojU3/IRVQ2UcmESBfRO2MU/e0XwqdQ3Gt9rmSg
VRuunZxuWhdJSzFMkbgNSaWRuxd7tRl+RJ13W+ddv46EOiKjmrPsAN/EwNyU26epE5uxxCBwZZ3H
2cGlz+scdJpzGIbJdK3QulHAVbipouS4uQG3p6gsz7x0dQMCmSa6lE45W77fYtIGvVwC6k4TUTIK
itGTedmkOHr4i8hr3FCKK4yJVzPgzaGmSTzn4NXYvNU3WmsHI3LAcS/KP8NmLJ6xQGE4h+D5wrsi
6kEvXkyeFT4oxedtjcHER0eOFsKjIShHOlXP4zDCbX/l/9xTMMReA/2DPuFIPBs9HR6JvKkDwmkO
pS1TFtdJEyc8oJ/Xk01eOHCaLF1DmnVesl3QBhT/MC+JK3b5F9JqxdEq3mHPzgd2I6VsCyvBlF/L
JqDWCuSfCqjSOdyGV7+T/j2/lzfizd0Uo/+diHyajHqFhNFPYDL1/mt/CDczLKiOdrKWtTwsE7cI
mnxOu5aX0BcUffVT3ycGQ4ue2xQiZa6x1DMs+9EweR0NySa4ibdDnjvCenGdNczSNRyiJL9cK2s3
mniYwvGcVIjG6GuHxNBd56C+M/8AYNYFVK31jfcnBXuyoakoAcEcoIP3MGmu1ogZRfU+SdQV5eK2
UJGlehSgesHYanWzFr4oxpPqgwlSl8egRJ41DMxygvkbJ+chK6uQJCCigxIBzRCZ8st/fZaN3HRn
jtl18oPgUXhS1xyN/0k1ds/3TjL+W/j/mpHP0/D1Qwc9PbjxCZhdFt3d8bJgDoBKOLpMKbuMYTqh
Mrffbj1aV4QHiDa47w7hU4KZKk58Wa2y1NcHdNxwekEmFu/qd4E1qv8RVNUJOU4D6+UNPnmvCZtP
nfyxMTWWWB2GKeUKjTMXWhy9zeOKDc99Fy5Bkz14v70icHqZKVnEuLLdWRrO2dFb2Nao1G10iXvU
vaMV5FlVWbJu8c6na3p4os9scG1qQwp7NHqIkWZ27/mjnf7/vGE/NH9m145fcUpRSgZhA9f04eMx
cu/U2AOVCqveo52dHYQbs7H24a0ln3K94wMyNp+NO6ToU87rhmAc8FmcVqolx1TNK8vXiR+ioSDR
IdCLkYnHLSt1P278Mxh2exDXAhjfgrA+flNxj58Gp9rR3c8FBNlTIFB6SIjqyCnfdO2YPj1oq4ZV
oWT7hxCUcTJiCMzrGO9Dx4XBst888st1y1FLlt0bHrImNN0o4fbVhrIdjMfhwCp/7+zTSM/k47Nn
9qcCDpA6gKq1NEcOEwVtAgSp+JPp0arczVojwSw7V0K56OoA/lHtjLJH1xRQ5EtRfpqn0RmIEHBt
mhnLu5gnR2gCTmlYyrcxJql+iydFTeoWvlplTss8szsiKNHZaxeRwttVna9TsFZ7Bv29NkFUa9el
+BicZATc7N1i4Y3T5QYk4RQwzxBHAJDrs9WU5OUnUPAHdvrKZHV4hqa6PvP++gMBIEu9Gw5SgPQ/
pBf/O69KV/vMvdKQjFvBhF3X1L+KbSTEbhw+UHg3o58mUAlWBWXmimHbheyPi3U/rRFFc5KyRsSS
gUsEETIA8z2/4jTm0R/tZzXqSRo1N1/reS1lFzA06aoSUgvMtygA/pLk2WMP5et8JAeVzSFG39BU
vc74DxV+0S2vbAz3tUYGK9t6ydspP7w1VKT3Rut+ipMt8ohPcDbO3xlxCEwKYq8JZ8A44wWP5j4i
57SFlRTbRGHsVEVgdFAtpNQ6IOh17vq4Ih7ao2F6ashZuWOznJdkqRbklh8MEWaSB5FAb7adGjwe
1jI3gUeVoilboI+6dAE5s/3N+9xx94dUMCOmqA8EAG68s3CNdGbCErrRXYkXI3wpYE1WhHzWAxy9
H2pYkxWe5wTwyyGPOIE/rXexkW3yYVkoyulZxYSAhwKJFOMx5/CnAbq2dsdI5oxLfzHPuWdApFuH
fMCc+5Br0BlT3JaJUqV261qcuXdtB06Qcfw6+49+FPHwsWHSi7W7bJ5JtRU1MdA0L5O85cSY6IXr
RR1lhVoAN4ijSjNByWR25VoTX8pQey7VtnmQHc5NmUh9CEEBxf5QCCo4lgbJRk2/fFiQhWZqRKPm
Voil2LzKZeKj5/PUWQluVjOO6UBN9h6cWlYAz21P7oXKV3JIwMPNGzcECREzyodKgeAbOGhS0Ktk
ApNQwL8kR3SAytqt4v6ey1WFTgKxHVNYxOkjF92PhcegZwMXRBDUmYtaTlwIvMDy931x4XBt8Xsu
mDpYYqj3Y3sCDm+ZkMEr1vZw2kpzx/cg6h8OXko2qC+s49I8YXPxey/oCOU2LsTi9zqKg7e8FBFg
DASWQx0Z41ue/N6DCPGqTLr/wofdQW79OaqxvsiqssRDazfWHklopu679UE6J2J3UL/6PHUg/PnN
yBTrLFTxMEmC9+IofXwdaIcdL0rARr/T8hNCsN7QKXn+Mchy6+xIS4t1Cl0MGCbPLJh5oXr0bWqN
N23OOt8VXhxViWCLjDRmRQY5QHIJJGZjkhMrNz9iDLoBh/AXGyngLDrPboGvRVDvqOReXtNoF8II
KvsBEjyAH7SCkRkuduAcEMEIsq/avtd9gpY8jW1iKMj0rIYwZnbvl1+4Al3Ary5wfWtw85n9fiVI
0wPs0Rh0Bm1M8gWgfXVuHNC0A7+oiZlbuh06GfdEEsvjyQgFPJeUiQQNT2erGRQ0APw9sO4qabZd
btSmULBhSKBUFAABXaF+4rvkBAO04GSFLYO7XwCp4rRPcpI6jx6C3FJbBfvlGeH6xCRiBw8mO0ru
BjZkEdGpYAUVLgOV2IEmBHXHUqoKyJ0I/WxzucnGBBdajTlHziu1MLdqf6diE2rB6rrwNgSspZAV
/ek+WaLAC/ZGlATz2J0I9lZ7zWLFfbaHgaYDynVIQSvkpXpSnIc7HVYimjdPhE7LCX92lgwddUq6
BkZabKUc4I1x3mPt/ylK3VWHxnUV4v1nS5Qacx5tnfH7FDbQpnSVr/nNoyIJNlZKEyWokPalfxDQ
yldNqeH/g9wkCacE1Qo6xAc4ZTII8HkNcJW3r96ldhsetw3a/CHevd+UE1Q5jt1RdcEaDbmZeZ3d
0NefZqaK6OIBNmrhTjvor0MZWDMlG6SVBlc0klQ9JXNS66H5NtageH6tzGeBRK8tS0WT9HcHXaB4
nQjeOp3bovC8uqE3IOK7sIZXT7/6ecApcgpAA+6wvOLmAuO8RTUGUAjXb8snPVwAt7ii4TR9mxL/
yxPsmyNCmmEY4fn0jalB6WXCK8Sw2jAU9xqXNmE0IZ/eSwVIhgxzqo0v8zj+NvPXmQgZwtAYPEw6
Gxc+j+SdGs/RnWiBHh1E0buinLuv66IQPE+WC9eqc2peVFrv1oC4nAs+NFxQzQsp2V3Mi3mcYaJ/
Wgzz+ymfTdmcmtIq0Vzkp/Azm9eBvPz8iETgPFKSz0pXtQXYDv16dCi3r0VtGyRe9EeCDcbjHIWi
N4Extxlo39SFr4MaeHUw3+VDH/HeHje6YAe414RIwluppzrpouwFcp44VZeY3hVb5Lx9ooY7AXLc
P8T7+Kelp10S14S3PyojA6Io7umerHOmjRCYxw9GC+L/wMYTdbE1wVWJDppLnF5T0xqadQWHgYyV
vfwgNZ4x8qeXZ3leHNVg8ulcff8vMO+v5xCf47b3k4DaG1ObDAKtKmzUAPcboo1rab+nuw5DL4IC
cIjHU/X7qtNeZQTYAvPf8XufB48YCT9OTATPFAUD13tLJI3jdVlILkYi10S18CTTtgelCh9zw3/F
vV81MYuJfjvU0o5EECoGyyuWJbY2CX3y/3r/lA9ZTEp+/yWS5EOfvUqDofejNJFKgwdYzBur5Q37
z0bGiGjvfl6KI45BUeO0ly+oa7Nd6JifmMSAlXvAmSy8vBeTCp9gYT48B7CNIGKcziHcaNI1nuuh
OaJpiY2Q4u6AkvqatqNv1cMhMo/zkP66XoAvYcvB+0YkTueAvnv9b8rFIUzskzfSUl3iTGVyvJy/
5EJe9b5TJ3ctn8B0/I6kcyNTztxPSBMKNuMbgkzquUDqaFLNggdLedw8aIcHG2hBMtm+uDDLXvHD
79kQUZONgv10TXG/4rTh5I0SiB5S/5cPiofhyBMjacFYiLUtM7nfckkLCd+L0y6RR7U54E2bIA+K
v2PBY0bH4+nEiPAYYTy3DCSl84EQKtpUZtbGqGbHnKUoj8GKS6pubj7rfiC2/iI3LtbwPQII/NWX
dGmbU4xjVmHrNRkTEF8G5SNdBU+Be9/yZ6LAmpY0EDFG5hC1VeemiHelYFq5jG48pJ0Y6qCgXWSG
Vk9W1F+G9HV1mD/KQhDKTTpm68qSpZk2fxHFDoTSFNzFyQjpKq8HHXoxH1/Aoixzh4K63aDlcY9J
eWPChB5qMaZp/xg0cR1eX8BbnXuSkYFHF799auqUnOo86CkkEXaO3leB++2LBBCCTer4g8vgXFkA
ml0BTaFMudD7r4dAaszsGpjpbxlooeUnwe7XtS90D5dd1WoVAcxk40Ffze2grLqOFAz35v6FQwxx
92KPrKGuK/H/d8d2ByAiBBAQdmerwXFPRngpU41PE2q/o9HzYx+ueD7LpszvPfNGNeAvsDoc9/WL
lFuTuyPhajFEEf55ZFvbCSKB1GLS5wowTGePnaKIw/mwIxE+R1H2dLMZKUZC330GiyDskFVK3Ir6
6xIl7hZbaJMLJKcMBj4HA3z2fa4bT/cCDV39ovwmcBGsAYUDuEA1vSmtaVowoQeLPEnYrHl2ubXd
cToh+jbJLvhp5xWIhwoM2MA8sfibNF69W2ejELOPaANAMw9vDiRfx2GhkuYzjWtcdaFLAXUX53wQ
D3QZlI8fS2FMxd3tk/1cO0S1hyyff5HrfTvmZvip+nngmuXhPgutBn275oZw6OMzwe5PNoqlCDzI
LevfxxL+O+MnDrsdaNgmm5zW3chf+G4Js+X5zI/Z43KWvsyHHaOiXft1pkmuC67rvKLlEM+Pmn1Y
TqdaZZWmydiz4FzXIySkydQlj9U9U0PBeuVl+hmXUemYobPU3zCyvZJfIZiSa1uDXaXsTRCyeL+L
JYQXTEVcdWuejgE/Aa67csazSAJ0dJh7SJX/pcciTg5yOa3zNAUdb2TvLPJbtBIL6oIpznd+zuag
B4mFjvyletdmq+eOXo9WpnuKm+OT+NZvjEM08GfG6BBc2VoHsfI8jfOLstYfU2sS/9nkCiqJ9md3
uBrrSJRYlThC1ZKmvMyHLRMELMDIsYp8Q3emRNF6/SAu2ckUyU29qSjhbsthojrvastP51p4mB+J
H7n7kXYbVBKhOTrU9NBxDfE07J6e0Fd4IFJhXoQhrkGsiuY0aXFQc6ScqyUBfOXRJxraToxTYVi2
8VoepgT5A3rLYcppymbRBvd1pgiw9zDx+r6dGdaWSgnY+8Rrkmar7+058BOqTetNnbKGMc4OWCLZ
NKbwOotOA0mxd+oCgBLQTLTy/Y/vawyxYGe2nwABPUrOg645O+DR82tlh0NbOVR4ixPSrg0aWwxi
7BR5DVt2biZt+d0OTtP0igMR9Fm10x3DMH4Ux274ZqhD3VE+oVh5m3gjMXGJ8SAKi6ufbu25OD7x
EeJFDQY/k//hH8Q2ThRUQ3cE5K3OtmyQ8dmIndKDQvU6Ae+ST2/dImYVDx4kNZvEMseQbgj6/j6z
lOv1ycjY8GA3glAdlhRKLQlw52ibGaTiWf/0J3/XHQ8+UKMPZZnhn9bVaMwxEtzfir6v0DDE8+Il
499vQMZrx+qPbEOD5uRhLBdZEVmiHg0sHsmzH3/X1/WGu0R5mb8vScbTDfzSbeqYKIBGi6JTAwq7
55FNZourn5ZBGIGhHBNoTwAjmNQK3UxYQ9llB/QMUU+hHYYDsMYYKwm8Tx04JL355vKTQi2sxRkI
P4sEN9m3zx2B9cGpoLmwiTqEXuHoTNGe2cnCTyTtPcL/hY5IkjSV1rLYY28i6WXLIKXYq6XtJy7O
WpUYO4hiO1iyTvCXhRK/5X+MIRJ5jlrn6fPUNXaUjSufc+LAynRd9CLBfyU3KtK2gowf+WJLQkJs
V/2OC9mQ8PBhau3DAlnShhDN91OFF7D+aUqxuHMYEGhlrFi8lHyZnJw/+/AMELocJaBP4yWgLqYX
5jrf8ENiRqOeeEIRrnbxe7iu9xgH0kAiTWyOguNj9nN0Oat4VcsD3eV8uTz3u3HpSwLnQa7TTgGd
rI844EZPoUHpciIzE6LdkEDWOSGV87zxZDdAoC6iPzdE/6kYESH/tRpKFRZPPqEUjhq3n9JDMy4L
0P10kjLX5o/7zp6IuXLhusixPUdM3FNbE4drPtbM1lYHxpd/HY9aEwGId6YW5CO8lN0J63iBOQjl
zXfVjT3GQM4Rl5y/gSjmu4xOQzGQ/aKhY+GOFZbXLr4VUpKjT2IVSjnGSdXVDmAUnwa1wjDtLQhI
InI223DcZq2O7QsEBZIRuc5ad5r9QWmARmBTjHKqZJqsXv1UEg/oM0YiE2FcHv3xhtDesTi/Cwgx
+/hr3J6iWjoW7EGEIFm6hVowPZHrgqV+xodlh6ScBQMgNjwZUlN1PTf2OZ70nKOaO5OIZZ4hf+6Q
TtuP+TH2tnHX8sAuCcyM/fE8SvptWaJXbpyuuw3r+CgC/stKmePDLRsopt1MniR6sjYQYGR6/tQh
6S+6qbZQmk8nuhdn6o8xfG9cmO+G2IRfqkz/hcOiTV6QhFqhowESpSKwPlD/T8qEPoAN0J9kDgO2
0XLX7GzI9Di9po1PZR9Rp/pHPWlIMllR6M7cLie+nHpd82MY/yZkycERl/FJX9GNjIbmY7ppThG8
DcEDUXY83PMbYPyaaTTMwENlT+RXuGUk5MZ1qE7GtTDSMMuSgXgQEhofpy25NRtxnbQMdl6Mndcj
VH+i5EZuAh30RNWbYKcHAYkmRcE7tRGLBEMLc+NNUuDb11DG4ASaJgdTIkMDnspPUg8v4ZByghtw
ZCa8drPpfymFqfTNzAI7jGMW6Hc7wC1Qh3iAnQbOSr7gaMxdfoTx9gBIDhnizrEBFTqoYWqxdMfd
yqJlIOW1jv6gmmTgMuUr98bTIfq7ttQd62zHSnIMK8fI5BzzjLysB2XVKed6dhIpIlR2Jdq8aUWE
ez10J//vW2W6nyRzSvhaF4vc97OryfTkJPpMMFaZO2i6DypIF/xfVLqCtimOeKw9t88oREjfE2fr
1HUL7Ycb08Csj71eQd+BEG5IKCtg9H9wyM6ymVIAZtRD7JKE9YaGJ9QE3Y9hsOMbRZpThp6txCoD
IjfXKrthdpuZWeS7yvHMrLF1cCPq2UNwaRlucnVnPPY5CiTWT6hvySMoBVCgGwFI3DSFBTSeudd7
pYdamaYQpOEVbaptqSGLdTtKt36+P2AzNHMYLm/SMFxsMqsYFQ8ftyUiXCqPLLTxNKXc36WFLbet
FrPPeHRcr/A7PKHbGbXWb3B5a4Zw5rDxQfDkxrllwktGCB+0ab/foDEJpRis7tFAGKjt3TqosYHD
uORY95mwWMjGMLvUFajpMnVzucFZjbGMVBLUttXjToiOwM/niQPlh86D1lQ+HPt/xmh+gskX9r4+
ejfNG415564VXASUB75s2zQSO/zsEH7CEbXkkzoRX3KUwGmWzWQ1+q30WKl7sttwmBdjaVwTrrPg
15R8xhY5kgPs4jQOHNFHzJBrbv0dcF5Mm/ZmaMgkL7iHVTBDQdRwbNb6myKo6ekKjpUs6mBGS51o
2n+NSDd6FcPuyK3fNjoyNuDQuk/HF5kUqksEeTExo0WxKnno4MfemVcRnf9D/sQEsJ7tqswhcBc+
uYVQCeUxSf3qyQTL7wKVcS1BerBcx2FUB60QM8iwEAbgg2Y/aw1FOn+F4vTw7vYVznBfUhn3bsfa
WYQbVEtKcitoR3R1nalZdP2ooo6Xb76xvvikO/0BT1+nnSKYtyRy2/BIQkuz2Pht2E/aT6JuS7TI
bTPvkkOiI1K53/T8yv9jQQECIeEzgCxhRQScmpW9D0jY+cJ6QngM9QzhWQ8KcnGPhjw8+MdtJ+qB
wAK/DISKcDcfCA8uhIAaV3JzbNzlUGiZce3wNjvDF6JhiW1qLHmV/UsOeBfkqzzzHt7NsPi9re4u
EQKduiiOxA6o8NFF0tgOdamaoPVc8tMRKF3Eyjhkoxd8kzNSWW3U1IRVfxjqqH9zUwvMZ/kINTQ4
2D4WluWqHuZ9gWNMOGK2FqbD0d6szEMRbte8ubuX9EYXBUmrIUpy9fzIl+kvjAiLOSf5+52kI0Jv
TsNtIcwEC2yQduyRqTl1QcfUfvWTrmRyt8xSBJyhCoTxJiSlOwQy8rooodwXq8iO849+QGg4aMrp
sXLuF//B1nfYmnJmn7DzzA2+llLcL9jlFjxHSjv6emX7nOsvU9QKZeW3Rg6bmlT6bYthnJpROA73
6ZYwZsZ6WRsWXEusZLU6KI/FUbhkr5zK4ddCMYGROANOj4HY4S5ki/Jh7x05N07FaNttjUqIMZ2i
HmFWzIspC92bwfcy3MeWx4YwizpAxcaDIEbV0WDRkn9GCfa2cnn3Mlk/lvgHD1cyVlDWjLJjiSk9
n5ePwnq2CLc8AQlPAOHY0ROaoB0UOfYhWl8M4zoDVhCVGdAHTxZ6cRPl/zk96j9Yolez28fSF84s
3UHZ51R+AsKg8uw4e7JeJ4wJgguiE/XQwGJp9C2e9O2eWj622SkGrrg2mCt+9ixPdBxuKg8p09o1
4R4lw1FthS8EH9oTD0CwT9Mrm9sggmPE2FsSaTd1AxdDYUdaCjBVJwPGf89crCKuwIcSmNvZbqQY
LWoiK7cTY2tzyVBA7PwFRCZ8meLVDbeJabUg9f+Rlp2B/wVqLsEgFdwtBWkJF0h4WD02nbPHCwyo
oRAU5KVl0zdX5cGwyCuS3pWOguptKJ9XtJaGPWZry9aRs/a/Zd/IXLvLeHhB4pPPZM+Di/CIHNPp
1f0h/4TJgePGzkfDyQZF9N+B1vOBfKl43a+6M6AM6c9YM98XjxZQ0Co0cv2Iqv2Jcar3tgGCmsrq
g1TEDdjLjEQc4hJEfu2Z7vPtzsEvtX8cBu8ikPWLBlnSIyidavtW1ZXhaM1cnTkrtuLcS/i76jPd
9PK1uvFqmYCsgvjpfescKMuWFxLe6w7XECOg35UELKTIzJH105hCTvQZa1POkES1spbwSDwhSSRi
VQMBgWTLwTCBACIwtmxQ82NjINALHnBPiKeQ+HvYQB5HwBkXyJoIC6VXviRcblAo1NRlI6ExerXK
n60e+hvV1W/8hnZxr2RteEg94CIL+/8GKp/lUT6I7I/X5I1/dyE6bXm9E789n7SJaueWX0txCr4j
z8kqjG14HSM60fzy+fMt700DRWuwunQIKimVieOMpDqsH8f2fMcCo/1ZcAeG/qGJAO1nkYsgVo6N
R1zv+/KtMF4bO7FyZ+XmHPdXzxJ6viNcz34Z0uWNzo1iEODfnF8UCtsGpTSqadHO5LdQ3uj1vUoi
NdbZcBBIWwr5F4XoAdDWLohwSfhE6zWKtrrk6e6nW6Ulj477diSoMyZCGeTT6tbCVimuTiQMdbHL
0gMOJy/jSxoUN7KxuLa6d92LZ7BlRTUd5XRVaxC6nVJv1e95suB8SSUyAH68W5aSXBvC9ijnOkXg
2/+ich4SocSZzPCRL65m8sKD3dU+H0dZWUxBwUDxgiYS098f6JOiecd8xGxIKo64lLENljkZKj5J
LgDWZvFL3qD1rn4GBdmrFn6E9rtE0NjWHvOGyyPuCRe8/+xhGcNwQ3cs9rY7FbGLV5+JcWgXttFQ
rtR5CejE/lmSFT3sEz4aSuKG8Y5USMhsOihFyper5USBPSpZDfmFoHaTUDIA02EBstuPgRIIwwjj
es2s3mvmBmCT5fMqD8BDI46YsUSS+tAT7LB0q7iSyaSLmCDj7wVH1lq9cVZwtUwpweKGtKwe4AOd
R2ry3DWmcn7Pg+ldzntQLuT6vuCS9qWb5MKA2XLE7uEdyic4Aie3J/4+3jH/lTRvwifAUkuLO8e2
VZkwqQ2+ibYVwjvTHvO6ggpEWN4f9/MHHf+vrD7KPSSVFJdNyEaNWDMegoAe7ZmjpI1U9i2h7dmw
p/Qd/UkOwA0+iSZESj7jM977EthM8HzZj7O0cv0zfI917K2uXNkMtUrX1PJMY1/Xvhqi0Y2BIque
l+OWSIG2aiRnpN0wMFPjjU9sz94uBlGnwbG9bNDzn8IrDm356AymVSOl34gRdMhvVVdEmgktOClA
u5RWYd6md+OwNIevkOm0KTEtn/GW6ek1pRjR+nbgCNR8j3dlaZLmBedV4bczS2GPxBqfbFqtbBsD
3nQBZfKz8ZrbUNjwBGIKSw8/1Xqm1ctkhrT3CjrpAq+54yzeZyLnHoOfMwnihk1Zzk1X+P50uoaS
YhbmzTK+w4pUpXNNq7en4h2EZmmtCX20bQECwF/s/RQPs5HzzRA6jpFjAScCVqv4hT0IYgLhQSko
ApmT/i94etu5Gg+b+6N9yRpQ7a/Pj3ePJ9hXQxJ27LTyIBOhOYKmGAZfc5yIs0EPRP3c3fo9jVNO
BeTsE7hQ4Gy45dxv9feTBIibtPzdLQgIjrDUQe/3MoUMUAE7utbmtdPAO8N1zD/NQRXTrjjqiANz
xltgRUR9ll1FFezeZmJs1kgMRsASws1xc5+lAaRv8zpwT+vPMaLfFAhr+YqkYQ1tRdkTeOvm7aHr
qtPbeopB8scPw/tzHAc5/Q4LzXircq9p9GiV3GyU8C1O/vy8lbXFFM2IhmiTz0IpUcv2nPRf8har
NmfJFOt+3J1nrqNSoIQFw4CtubRXlh2cAW9rFptJJefBJsScZ0Kjc2b+IBlP1vaMCnndXCDjEfos
gqGtCrRhegi30e0NtOEt8J7iplnEUix6GlBlLhk5Q5psPyr4uajRMTApfZdSgjwqU0yn7mAHDlOR
VTbsUiaa3Zd8An3nor9Z3Ou7XOGdR6B5dcFbftdfjDB2b+kp8lmxsrTBLIIPWgy+jXf92wSIyajR
sEsi+Rm1OcmjJwZEyCJOmMCHPkV+n3e5oasEd9KqoQT3qtLYVhky/iyTIXJRHQm3F6rC8DcSirbf
haxbtB2D6OejxKtcDVKUJ0ClNulAG3xbSxEs0wpUR1ZoPyJKowO0fm62S9RcehrzD2Hzv/0iINZg
4ddZrGGBKqGiryYu3vipGBshg3Z1bmlqvU5+gs0aI4xN4lprngXfgu+R75GxxKbixjIaloa7xYp/
EMwYpBvB3uHRy99ehwswgBxVJVQoMo9dwA7vxMJhfrNFf3aN25dcZGnl1qf2nHq7XEV5Ff4FENdd
jcUCN1PVDaZcFpDUKkurO3OqfYd7lsMVNSKuux3IPlFE7iHMugtSaKfBNQ9qjNY5ElZGdvEW9fSS
s3/asSTXciTkhuRK3lO7cm8dOhSgBHL5iSY3fvmFX8IR29b42rEM9VuVNL+zGuNUmhEANifgNI9z
wn5jdTKn70+SJdHJy1SWawp9Fsumc3yro0/9E4TLAtMh0ZW6O8C9K5AoDosmvgSkfI3G1WEuxaXX
sYzKoftUAdNKTX8WK6i3lH9OPJ9V5pkjVD1GxnBdmOy+ZtMLxNiPp9C8x4e+ZemLJ4m9PgdOGPlP
/cj+11RwVlawEO0WYlflzXEcYHAs+Jw7WLqYw9cQOip0srDwT4tYck1It9xlM4WnyXJ4KiTf4wSu
OIp47ZKOONEPX0OHyAQLxeBgsw9xGJdBbcaAA9ZW6lINpKC3T+4UdEDtkqlPiP9Xr13oIJ/ellyH
1covi5kbq8dWnp2vl93pkJ/Z+KyBPMG0tjuDaE08CjavAi8QHdmtcJS/j8n2bfVEQ/UW6UtbsE30
pSJOyYkreiL969OgIM3tfm8dzo8USsz/ZxGPaAtujFPYVCgmc1PiRjUUFlCBUDSWiL2hJ67LzXRU
mkVrguZ2PXdP/JGDiHPX15RO4R+efYdE/Y7FjFemVwJgtxYF8egRcfkrCRAyhu9yjBdmOv1aX5ke
iUlUAaP9XE+iPewNxYWoXcXIxiGk/rvg9NbcsjwM7ThAdXV2HjB4UqW2/TP8jheRK2jj5tmPQwtW
Hn5vtTbJtElnfDveM+pxBUvXgc3Xj3zVhLEmhlH9TKmtG+QtVcNkcUVwlryc4FnMTSUFP7RCt7iz
lwdqboQdFgH3Mi8GxPPmLlyO2TgZtkmypWcAKYfBphxhBzMv2NtfgFqYACEN03LjPzhpuesB/RBt
Xhe/xgIVmGe3PciKLPDvKjj3JAxeotcBbOqQj5h5SLGUwoiVLO7HlBiyqWVapdi1p5N1tFgwg0tO
VlXfiDVKfN59YK1xH6HSK/IGTtbobsrfDh95ZcDU7jUoPkPYccu4U9we2GHIoT4oVgnAd1xSTixo
lq1Pm+XNDKvtzncoEVgEg5m/Czi0Q4GUfYNumaSm1rooKO5a14laSQ8aqVOO+ySER099wMfbvZPS
dqwOkH+A3HCjGGB5sCzPYtaTavUF/XvoXkurIgVGSYs1NKG93CrzgXLNKFPBylOaj+Y9/1+PnBSo
7WvgBN1NOnu+2+PfyygIzCzWU6gKk2k64ua3cJV7KzW02R7LcHbmPGOKFZyoj9BRKi4Ysoiv/iij
isVVEjECnvgXFDmGkoqBpCu6es/l6UBWO2ny9P/m/qqM7klEC0SEGkvTinu0d4/wNBF7Jur7Zs34
RJIKggIghvNpF3btK9SRF2o04cFb1/1cR1+J2p981PRIsvCo4lTlPqhQiaedSXYazyOSE6sk4x49
TU3M+UCR5tXvGenyAU1D+9mh2vFhgz/EFuftRrAZFx6spmmUYTWztAZvXxtaLO2XFh/p4wesHyqD
5vtjZccKmSLnPst4djOdBJnvZQ3xq9BvTiYLBQrJiNnPkgcI5mSI9lyLiJjcWE9qkTaEbyvso5fc
denpTHlqzgHUFfJ2IvekvH7aRPNuMV3ssL2Br79xQejJFnhujg49A95Fwdk+LzSASUhCbXKLysr6
AVMLv6aL+ISJBCZB99fboV0FrpsigiQcTCcs9gX55EaIqhGlKL26UvJ+d9YcJel07wL+dGxoKWwL
Sg8UR1w4viySNQkDRNQdftAMafWw12apiQbLlefQmYqdmEcCJgxKvyhqfPwybxjFAU5vcRH3qgnE
4LVEbrG10D9QtrJdxmdrjPu+igwenfMlU+G+FpGuENQHqL9eeZOMtXv8vBnBd2no94n+f1tPMvR1
0dIEEwF26Rp92t2vUEqZ1Cyz4CQHOODZJz93XzdUtfohmSZVNOxWzfBBa0BuhtFG8WKv+7KWpFBm
SowUi7U5YbQP+Jl/pQ1W8CptqsmlKADUgBCEWm+IleIaEKH+X6+kjViEk9Cl1kyum9nMeEgLpuue
9qlMpXZTvBE0oRtFlxV5ZOvpPoKN305M7TIQJh/lir6lVrpNM6W4xCgt9UXNxx2+79c9X2V8Rcyu
3kwF1cfIByHwuIpbt9EhI9e10cfWZ1L5QqQRnmIx9ftK3cSCAasjo/HZurJ9dGf5KPj1eQNlDYYA
hNB4EjisOkTkeMj+VV42d9Ne5lb3JscbtPniBPjK9Jn9+NWMeTVYfA+ANdma47YbLt1Nnd0Ielxz
VT0z9TJVsOxeuoQG0bGeL8PtIP96RXYCPi6p/utMn2Zlbz2sTho6JT4c0O7W8LneK+836fD7GSU6
17XPVphWWnl6Y12ZaEDsFRIqdEFmROmnj/Z2u5na+OGrWF9yFEwHOSRZLtyKaY/OUwUKJ5NdgVoH
4CEIuJ332qiTr43olEn4urF7WTOt+weLIhGUrgMBlcullra+w4ISOJMGP9HJb1Situu8MBLYPYU6
ttnXje+13+96Hnd1BJ/tEJWtlCtzmZZBkyqEFTYDjUsMG/m8GTyiFip8XtjNGo51WwTmSsNB8xTh
2n6UoOR6h03Cn8UC2H+KJN63Zl4d/PIEvo7CulDPNB1IjMUhGcMgWarSnDWwSi2dfBFBcNWCtoul
W+aLYHnjSVJE4Tu4sry3HSKDIXq7OqVU2pEaUz3TZ9J4KH1cgA3y1jxMTVq8SSHkgrv6upw1ROdM
/5AEt6xEm8wu6rEUYw3mqA4Xv4BYLHT7s/DR+zLEqYivtGlEk3svvTZI3ALBeiLtV/AqRd5ioKKy
88EL2/lVi1Buz3NgHfUfddyXxqImFN25z68uPO28UD+dLN2uKsB/3u7OAw5cogzA1YoEe6MFLIIW
jM5JeL+hssKkAuFxZO7qUP6lbZ687xe0igWPNZ0IDxbibJvL1BSeu82nP2OJ420wvBmcy6aeOW30
tZIFr5V7lUupUtiuM4A/k/lPZRLGNrRosb4lR61McID02z+alXGkLHclp2oKIJVNqKTmuI8KC5tp
jJ/vZdFYIZzowTMj4m5Px86deVuh4/KOURAf5wmRZYUxJv01eTZHiCkKxBCTwfwvNt+vFd7cq9UF
wvxeN5/zyY9BC0KZH2FjxkShTNkCHOpaPU21ruxIKue3pm2Q4aLNYavOdiSrZ6fzI/c1u+48n0Jd
+GYygtD+H8n8TV5SUGE9HFD3IFB7S2ljXMsYN5UzuI4TyLMIbAzRzduUShOrCyxwTEx1OZFHGJtP
9ZaY56gV7sIuIHDpL+Bxf2krDe78rhnNQRJW0tU17STQW7vjB6XeJMeqE6ctxVgKyGfudYJFLWQE
aRUMF5nvZydNgsCm13v1AUn8KcT6vCMYUqAUp8eCAlGhGtmMCbG7D0UE5jfEFxI80uusSvz84Srb
k8HjqiNFDx7aVaSkf7AljXaRgKLiLbAsPK3B8QW8QnLVRkCjYppqRKNC93d/BRvDSU7zlAnHmeMX
s+KmgYNaEY2jeYThX+SVZLsRsRqsDs9xfwRPEBBJCNtBiY6C+THf1k3kKdK0pyriOg6nO+4ho7+P
6lzmoAqQIgCy/kxrKiWXgD+G5EL3bUphv5yj1euhQcp6DypTcxwoWxhk4fjagndXPN+aI4N0MRgT
8MPX754DUpcmaPW/cklz7MmF5UpkO28eu8HVJ2UW+M1gqL9G58uAcqOvxJGvPa/kybtuwrZMsYtp
0SSf/1WRrV/nN3f3DcoaajEDvJR+fwx84ZBAf+12vJf2gpXVI6qVb26hUUXXSJFrhmwHLqtcXdDr
BjBV4hQ3fkIWX63/BOXW24W7Hhpuq0av90yxEgd/ZKx0SqY6r2yjU8iIqDzuRG/ckdVdgluOm8CQ
vbb8D2MIIZVgcBf2/tyQvRNCzsY392USuhw/OpkUYfyq64ezuPN667ICABBth13WR5MO2X9QVnC/
eY8J9SHT2u4wjGnTvacnACx3WYsry7WPjujBLZzf+c0qKCzrwYL3821e9yxJtNcM7HS6QQWUBOf7
TtbAF2ze1pYXv1CMBw2CB5Zr7fDXw8CE31n3kN3QUNI3UZhmPcPFQBDGl55j/51RuXocScugT1uN
4gOmtNAayu5iLUqZfTkPcgcCh8ryixCahgMmZqnKWS/nzNgLqW1xSWYA/fvXqk9ow8753fuaJonB
qZr5iKDdVWF3S3/doHC4G+ODPfMNWy01D1glsCvCFJL1RvN7lsvYiyer1v/KioWN52N6BeP1k3N9
oaNVWimeWsmacNMcWGWMFQ2t7KIdeiC8pNrwexoWGeS2K/BE2JzIP3vPmC1HDMNmuwGJC3pGiwzv
c818wH4qisBTsBDlyzbwWFxvjZGFuNveH1AxjeShBkdeDhAJdxMz7gr4PlVYx3qjjwzNWtSrKUfk
/sfq/45XVLmQfjLhyVfscWN4Mv7nNf39+AuHIrw7NMxw8OZp0YcWLmG1aUTI7UrItB13Jj85z0Q6
k9xDHOJsAEX6RUhV7uWx1PqMeV91h6zGsXn9yqXVtNvs5N/YE5ukOjbkmSoFdJP4sUKo5p+eeG9M
HXG2oSjyugNrZB0VzIhCGFdWxAF2zTGV1L94pT+9vPhDsXzo+i91bWeiMKyfmUZGWfgFakKqXS03
3uHSOE1SQTzgEO1RnFwRrry9wQTptnyOX5P/tr7A0gM/PB8AJQNNTdEEXxixFyw/sSYmGw10GTK+
uJ4ZKrEEp0qkSSZdTGzoh2ls4vmJnMOUYQ2/gQPKy48A3J4RX3ARZ6njt3qzjjuE2lnfv3SvtYNw
0AnlePTOpdvWisVCX/Utp9u4VbXUDlag4wp48NCRbuJSrSbZ5SyBGcexaDGcTJ6NRs8oqm3nCDQ+
WpUsOvQ8IK60Dp7U7cssi11D1eqX6dBmTU6uUMqoJ/yb5OY3ZeAgRr9eA1uhrU/CTKlqjoMLggM1
mD8bGrBF3/4yPX79BdskSXAqvjUEtgGq22aeKWWZQ7bvdxnHoRmIQ2ARtS4cfbeiDt18x8iWUY0K
Xbjv2AGT1/68z+2f5DzvKz1j3q2w9is0g9W1fIJBHCkZi4E5eYBg18fSTnorG+7pUjj71zkL9jB5
XVffKc4Q+UX8VekL+BdKSjcoBV35x8t5u02fOBYqaOrE53ExRO28AluzeLkmafHDDnG8zcstGgrr
FBmZEUPOSDeAeOlg9sE6Nd5/Y0j5sVr3hxR4ELxNls1iK1mEDgdrrLGz4HNatyp/xGCyN5A3osKf
2tkCl2aTHAj0aFE3Ys1IA+RmfWk1SErUQO8hIXS6LLx5hJ+pAXaR2a5r+EHwS/qbEEniRRmm3pBz
w/VnMv+Xh6C95eFzhxeCzyj8wruJ0GWlxyHI+ocp/nLrdSI9BIrITe4Yo3n6DZQDQnltZnL7e8Sj
w0/UpkpGaO5AxzW6QIJ98srLj4CjWDiK5m0XNK+ldpUx441jnW49zi570iBQ8YRujuQhUmoEJcsh
ylxJtoQMtQHpzbDPYJ0grTnndJzy/hQlM7sVU015ZCDY9hHva/3Jo7q+c6ezGaAfCh8RXZpV8QFD
TwuBZBckvRsz/EP5QSvsMz5u+oDvrhTu2X7amgLYXX9C1NYxtqkF3p0YfbK6kMib992w0rdouFeF
kEgIRRK8pOpj8GsAn4QXuCbPEtLHgd6Sa39Vh0aAzfa8nZigIck+hoqP4/riu9B16sw8rN80LnVc
zOFW55MudS9afmVzSXU009n3/EaIQTdhPeKv0mZOz7X+cBZuScCgNlSMRmaeKCAiWePR15Z8dDjL
r6zYMXa+hvvhP3YN8CnHie5mgxwc4oFUUsp4VM4JQrtuFA50C52ftFbSvaXPpKuiQKC1d3QI7KT8
Q+7kZNugwWLrtBCS+9dlVKpybYhVLeg/X6DGerEHtWUknuAa+lCrNnzlHJn+xX2X2ncZKy7wecZj
VJp5FEQ1b3JDmGTnqmSDMEOEbTVAOZVvB2s2Bpr0RTmBAtQEHNxnQSbj+/ocwgeqcm2mLBGuvqAp
92nK14NfHxqmLCnZxx5pgkUOhrNGhIVOAxlHiTxSOUjLM2zAQcxRsiOA9pWhr/LFsgf7rb9AMP1X
CysGC1I9iB3IRn607MEWpVh0x/7DqMxyHWWa5TstEDptU0BFKFYgZAfdKlH/qF3L8dWtP9agSA+j
fq1EmST1VTD+1whnYQqKobZKRJz3YSW7A1xFcMq5Sa73UFuKbVUY5maulvM/FmBh6/jTJNYj4BXc
f4VeiQvs0ExNN/vlGodQthne1jnjDsiLG5OuoZDM2auDzstqwJzKxQ3oq67ap5/8hEiAty5Ee7LX
Z/e/Y1XXW4n/QHN06T3jsJBKrrixnYQREPw+SDMRM+mgcr1flnhupk/W6g076Ks/B88Vk185PkQU
WTpuZpd3+IV9whc7qxG2uPAAGr1Oz29fcdHx/Yzdgx/cCTUnOEbSw+j41wdlGDGwDktisDEPl4NM
rlOiEYsR0WrfNDxWoY3w32qdk+3xztiQ6o+M9G0RTgg64sZIocUuf39DXgIem/7UV530hIp6MSkS
u9OX9V8bXO0SXlDZpNT5iQcqQtb5vmuYm6WyAKh38l4nWQijktTxnpfq6J1SGLN7v76XSC10/SWz
vm69EfV8dgOLaHe7Hb7fzGWS7q8UcL/F/hbAS/ddCxRT9TjH8TH4BjG2oSToJejGJUeqVqAGbpbB
Vm8zttvH/zo+VoDivi6dLpl8xCf8AqHV9q/SjwXT4wV9EURSmjFajs2Ue0xuehHLKrvEfrZHTBf9
6Yx15zer0HA1RUsP3z/0/VOjB/n4o1pY2xkng8/qItI2+uC1hEIk4R867hIUBQIBlnSgsmEKtTwt
/JLvf28y7E8L7ZVkqsgZFbeSjRjo6CKl0u2f/nSjfJZKVtvj+6obY+7/SfEaTwfarlzNhvLjPgHZ
nCLDd6iVlffh8CCALx+3UW5mGIJrHwyxxVgo6Kv7OCxlpSuxZ2Sm7kKprabpxC4invy0wonDsgVS
EKs2r3Jhny2CBSgSiv9xKrS8rcOYgLxwCEtvYn3pXQpQm0iucWgWgeTjYgzL0969Hpqbx02lTZnw
r96Y8ArTrq7ljVUKuAZ0MeUZUikHA22yuEKRMxfMXd3zEx3dRwe1smvD0MgLmzqqCnDIG8ighPRf
3VboQU5SbMyCeDrD7DDTcjWokIZVdhg5B0fKs9oYkidnNDZ82c8YqIMNPxExl7+W5sLF7jtDuQ40
46UzPmWqRmgCfpUKIx3v4lkIRU+E/dAusrZeW6+a8o1+w0tgJAo9GVtVeWxL8BFyCTmv/lNeSP6T
niq+2lm49kp+mkQh8jHN9GZcWJjUbSS6MRhEpS0gkApS+9NzPZBojKR0i56elT4lvRBtbBOQM5Fp
6Q2ODD04Kkbvesiy4AlPdu+dzhJJ4YVL838LzPzLW5UP8bE6kRwMsgN4aAAZyTg349Yd9eKUZHLR
mxzL+m2s0ZskrZfN2Uxj2oyTQbcvNxFAPapHmeJMuytL6CCNIfoJJXa26obuPMWLtyutQKuUMAFr
RevzGD2O0G1s5AjyDQnfebvo7lPvEMKt2kBZ9WcbELSpReGOrApsjgzMN6lb182gL3SJbHUDiS8J
PwCfWNgnNLxfXSjHwSKAL8jwyY0BFNRkgGVTKX2jRM2oedo9FmlZ/3wFQq9qdh5FQ67aUjE31gcv
b6Nunz/6OsHvAADlOeqzuoEk+0qqgVvN8NEE2rXF/SihgP4bBIG1tLMkW7Ie8hUVcDbuBHFtD9WN
XYvYs1+O80qoo+nJAZ8BJCzhbyVYn9yOfEkCw+3ZYs5IFotz0wQA9RHa9PU4d0RP0+o0lwPl9GmP
wr4oOwAdhnt0kzOTCIspVCo5WID8kMgAQVp/X8w8jzgW1MhgEy4fASVRCHxocRR7A4pkwq6oflUd
vnU0oUCsIRmqX4gpAGNeic9WNBiC6uZba1iCGvNlHJSGAN4jqQosqdmP2YxdLgLuK633ZY2Q7QgH
GaBnDknfrjMpitZb7GMjEfRYu4/mohwGx7pzqPPCo78aPg8BWKVAoOXzvUDxZAkOmfsENGGJ8v5z
E7UNFBfEyZzh9stJllgfiap+3io4SlWnB3efdDZioRhmpGBJIdyUTv1meDofZmwbxcuVLuEyDB75
mCfjoGlOUlG1sIN+NQ5EHZuM2qhdaDwjeDTCtnlFrojV1aUOWwcGxjeu8oCnfSxdgvPDSEGQYYFx
DzQEMZ6KeGSlpcgM5sSQeMio1GfBrpfQcUmElEKnUKD86qAMFgeINWqWxHXofeybAeVCzYf9kvJ/
81KOsLaIHaLISjwSMw235NNqgHWJtlR/xCstnpO/CB172mJQTT6+AwP9RWrgVxM4Ft/R3fqwMPzu
ChyqDjleNsryvZRxtUqmSzT9SutWpJc0MEujnXTBtUowqo9KNdm60W14Wu09M95+ldszZprws9kv
ksrQKt4oSa2BAek3NpSxP/A0xJc64CU7bwiXF8GVYT7xslAdtBfXjBOz91cC/85F4DPrpUzz8Ca0
4Sl6aoDo2SVhO7c6oKs6uKPKGVuqD4iRrFtDNHGiaypvl2ys9zt34JCuExbh1+6DoU47c4CFYi50
4HFvKfEiHT8vPAQLZ/l3g/auT1jaqBLb6RRpUbaEUCA2EHglsysG4t8NWn5KLwEUcBTItwlSK5hJ
weJuCARE9YkYN4JZWi+eH3WnkB7RqGkG1PvZVy7DsIFo2EQgfA8ciHZXSku0jdNnwd5uISGdo2ex
2ylFxhB6SImCqlcHd3tW79w+suoITSDzd6M0+KBtLolKimILAI3+hb8ucR0kJa3H0OKGLAGXYdHE
sScB1mCMLJOUmk2poadFOEfMfwnwM3Ent8N+Iyp7HQlgjRpWiXFgDZx61jqWg8VmXT5LRaJsuEsn
ET1HZPJQ0iqOFdjwxx4jnEwnOualrPtk3GV5kRFsX9R4yL1CCI+b8vT5AgstDggWALjVD9Oy4URE
RtEk4UF7c4kyPQfcLepkBZD1VBm6W1QzqbpDoSLlECMqmkKbWJ15LXVIN0miFejuMLgLX6TczpOE
JJMunMghPvzXUhdRV+hMI9oAgPJqVOTNFA02Gxuva+3/5InzbnKXw2uvrlZewQG7YfL5ONuW0tJx
p0Cajy1UxAc0MlnZ1Ea9Xxh5lHDw85OudiBtIB6hWwd73VuzQdI3rjUrTMWfA/L8ZtH+kIyJ0pUe
a90arRK5D9fSC9tkQr2c0bxD7W5Xz9T4VGA7CEXr9hGiTNWXME07X4u0I2t4tdN/yns8c3S6ofwk
6gDz5cygc4RE
`pragma protect end_protected
