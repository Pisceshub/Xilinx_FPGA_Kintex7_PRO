`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Uatrsv13d29PfrWjV0xBAuQNRDsPbF4aoQzxzjV2rs48Ydkc/R2QL85sFEXhAqHe2RcyZbml3v9A
SL7mZzQHwg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BS5HLsrPAulryyaVdbkYq0AtWS73qj4S8HRYqdhOuD5vEdvQLRBakqn2wfNVXEj2qZmFQUSo/s8b
xES7ClT/lyzciNkdcB0TK9TaECYqepSgJucz+cDQHr9JLL5et1clt9uBTh5hkZf1nO/JXLWOgi7J
cf3zXYFaRbrnI1iGPDE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ad+85FI4YSUlgtCMKb4o9ZRNpzaM267BxC2ORKVlmjYD1L+nR8RxkNYIlg11JVM94kc/lNBzipom
feJEYOBy97bdOzoAaQhjz6lIrNBeYMPDqe9su6cDDFwX8jn6VtcDBLKJlT/2loGhbwK7w6xbwKe3
Anqid+3se4xm4ouNtpSqtuKpiLQMA5ThJzkO4KSNSeTZRseCJajZNXZpY5h8FSVZcnLutC+OlDQV
Hi/bbqLq9TbNEAPqCmkaiv2nPUQb2Nx/2omioRSxOQZOAkkz6BaIWc/5NulcbeyDI754+jrX1IzP
kKIucRZE7EQ47vLczhbbeWc5k2wV9CRskzVzMw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Te56zBdwlSzrkgzOJvdgD0vMQDPNPyGWfW3jfmRvi+yNfSdQene30bK4eS+ZgP6iemEHii3kq3uj
7ceRBJov2lC/U4oe/4rXSZ29SjyDjP1fHHiJUH8WIoTPFNrbJG3/XaluVfig9ifZWtvSgpq6uGvm
JiTJlVCad3bDL5tTY/hsKCYBTmgqQYc4vyssul6eoLmhpniVCsakmKkNy2WAO9U5Pz6ioydZ5QJ7
G6FZKw8t/hxhGiIRcW/TvsYz0wNi73X6bZ51Jd/7niHRWGsuyam1u4VWcr7MPza4y9I1jA24ifP6
9OQYJRN/cp2HZfNo91qVH1hODGTVz3YoCuoUVg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZsHbUEaQYxKsaj+XZafU1ONMpnmogc7FFymoYn9XgTapjD4CsPvjrDrdXnNzjeLnhWOGyrH0IAqJ
LUzE3ZWbAtMVz7XNgTXJaqKh7FGFvTuIxbieM8AvI+4dCKevh0d60VEY7H7mCdYYDokv8Do/v6ke
akqH39hyi5wtcsMRUYIT14a2tBpJo1YnUMw11nlU/RNJ1wANZWueZJ/oubglSkSax20Pl0IY2zlc
G6zM/mwAfWGM5XYJuZIqknUgdE7jcQ6+AJDECa7ExTNxZE0LQRN9GQAg05sfANLruqoKYM/N5gLe
NXO4Ts+pgESnJjZMvEO8VnUXwgK5tNzY06+yvQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
up68nxOCdEG7lushuPId9b7zLfG/wfNNF9NWgUqYGWUspqZW68zcWImE5CW/bKZewyvCtCQQJjr+
E6b9gvlOYPC2wNFlIycwitlNbLpoQgEjCKFj3bSK3eNRaGFXxXkbakGzHwR9N9cOKbhGCwDwb8KW
nih0+eJPhrf7MJzerfI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nJFjdJVIChMGO/riX/ZCL6QvLC889wkAgevfIXFpF9k02Ah0egIutv3VZhheNQgNKYvYU6c6BEWN
XLbAKll1pzVFRRn60Xd28BJZCDbDCC0I8tLjOtkwEE3D0Etew3E/siFtDyeQUqKo7oeRq2Iaao8G
4SnNM8GyzG+9rKULIYE3Et/PZT2jyhuwXp2gzCpvprrc73WUBxM/AhFIi2JjZcH/6XZMQSH9YI85
h4ftXwmVpwxpvDBDHK+WV5hJB9/7yXzO1rfjQZoRYAkDoP1IiNCwuHOW2rsQih9pu9lq8pVo74jt
H57oUmbT90kyqr3Rs9rtTofOLxaaJ6LGiEzcyQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432)
`pragma protect data_block
sDpKAcOHY4L94t7LfSDHshw3fCKo16vSwo/K/qaUuO1OG6rab49ftvRyKBdK63jlUQzJNnlYCX92
vtSgAQjisTpdvthYUpkWpxYIAwsA/kj2vCM66CfRPTSMCiu7MiGR2roZoGdLFJqdgDpHrttUp3R2
iCwUvcY2yfMh/JwrjnTQ9V+VRuFXHRDCECfd5GlPKxjDr3Oo7RaGkrITEiJ8HKmeRRg/0n1hmdQ9
bAhVptA86x+Ku0PcFhdHCP3YS9oKtbUVJ8p3Kg3N2FVjFPbkN9yE7otG/W2tqJTMRznvZEoFvs6D
4mB0NDZVnEw3Md58zwpZvwUKY8YSkJVuVc4lTDwBmJG2WOlHNgLA1XMLu7BOJMKu5k9O89amWjdC
vxMxJ6GcYt3s6vdna/Ulm/jLdU/COSeRGP0+sRFAEXiV2Dm7yUahbNlzX3Y9ntqWH8zBZYLeYRkd
yY0rCHate8mEu1hRI8mLQxSqMyJREnVz6AqMAqux2CcNjQXPn0E9+eX8M48TsSsbsBEQtQiEI6ip
+ghQM3Qbduk76V56VJs4k4x5mYY0F4lShdG4jU32YleK
`pragma protect end_protected
