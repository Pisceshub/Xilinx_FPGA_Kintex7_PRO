`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9712)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NyKEG4GrBklyv9bfG2Mro5OaKdYHhqxWoa0
t6DivGOn6r0xxgiHDSmb6hMZuG6355NgFRaSx83IKAL0YY8m3frBMBxHGpd7Es37k9cM5w9LbLpX
ffGY4zbm8hQpsW3xpG+E32eZXP88eV5cYBu26VoRjvMjtYOfmBGQ3WXOhdwvQ428PvPOVvSgj3MY
zELpk67Ar2roMHJhORbA9HFuV823ucKAe8BXUJMparq74lvLr/dnIoifLZ8dhcixewf0R98pBJL5
6cF9weCHiU6cHjZURCKpYtj6eQmR1j1sivtaMsf+zDp86ZwtKpeIp76ztbojkQcAWMjJu7KY4hq1
voCaibmMgqtnvAQob6xYUj4aX3jrgMMQRqwK1zmXJ629WgcgUmPaBECQYfDnsLDbgrMLqw86p39V
7RyEN1up83/G3XG/n1HjBUhfR8SIWR+H3nr/pDDCaHQKLKE1+mZG9dZAysVARalYBcu0SZeXjH0t
DsMQaj0ArUe3FXSYl1NmehqHUiX/Abi7B+nbYekyFVm2M2qJUcKmuSTzBHFw8errLzJro0+nZmCq
Sc5OtAgqwKFem9JxoEJEC+S7QGyx07GXTk5EMK0P5CaAF3pB1qukNLvG4KIGZPAbxDbsde2JU6gb
VQb9+a98cw3N4ZWNpTV0d+zYpc5kxR93MhgWlVQxDybRP9rluOTfG/pqRvlhBWn0TK1sGSDa1r+i
pZ1XT7GqffEDhKLbbmBIzKVc9pzt6s4+ks+Q/nmb7zEUolRZugNedfBLJpsiBGPBd0kpJvSimL7K
Ky8MWeF15RmBEk+VdBlI6qgww3oOD6ge/oVXnqcZX8P+au78Dk0Yhcn3+sIt4qPNcxOm7ERiXC+Z
OftOrHEtl28KsFHs+9NMT8I7UeBEzu8aGg/F1g9fJy0a8ITPh2DDKfneNpUrBCAxECDwK11pcglq
BZ0+ucgacEQrjpyZsWkGQbgkKBaMuSK17fnCyHjdTMXIosXm7NrLjVcYXu0Tr9ZukylXkr/vgPSv
GOlCi49QMNkbGEUFlNyzEFTKKTuBKbBTfwXzSb87mWVB9+SW0UCaq9O7uqyjy3DPUy4NF6ycNpbe
biQzzb7xOP9UPosxkh+3KxgyrwR4fGAEhkBfzTFy6Co0/oNtS8bJ2PI37ToOA7Um5xbpsiC/6pgw
jy2s64AU2HUCOMNMXsTseOtbcGZ1/1lp+T+aTUvrKKjBAB/hdIQLM8jodFVrGZTeNuMK/kzk3D8a
hsNCWQu5Car0elDj5dSrq103ivKBkKzHG1W4qQmJ6B4HjjofGlKeY3IyTlD7+0iXC73wW/WeYdIe
T3UhhFIFdrIz2796B1MHI7iYRJsak4VJbT3l59izRD6W0e/IDYlpae64WJWSakitj6BXVbrpy80B
tM0KEno04WcJ4RNmD54NyZ/84vndIfYNcimMRYCU7YyvlqYckkfJ6jTdaf6Y2yL0yAJjt8TOAwy5
Zmyx6pUj1PLVYb0/C1LXdzHzfO3HDJP9S+/WkdPm0p96siGuR1LnOB/fccSKxyQW1TycpEQZWvli
M1WQkBiMXIfWZIMkoDEbBdQfth9eQjRaYdzcjAWW2h4e4FntmrNJOTbaFAlQ18YS9FH/QhNJRRsg
1B1/SenOLRY5WLgWzxxUSzOfx7ec51J7y//QKNdPlPPJdTUxpp/QS3bIOIzI2vhJW85DfRQhuViM
4ITQWS5qg1Rr8Y8pGe0TZeIzlIBcoz2kVpecKpKTt1lRkUrOxJnDT+vGTc5UC0IEgb/XZ6kTyT5R
WFKWO+WgpSM+hKfoOiQLv8uV7W22YT40f3GCAY2H+f2FiqZUcsaKkhDI/W/cOczhxzjN+jYa5gWc
n8WvtMvqMbr1v0yi8mppt+klOFOV3Q7UbxesjbGOasIFjHjnNUP5Z0wqMikP2oXjmuUkdRKsKTVl
XAkhR7fvQheMAZm1PFchVfYdSDlZ2RoOLlYW1UhSonUZvP9AgT2vTxyKZ1q7RCmsrEP/TWg6lZLZ
Yiwsn5qqjviD2IafdCLAjbIwbu52pK832qkJ1SSeJAbgp83x3OHf5dpcGP62ggfFDZ8vp0jpgBd9
27RgI2UhgXnnzf1xc6tbOMOFXKLbXIJZD6YuVou8gsbfYtEXD564IVW0AB+lB9Ckt25gt/gYJi8v
W74YcQpa3J91cC4WcJNMoye2U55JqV2T+IQ7fTmA11EZSSjgaGs4dpaialcUqeoYLmrLvdn25Gd6
no2MXg6QvGHzz7aBkjWuEkBZW0LucfSGpiA5rglVCs0BdY1E7299Bmjt5WfH3gzUanQDlgdxwWpC
n5DsiiUcl4TncE+pVtkdzFYTY99cZOkG4WSKuR8Ccw2LuB1p+PdksNeNHDmOe2816dYQXALRNOJs
0/0ZdGox6JDSV09n+BFMwJu1OY0Mf5yiEFKxmxsO0vE51GCDaYOKrLYTD9qoAnGhAtTGyLBtWHhD
Vw2dMazVY8Xsk3CH4ixsCUdz0eUQbnewTM7p7yhK7JFIr9LN3L9VtV8SDxdPuvtOiBbjc52SOdOI
37BtIDnNmzsP78j6KhfkjNc+aPQSbh+9fvdcEFlXNlbNXFlLGDKXOVoe1l/a3ogYKGHcFF7h1+gc
1SU7e0maFZgz1rFO2S48UFNv5B7vZGSYTjRZqWqiekqKcJSqDOacOrv+DXlmyAtO/vOLvi02FUvC
18YsJWFTzrYA47ZXmywdQek0LVE89BmF8XbPA1YlPQlcxjWGqe+SO8pUi7c37inKRKMH0VsbxaGd
mAwWqy0eR+rn5n08dldeITmwolqc6/8n9MfcZkyDKZXouoxSx/jgfnP7+zbLMFcdsqK2CuvPwrZ2
SQ0IAJD8Xz9jvvcbpKDOaswR9nokWD4RosDFKRRcYlproEspcp+uyvBewp8A9h+Z6BulR1bB7lky
B6/CTigohbu48gI3N59OLXNp4YJOfRzYSv+i5+2wjol8Tem4jvtqBkAW2RWyZ4QieQOx/5CcU8TG
CRFIMjPMOOItKTDHleDIm47NRiHJQ4aSooMBL26GzrK9/pXlqazcXc3mewp7CmDg9HA9+PZB6ZcF
F8bECZBT7umM6CanIuvPwf5iJtdvgI7YLshLmf3bUI2en1uNc668fmeocLHXRPUQ5qUYfh7HKbHJ
EEffqX9flYglkkoM2PBekIGpqud+7pr/0PzYOcbW7otjHtM4sWK1XP35mvRz7DpCYYyk/5lwFWEM
Jlx94rp62ZKoc7Emz5CJLJnLV/RCAVfmOOHRmsx7a4W5NTYw1VqEEkZtkixCrTKRWb6a7s69CpHX
TzxNb56UPTtmCXH+QonhzOEfCcy4i/zJbcgptttI5BKDJfAac23cl4xcLjD9qKPKCQxeUm6Di3o6
0oibpcQHKUYs/jztAzWuot7tS6poHuW2gxlcbZtF7VVLz9KbxaiJCpBR+MiCcgrW7Cbdxm1xXLkx
qQC9QSZfEJ2m0Spt1EKTX3cMXa29WKg6lAmHhs6CqbMaZoDtdeAjitaSUb791uOE7SWp6MnZpenK
cu7a+97bSl9hyaAv4LeKavz0NNyYTc2N9r3YsiVhuXY7ZjsWs3o5cxggxLlUcDtSqg+R9bJzChvu
GxngChYScjFgo4/3tq3/liDDqCJon4h7Q2Ffs2sIFigThqVA7BGsA+Slwr2zjBgAZlf03oX7CaEs
eCVCv1LLmrbM6BZivQUuqJAd0FopKnK+MS65hqn9AcOlrJGpCfm/OeT89S/6yqG11evtTEiiBreL
pHcl+CG7gksar8g+/aQzv4hp3yGUtUR+r+yXuXT1E/i7WpH2ypRhu0GPUj8u5B5Rz7AbMol1V8ho
8EGe8L12/lPBRqyKdyia03ndzw2zJhyVUWHDuQhP+gTnipjzQyqoMLTjWaeGJZQvnvbqH2DzMf/3
wq0/2zVVRObl/z6lEKpFRIUUafTo/EfKsIMbcggIDshdRfCODoWvqeWxXn8wzceXFZ57iV3AejgO
G+rpA61jJs38qsUjxpgFTJ46elK/vAkeYLLuap/a7q+vh3KhLds5YyvoU+o3Z3sh3cVK6TSVAgAC
17H/C1a1H7OsnA5XyVkuejTA3xadU1DLuxOrBsnMFTrEXuKGHMbBPF+J2Z5TzFCuyr7d3J0Xv1f1
uFD6YqQmDM4PEheFKO+JlDmmQyiZtcC7kXUUcBrHj7gIzezKjwLBStgSnqL0emkv4yrTHWTeFn8N
W8P09l/apapPbA3KWNIozbipHBkzlBRo/gHEbMfWLuAWPH1uC/68cfJkA55PYyfsNHQKFY3DqwZY
jTT9MRDwD1m6yY2DDVuloV4YAc3caXFfo7oEL9fziG1SyNWfnKN/tHt2VrlwU5cV1OmIGtoF+0OV
L5JRYBPG0A3V/C/xLdBNBjDWjph+eTFFSC0LG+RHGC75/bA/rlIguHXOFmgNjTRM0q5iwQ0MVGhu
NaMAAIJ0NLrFvrTiYBmVccAvZ+TDTyVUjKBBAdw5ahWIi/vyk7k4WJmangX8qfUZMJFkf3NwOxby
QCppMZnEJ1Pz/Qo6vH+iKTkpbwBpAS13oH3PCIGkyxnmnwC8tPyLhzBqVngmVT5DnymU3wtVr4Sy
w3MucVBM81hY+5kgRqf7UulWOQPEfLBdwCD/kJQHmSw5FKRUuTdA9M66ACriJOHNphT21dGHSTcE
H4ZqOmKpGaTzkn6hPoYsasbq3aWGcusQR1Gd+8ubSKSN0W0OVm1resRE1vyafw3chsdc1z5l3pqo
rXElWypEJIYVM8GNYXMb8evYMJVo7XMlHKon/fDzbBfXrt3X6VJgGYgb8SvhMOrlJlgE1iNX1RT1
MNRLjBjEYVU/RKjqOBNc5nW39pByjJH3NZ6xvE8jH32YgfJXGB0KqMKJw9gGRXD41LR3VJyVS99w
v42W0XiK+7muHiJYXDlDX/dYmHufbPKdSYBAcNdGqpmPOKSMvFVS/qZ5TGEpSjLxHEYHoa7/6W/1
Hz4we+YQE2hI3tDVJQ1f+4DKg1TifVETOjahkND4gIkZr6peUW6J8JWko35yDMe0WjA3DPMwFwl+
/XSrQenWgVcuaAVMjP9/d8lLiEj9SDQoqgsT4FgtMFxIj+CsWlfhXzSXEb1ov6pRYbH4F8hodPG4
SZbJIckcdgxl1kkp6xwxr4SW2pMlOJdnrEjln0aRUwRAtGA6bEYoXz9jAFKsQCfo0Gi/FWLfVJ1I
m1sW2FiVx5qHhCqx1/EM8s4CkHEEa8/dQFIyOUg3sfYv7SWTTe6V59afQeqo86ZpPC5Z+PB/Gh0c
hTpixVrp4ZbxRBzA8yFurmxoCtxkaTB0XzNLPU0p8sdlJ+Axf0sxh6JoyDsZh+RLTAjvg9X/M+K7
p66e4SX079DWnVIZQS7wthtPFbEvJFmG6w0cBWLi5sBS6GiZbQcjMJdjC6vB8oQLqiNduyN7EQd7
IDOdYs3UrjPiKLBoDL3NkyiM6PrCwIGH6pMxE2nVkyHzuJzb7nyR3RhQFfS9zS3O8plNtGX2G2KX
EwlyoCOgl5lRQ2xdupl4cpyzL4Q3I8bZ+nfv3ItXOzsvger2KvlFeVA6OEB8eTvFjDsLExtzQkdw
SYsRT3RY54/CICi5p2dMcrIlyMDNKKqfCR6k8+GpdnFDnV4VcZI665Z4RyGCIsXeefwC6yWf/6yb
S9+Kp3kZxSTD5Z91V8kVA9hfUOfz4/q/pHEIuEOuSReSq/nO2AKf7FV9xkRN4yrJAvoM8rbzglLG
3MAItVSMEHv/Vb+4ANn7FwLpL+x0u35FefWgbltnU3kcmmdurNOJ/x9pn/AiEoaOq3/c4SF2HPNu
0+XFt4SWneV5rrJuDdEeZ4hAhcCrU8WgWhHccICGcHTQgLZhPTEy2HMWjflrzZ9iEuSklLXy6Yqd
0geQykgZFNhYD+C32kjSddX59CqktJ4/mFW5YyFxNz68o83DXXUtwEq/CKEoMqWRvyjPFOmqL70Z
20C7ZtC4zv7BrYreaI2rYwyM7WK6CKdRTPIS/ejE/hZ38R2b6TECnRKKxCUNoQ1TnnWciRGEIlnP
z4RFdJie5HCrj0roiHervV+WhMd+jszVqt1IeLQHSVrGg1GTBjFkbii5+75ckuGvML3scLUt455/
NJV2GhW13VWB+PB8cRtcqgGqWckFYPjeTkVZUAXauNOM/Cvod1WyEp7+mdrJW4D6Yn1VVbV4o0OM
j8SuWdVpchWG1IyKG6gdoRKZNPWh8mcQZCFzdW3QmH900V9oLXQE2yDAE3J99FRr9GpsecxxXWBb
fjP8x5VY53UwC7P+XXkILrr7RrKjFKxT43bwEBLcpHc54x7EMUPUUgoQb+Ijxs5QpsqMbQjcrEbh
l2q7BWYTPQVkz3MTAfETLcEUa9xCmpcsUCeElUwrHdYZjDLFLJAc8jh0bckp7mos5imEnzXXGl5H
dZD+HsBzebQUFxIsknjqDc1Ftq2wt+fNBLpEJ3WoNvbK+JOxc7urSqx36BfrHj+5H1hwN92ha2Tr
07xxfQJ/CZ1YJQc2LYs29Tzvp7vyOvwu56Z6TO3VX+C+OyENXeYKU1lx76HHWG39co8A/nga4HcB
ah5axkVeHKCF9e12yaYNoAFbBMs/knxmwU+NbjKUy4wm7HRsuf/fLXAwvXanD93L9BR1iNQWzg5i
EFwm+Pz9sGp/O3E/b2C2RQ5jEweHCONnHp+gMdZKq6UCitRFhhhyZIeGn2iR1kXktlhMlZekP7DN
flWGCDCV5lBC11S2+24+6VTWyyAKkUnbxXEeTRSEf3s+Ae7qE4Cnv213hvWNOhLcoICjMwGYiKWG
5vBgU417/xWbIj4/0r6K2V7+zTxGuSG0Z+4uL9+CzE4yqy6kzQiv8nZVwcGoby2uADdyucx2B5xX
m7ce4UpHwzD+Bk9YDxqpkuEqRhzIS3rGXUbZ5D2jKTI4qzeHwUlYg4hnEsKEuu3rkQacmtX2IrtU
ENepGIniiIrwekCkJyvoI7mM76CQ1h9rkYJrDxZinoRnvBlB+6mccnqq/tuEOZh0uBNbu/1aKBYu
UZL++kE3hpP2gG6mR2lU7jjoJGfR48td5IqR7d3+v1Z2JncJDuy+HvGTT9MzF/oWZeyfjBI+UGGX
cF/VgAFox6qemI5dyjlq8Ekpq3iEynv4T5KQxFQ0w0jELxGFQqePHbzolZQvYCnSgehP+sKE6mrc
oZTJqFUyq9ftDihUol+OjnFtFXU7NLobNLsu2cOQqL+S3aIFH1sWJB6AMtpy4sFStmzbZMYy6A4j
bnkCMhN7X5FT62en+NbDfoCk+viLIXPhtGxF7qZ4oFWu+UkNONb/RAjpJXZ71BxrmEhvOb3c91q7
YXgdTl1FIhrT4TBzwVSXmaq44WqWvZ6ZZ0553RtITd7nlxG1zDXZm5CwnawhTBLKpT5yHn5UbnAz
TgSmqjDcs+TIPwbhdFtCHPiUuXgKJ9ZojLbvBq6wAB0qVdYUprFYPOlX1ybPrhLa7z5KK6BivV2M
UCFVSPxbzs+RvDqW+ZAmJM4jMxv4NzAqONNg0V7k8N/Khou6J87Be/QAyhaMUJaJziXfg/pgLVSe
37q+2AfSZUVpwoJ0xjSEcHsCGt9vNQiDnrvIwmlR1h8LueXmH0zh6g5lMpDsiBSjefF16wndWwlO
FIXP2vAEIbmNFb6svPFZH0bSY2mZzEAmfebwEGVydikIBNG4c9NJ0H/RitSUAKZHak2ywiXshFYX
J4K/gcle3iTl0zPwc7uoDNsmxzgIXEvx2Zz4E4EbWhlVs0HnVwPRif7cwohfX4ePzNNgaO+Z4eDF
zKinTJ8bwPya6Hjgm2MBMHeaEIQaWcu/bWRAGhpaGllPt7HJWrrgErKY84e5c1eQCBKYAsKzrm9m
+GVT42Jk9UMzjOLtZOgdC5qhpqrcWMJaxuae1GbWE5B36smQTZxCnol7i1TNHAn2Nc4ke4ys4NuK
clz/PUFmvRGbbStlGJ+nTvhnLyA/XwZU8r++f4cBRlWvgrwDSRCZ8KEfe5hX3+z1E+L9bJKEoyjq
wjNNlMRVs+kds7cgo5BtDAhRuPKpLVW997Zt03tgLbneVc6oJHYVy5lOziXI4lyR/wH93m0xrx0h
E0jyIpGcJc3Q9ktuzhh2R5Q4bQmXVEd3S/xUq1+3MOcYnU4wnIQhplOhpJZyIAz2/OH0oy5e7NpV
qyNLDyog80vQkOtaNj0yqqZUp0lG3lxj9Hspd53R7WTH2IYh2+lH0boiOtKJpuqp8hRLQgm2qwFM
Xh8jMwL/Imua1pMQK1nveL3+igiU7T7yXxx1/AIPD+JKtGa3yXW/tjc9qsm8V/bfFv4xAnEWXewB
frPX6W+lib1+0SpDhs01tzixQPqBZQypv9bg1FkAkzcW4tpGk35rfd4sFsqUYxvSrYniapZhwwYm
TsY44fW423PWQ1mDpSzNYw6qIG2zeaxlRYy0KLvLFeQpQgoByfBOe3kncrN5BGY8OhNZUwNwQRQ2
47l0krMt3JcvmEF2UOOMyqP9T4ZSrGo5tvpWYcHwz4pumv5JtZcz5vyzXWBKRDDM57dk99F3yt3s
e3Xi13Am+/2poSlp4sM1CHx5hauvLM+8c0f/Mrfc8Pp7KiDjqVz4Y4rENoK0gdEu/HqPSY5ZT75H
GQRGq/BxYw4h8BckI3Gko8BVqQXfC1bZYZAhw7v5EfSnfrmYYE4To85xPNBkaH+lk9O94ivACDMS
0HMGEABoyl0u5c2ONICH1NfGEzTwqlMrSzxfQQ+VIHVp1w/5+XBuzCdWGXPltls/Pl4rIJvhtqal
Lq8gboYP1NUifCg4JfNIQhyY+Q5gMCfQ0HWehL+zIqutWVtyXYOSkiTgBR66pd9zWP7Z9VT7TvIy
o3ib+tvW5FbR3mvVWvMo8InNVKqohpLyMFDmc8OqNxJOekL7zy4WtM7jCz6Hw/ZruPo2/Q5XNKxr
F2tsPjQJ4ISZ3FAR4r3iToZSsc1R3qGcvogeix8089EP/JFOv6cU6U8IN+WT9c0ToC1+/ZbaPAPO
MXGhnGHarxawCKinjSimTy62ph50psnoMMhhyX8NoffFUgOgr/yhkIqDVYNfCARVxLtK7YY/GqqS
U7CQimyH6NdgUnbS2ffG8GskP4D0i0CAep20wQ2q1tq+OR9lqEg8v8XwjOn7uwyjlVY7wUTqjyXS
TsX9Yo28m5ZBEbliFc7BfG8qqCNJUvPOLQ1TvdJBdYo9ekzjWKdh91Fl/eTIE6WH5CDrDoq5wTzv
MEFPNFQuBKHTn3E2CtYIq7cK1GeL+ceegVeodug40DVBSUfViATmqIdHfBXE7QcnUYuBqbzmD+dL
8xTPnIPS2jM7vl1pc12JbXBUrw7pB5uJbMEyStJyDpJmS9cxlgeNP/vstsNxj70Z/ahm4wqwRMa3
yUPwXxtR5RYnz+Za1aTTFcfGHNQ+3ZGK2PVjhbrkmqVOzkG/yiYj22OIQ0NW8MrN0cDbZI4mOwM6
QCkvaXqTRvLVwVfIrD+j0UV581cHVBfSxLzrfwtq+MM/MJtEIPGBtD8Q3TIiU4Kq33P9rqYYMBQ6
rdc8DdZpHLEKcJ6ry2nreoEvVhh4Z8748Nw9pXHxGzqoiUQ+OwzV0mZNKHZZz2NPuZ+QEviMXajw
at2Y5g/sCNfKROyaICmfmb+tBMJxGaG8w3tMSItsSNihwmow7rbkxhMnkjwYmMwwrTdn8nGoqf8x
5ZRxeCvDov1hIybT4PFQVSAau067eyCF+hfhNBdjbxNftZGAxvyi9xVjuFHclu/E/BMD6tPsjatF
7hK99GemDN+i2C4U6ONyguqUSrJ4aiEeDgmcoIBolgBvis1IJrM8QDYsKq4bSDjBYx3Zpw07gFc3
/XIqROxWzYiyz6j2j4quASankx3m0W85Zx7OmXwgShzAcDOLgkD21Eslgd5z2113TAfg6y2Dic4H
/cg0tt8qecIcdx/Zqtn80bXh7Ow0tO7aoQZdR/Fzaa7/cjZPLS12+sB1iwZayBI8S65y/CsshJEy
dJrEmcKin/I9cqKUn3hFTGN2hlBxybVAouJJxzt2za1N7oSqF/MghOVMriHkSmKXQ7r50UV/QxVl
ZugARzWaztGidtsQPeaf0uIhlQ2x1mlmnL7KWY6jNk7Vz4SVcKLzUplr9C3OPu9JvwqTH+vyFGJV
B0VNba72mymhFYdWOeyLrWbvpgQVb3lacTE3HDkJ9c+vJOYAeY6JYOthRKRwcIjbubmjBZrpbvpL
UzM4vFeAYIlzMNc55fHb/SqA8MSuX1QX5ElV02pSIkAeix5lBybl+eMHyYNfnxOzjB9/OWk/pDBG
UPwQCJxKJ5bYuSSCJD9+e/YQQFtPeT7v6x9R2qQBGC/FATX7/4yLNODWlPAb3oic8OR+yXWckqDi
AnRIrjNf1YMk56dh39AmFaZo7PKAuPzaKysgYysG6J5BRbPwu0GabQWaqqZLcMBBDQIcWevnnWsJ
ijjlwznmTT599E9Unnb8Orz+69p/MJ+lr0HK6KXn7+uVzmIhsm0fKA//aHqaC6rjta3t8mwEULfu
n/il0ACV06sPQZG7E8WDrI0FsvElYbZV/rcDIRqikOTYKl5mXgHwifh32l/1rY5B9U1PZsX6fTag
fadaTZVNiwtwz5l+C6AFm8Kj/07LeFW8cOmB3RwqO1aZhxYbpk2xpg43/B6PoUlcfpqIz6uHLLT3
nROcek2kOO5PH7/l44lyj0RMM7USRboOe6xz2m+qfI8pz9167wvtkSYrwpH/KY2aQHwMqVzcUWU3
iZ1x0KY+7AqlgukyE1pLsfZ/igQUKbgNBxVZUdo1SICa06HOk0svTTsXDqkQl8wSp2raQFM6ATZK
wLtEZyOs1U04qzM7bvhFNwuSkyoxfOtGH0SY7yzBRg2JZhz200XxNCwD38ya/vO4Nv2+UUPWFg6J
rF1jXzZ6EBpBxcpZw33QjGvRgGKBJsZIOxd04sFRQQESlveAn3osWGJKzXgnnm+AExHRA0jKeft2
vPhP/+re5CtyHscexhsR4hvTsXo6vjbN+h8NyvcFtOjK/D2QD2P2a8HDLl9cemsbT+SbdPgmrVRN
xoYdj6PAwgS2g0qWMISUNQNtTMgFRGCPxJvAhiPt2W9zWKocmqsoltq/XKwlA9BWZ+hgr+DRqPXN
0JXXOX+kM6jzBOjo7PjN2iNoPwP+5tRVH7LWvcon/xhSdFTF8v6PlGTysizeMyf66GVtuXcKK48y
f8iqD6F224rGl9T2alj4Fft0GaspVkGPP99Dg9N4lLIZ8sQMpdHb9hCWxWMv+bB3mrFrRsGqyT+N
ugO16BpK+5EeFykyMgf6zSTw0789S74dif8+8BpSpOMKlhyawAOVjcr99xqQMniVI0H1UC/HAUHT
Mi1qr+nf/6ewCFHxr20GGEmNTdQXnu48arsZYD6fQMLmw/S9ECe/kl3ojhOJne2CgVxPRBa5OkGo
lBx6Gf3UooYGh5kTbJTrt8ScS3kqVKpxkDqJa1iUsdsQWuarzbc/e5RTctG0wVdma3mMbZwi8xEv
K+AFXuwHtr9gzF0XINO630KhceCNoEDjs0vOcB1krzSTqMtP+eaFz1y0JmvuGBmR9u+jsTpo/skP
4pTtLtd/lP3PvPg9REODjg3LDa3Zeij+vL79lYRtOfGlNa4w7hkMFN/GRhZOFN6xXw5Fm8Y2Ghm2
tT/6PzTgLb2Ut6JnHZxOQYpaYRqsqnN+gJFFAzHEHCsmcPhsmxHp/KzMIr1toqRmpCSyzO7ZauHA
0i0UUPePswZZDt5nXm2G/WT9b+b3QhYupSEG0XBEtQvRY/+JcNgCEbfBfSP/y8YBjinNBO8LZg/l
lPGhB7gi/oNE8uUF8pGVVMLhkgS3hnTxGOLGGbYCfFLgSxTs3FVMkiFUYhFbwLnCaDAPG0ulfhNp
fxj8i8oPXbPUncv5D7QD89pUh7OYJCsNYAaCGnKgTrNADoiYsiA9ZSg/wgJjx8NMCXgTLNZalWVk
jLMqociz0rMfJvfzGNYIXGHrp0igdC0hAU48if3gAuaa6x9VnA1JgDq3aMsLXxDF8ZLFA/+6cr/6
bqUiV1RnwFhsCHMYFK7IHg/gA21A1IAxmDyPVywsfdRs9BzN5BXvMI2aD1zfJUCX93Y7GPRBxSIK
Vr8KyO3QPem5uKwuWeuAwIunBO/Uf8ST8/33SMFzYAkoq0Lz9AvLO4k5wHxnN1wtFrzNj2kXKVWO
+Ofj5YRTfq3m8yyh4TGPFtXiV4JkJ7lT7xvngEiKWlpXgZosYkpB51qtk/B72IYxdUGDdRemHCKe
hRjYuPvuNDwDIGZUN4BqVgF3VCmuwTjgMhx16Wt6U+optbwTwHadHWQPfLs+dPq3+/Yk4KTQBsTa
eICuWxYtRDSh/JOra3XzeP1hQXQj9e1wkrN3FgQNCQHHrEeNHLO0kZzBGyQcJ7giW+VMtF6Wp96h
FrNBIHlK7Iujej2UfLf5X9WPbP6zgmdx3sNNRghLLHjfbOPAKOrWnmtvZMsZTef3r5NA2ZZzO1RE
70VO6UN5N5L4c6CXdCZlv46c6f/aYoh1LVFdgh4fSDHglcSvv06XZps3Qo4bW1Z3+pNoKpynH+MG
4/xmIOKJ2FpT95FAfyFSVz9JHTCoSrnGIqrh1uA8mMA0eV53EP+uwIgrQ/Yo/OV2XHWFK8tAwPkp
gyTSne0aNkyhfaqJSoz+Izscp1paMcXti05HwfvqQVNmCTiyH+rd985UdjjloA0u7U7CN3SkYle8
wPE181VxL06nA9k4aqmUK4poDyEILr5PA/nKSR0dgvv3J8QD8BITH0bQNvhNfxSPRZTw/7HT3AMV
8xGOGx9cGsgQX0kdcYW8qsW0T8VKX/gWhpG9qJIDr2IWl/9unPHdFWmpvtB2jXr/IYecS1TUbgAL
zfIMAI/M1nj5Wk1ouUtN+QJnmEP8gw==
`pragma protect end_protected
