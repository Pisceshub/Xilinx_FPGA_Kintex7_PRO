`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9216)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEL55eSAuGgIack1mk28EiE87iRpDqImXiVoGroOK+DVjMbWY6PRq2tNZ
hh6R4oejWnGmAwz+/MlIo7uAZHlWMcdQ3jnqpPzkskLd+Cypvs0xQcT503GD58T243HboRiUUK/r
0Yj7XpMRvmW+e49nvpBgeAn5dG0lyucwTcAC/0/d16qg7IQCBIBB6MriqlgvhAzQxDdfL78TPhmh
GdgVAw60V9BPsQOzLT2Ojv3dXdwgWnuwIIUlp8CA3QcwSVxfVfbMFnJzpkODFHiu1IF38Ul94rKf
BCGMoIDYCTbrrYg48MzZwKBJRhkLwtS8EREuhon+MbqgnlZh5NMtr3AN29FYBslXmZDDPhAPMdDE
GzmjykjRGNxU5aYr3ab347Mok3QszAT/uXCWQV09h9qwvl8X9Qd1UoK3UeB6tbxSMr9u/XgZQ5ZB
lPT5i4S4/5JVtAGXYkec+dF9F8rQ8KIViUiEDPKgrzhdTwVSXwop/qrFs25WaTwsa2utIw81QooJ
VCgaayQb23D0b8zK1GV1eYkNETxdcw5PH2DnY/ViSby7AoPkb1B0PU02Lg4+Bq6CA5irzsevYQlS
sXIkl9dgz9tQ0bknnZDXVA1KBVzLe0CAcVtE66Uw9P8W5ErGzQIbrSTQeb7q4jFUuWTsCSxCFUSA
Fnh612N/ejs2Jb+zwgPG77LciKbjxvTKT4q3sjjzz5hhUYhQ4COREKcHreRodtrO//p34vEMuSpf
sRwWgJbMF2joA7RSe9H6g+2UqggkaUyDVQ3OT6MBWM2PV5pS8hp2WZa+R7lhNBhsIL5PY2KT1hPj
TZRjB5sxu+2GwP2qxNjsAmWGVSf3RuOQrq5nM2cLwugUcrk4ffRz3jUj/6CmSY24ejhRDgxfY0FR
2IliknmQUE3heL1VyJ1HVFvmaW7yt6V0AQcHKE+6bd2oUd+XktiGOW9JTvTx0mGvAONAHZ3eaqSU
H928hzI9O21BQgFMyqbzwpR0f0/Yp4PKD+8D6J/rJ6sO+JFgawedkJf00bKJLDtnRqdPEpEGWJo2
LY36+cu7RbMfzjupC608KsdM3tpiFibmG+Nrj8d8hjW6+CwiSpNvru4P3LdNmHgCW17tO0/0xp0D
wpWgkfaVBIw2urTW/gXEh/Dor805jPJf/0ZPYjQUfuCniG3E3mVFf109shUQfsId3261SLgeEuKM
gKZ/YQ/JFXFUxqwxTx4ZJw0SKOobFLDyxOqzUkPYupF8gkUN62mDtT4RO1uaER1tcS/fXBiBo1Ej
w158htt2De1G68AVKzZUpRE4XPeG9h8xCCg41r6xo5AE5q/MIOEDjM/HIbtewP67VsBEvwTxqcdB
zCDll0u0W+CmHKa4Mc8eGJPGPUw0zhNnDSCCnn0nc9Gf8RMgJ+JFxWrPS0SdxSNw5N5/RR6nEVbP
sxla5gm7m9hOQ8Yu3+y8qOZ6jKOQDn2w7OpAeA7R6GZrm0SoXme43DYFzB/NSnw+KVN+uYDCmLH5
ZihFHbvvaa+iisznBCVCoOG3uMnnxwP6NxoKl0rYSIVH+FxDW/9+vml103pvrHPjWXemhZKkQaa7
pVZSuUdgztfJu7b6Zri4K/5sueRnsDO7Dg1GgpYc86bNgqhjkEDTwQIm8xkqBw0HktfnsAjNYPhk
I0ZHOWOGXsphVkiBc7RoPaydGsYTIVcIKeUT+pEEJpw+8Qe73QVqBGnFGf8aXZlloixpoX+7P5J5
3lRTPS55XadNnCLAwRpiBfK05CBi/9gBe66dSm02EzEy6KZ6PUacN22gMi/hLI8bqoi+J2Tb6KSt
O45YMkfUIKVBgo2fHi8Qi6IbuVXqA0OhtTtHdQWJdX93uuBnsvlSbTa2n4vEw9OOtOZmsoWV6yRI
EECcG062D0CanMYNukqDULyhWkaesliATYHXw6an1py5vnCmOa/WftZOLevqBm4pmqP1Vzf+I+AI
V5rm4aY1utIyGj/lCnhZrlz0xaVxQM8J4Sblc2GZoiN4C9+0d0ZZ3Tj3zG8VNti5JCsspjzJvvgr
DSfg22gc8swgYveE5/rLQvaip1EGT6gpb6zfZadxRBc9K0LftbSQYF0hqatQiC1cYq2tMK97yt0s
uspW51f9cLQyidd6qrNRWIcNnxJbvdS2gkusK2YU2N+U6ze64a4Z8M/ABfMDI1QBRgD6pBk/gc7x
6Y3V1JPCmhwbJC1+YZQ5meYbtshTQiACAEruiEN0k18EVMzTyuPL6COQUuSrJrD3VRibiaFWC+x3
QCHhB24LSUFEq1Z/VUaofsiRuMhTsW6Krjyn93nKK6Ya2IXTHMwCA7zI8+EYdskAi4s9/mrUOXsm
v6g5vvv/RgG+BU8v6VGRVdH1eP8RhxhgIk401sekKzq2iX0rNg5NC1159d6IUGwtiEDNeFc+WaCR
mtDhsU2tOegxoWfrAWw3AV3/sPLbdiIX2S47zubxlCXyRs0S+boeKcmqZY+Y84MRPZYSliU9CSKC
qBXEzFdRjie22Rz6Q+b40jsUsMzpxbdbZl4o7L81apS2BED22fuzojg4TNUAB2qck31h6JL/YIwe
ezoaJOcqQVlFXUjRSZntxPWHmkuRZWgcizgkIIosA8c9tHuvT9+X5lIJjx1ncPjAL74xEb7Q765U
ddIiLvStzUkw42/vP786ssRdkLmBXVFJzcckzFMRxyBgpVUgjyj3ALBGoAdq3Hgdp2wVtw89GZmr
s98NuBl5yOyZaWRDC3SnmSWFCcVnjNXed40oFUJaKSA/HxV1AJE/oOUwEdJ/75VFV+Ibuj8204pM
AzbRFVNG3vSusYQGgfi/Q+SntBu9zWMdsLREF9F+MMOHfijLYKw0lrehJN4c7/D2CYpfyjGsToX2
fTf9abqGTEO6qLnp9o5v5Gz/91L6VCTKylzTg2I1/H7fjKCvopqipJLoqO0LuW8zosUbbwxp3Adu
agoepN7iLznigFlPyCqUc44kLSotrGFzG830NU7YoNKBlf0/m1C8QLZrLbd2nkRIOjW+r39+oSMg
k/KYTi/wOu6Tjrq1gso0CQV0rrKZZ32SkE2BjsFZaC5mSSfB5CRd/czDYY4brenBcHaui0f+IMcz
/DCQZqV/MKvsypb/M7GFJr+yQ/UfmqmLPeSNXhRdIxV48gL1Kp2fYzRijCTUuLYCWS4uqfnNYfLK
ZeM1dK2q/MlMthFd64JmmZ3G9TZpuFR2IaYNZcIEDhFoUtQvjMuhoBjJfqO2i0q4L4LiK1vT1rju
EEVeqynQn+iaRYdnUfb34fJ82L+xskcqQEzaulCZ9hofljyJcmbK47cfWomU3k/YA4chonb8BgzN
5PA/tx9zg//r1a/IYSNvAUts2wM64m7r06maipz1Ofq8c2PIUh0Jb/u/d/83aOWsVxWaolsiGI+p
aSr0MjM0naIfHd3K3Q07NDhZOTvI8qw1h+GEIOLO210n+C5gb3UAgpYK//ymPMLMNBsWgdTOYWLE
HmXQe8pUs4a6+xSOWIATeOr3D5W0rumVKHIolr9CONnrBrqp9C/ngyW/WRO14L3GOD3m6i1Mj0re
KS0J95dGb7NVhDFUoEpQJ4kHBaJ+kGY9oTRsZMqEnmKjFF7cJGd1wsi8frLMiN+klgafFb2OGLw/
MA3GolIOCWdc3XF+vZ+dad3ZAIsltTGcS0FdIAq15PtbhyGlkJBryNT520J9wlWKFxClNeQgiHWL
4l1iDSgQErHb8hH68LnOcjxgydXKPE404sSTuxd9DjB+MHixx13jY6Fu9PnufxtygzdB6lNjZ9cn
G43Xjq0cFM4K3Sb3RZEmD1vSKkjf+0cUqFrWJBr0sXHEATyV1Q7IymoBwuBj5wyBRFvjO+gtnTTZ
r8qHWo14RMm2ZAfV561wQLRVB+OYldbpDzzjBsGY+W+MuuXGMeCuCow3ZWODwVKSqGmh8ltluAQa
6xTp/Dd0FIfPHSEkhlD5+LLywxUpSnWbzou56shTMv3UsgMrtnTd058zJYuZ4z6+7UqkCdNRSD08
/B/axz+8PoHuuCE2/D1kFkN1WSlX3p1GKbBeyVGWfZfsdboiMrANcl4k5m98F4hkRtdO3phnHxH9
YEyvIpqF3+PLT31HCieoghaEOsZxzQHrdP+PS9ao+UoblcB+HRF5rENTxyulS6XyXnFAJ1QevV8R
w/lQ6eFpPYjRxZpNs3rLKyEmi7V+szYseHuN05pWGwXLvjyWPjzPMqTdURmCKk8wWeA+3fwLYZXo
HeseG6idSwCotCOw4umrOc6uqyxNpuybPsdtCjaVtJsrXpezFqxM6AhJdhheTjlOlPVcLrUKY+rK
/YwH3zonwrOqvL7tU/F9DNz2Wci+pQ6NQm+4tAfKcdmmOTm0HNBHv7ZPKHCM2gpKd1FpmFGSt/ZR
RNO+HtY2GQ3d9GYedsyEWoTYo9JR2VFrciBfpEeP1JwEtQ9tycWMAkvoiPjtwmm8Z8HYFUce7R9I
znvRSamSKrL+csywS9joaAHP4b87smHYb/BfxIk5bd7QHcDt1PIDbajg/H/XoNltU9wviD8PudSh
sc6gp7eVwJq3juyL4fFzkPLLkC4CKmQiSV7jipTHzAaj/OmAjcZMsjFEFq302fR5RONAOMvhNEq6
h08YDZX6ToNhQ8ByAXt1bICc6qYSLGwYPD6eKsYE+98RouUVjg9+0gJ5fVfnmYcIKQCS53K3ueW3
sPCriLRijWMW5vDfGuoe2lMzr4JxA7kx3DcMJVv1T2jJloGgDg8mC2+UwAlLJGZU9PnxiNVm1m4j
7iXJKVu0yxFKXg5sT2Znv8UlMLtt4cx+P1b77vDW1CQOivpvbaWBxtjKtJ+7oOMA7M6qLqnFECwm
XjhQNKIxERLkMEDnDdpfT+KB1A3YtXqlzBiRpMBBkVAFooqSt2u3qChGjqDJtYNIISXcgWkzTOag
D+mNLj9y6KbhcEB1KIHX55wvjFLZloe58qlNmkMxrCVOPIXVBDhETkHKg50vNSL4S1z6vr0aHnQO
Y0UNl99/gRqGFpSxtjgixnVLLIQPYwKH7nYxqcBRJ3Gzwz9HTyMarrLwQLH/KPMAhkcBbRLWDuI/
SZMl29ZR2pOPRbWl8UrN1PwZHOMlmJK9DvbhEVaDh9I2FRx28iY3u8IMtGKBdk24tY2ZnJJ3Y8Fa
r0840eYjYqCBumzIcBtYxEXB9aHsK5EoPJx/ui0fD931/icUGajRfvdbsC7skOHQgX/OQa1f5me0
0Hf9CIh1loXLnpF6F6H0yaLYlQjDBx9mXKL5Be75xKXvosQxixcXkN1t/BEag4mkhqE3F93HeJAW
1gupVO4Fm9OdoCyC7D2tz0hFqhNxHQ1x8LXhu4hnwh1qUZLn3lLRtfpnbJ07wIag1WYx2of3H3dl
03hjYDiISksgCiydftBye/r6AUs4tP/RBuN3W+wOkFmef3iDWjsdBHngR/zX1xPz8uBoT8IyKkQf
xL61tisC7s6RQ8vzVAZh+/2oimnfUlnsxNsGSCGLsVF0WFHDVoPFrgSu78+JRAJ2uMHKSXxRQUAa
4bCenEn+j3yCBbP5NBBlqXNBtz+D34fbLLt1vsxqjLBaLozwx7HEQBF8HVbwD38KiFHudbcN7y8L
q6mWehtTugrlkfDOAB6XCHB9mvMXJDkuhXgvOUmAn3swM8gNaDQ+gtQG5jWI6vZwT+VF0hh1i6Jq
/tTSiA4WD5+44IiGrPKsj/00onTCefGHCvuQ+nuSTrKJEzpkJIxK5a5NIpOvJqbpn7VQBr9Hy9Je
5RtROJjdurFcBa40WEjaMOYi31Xf4u/UVHyLpU91jvP+gQDmol40tKzz2CFQW6vjqF2w7PSQaaSa
by1IQJsusybcIfQUh2GE4a0S57Vx61z4aDUUgYrGR3ZVrpwRt+hO5JsDLQXr2Bbho9JFdZIfxuTt
0v307Z7RbyBgpIGQNTuAm53mO0j+sGC2Fu1Hy/H8loQiT6dwsE9JGpfCqOyj6G2/c9XqVUC7O77C
Ej10TlcyB0jnSswQA7igSWdvDbMnPfBtVUxej6aM6V/X3RRiinXSthgIBAceai1IgO/1BikJho3E
DOK1DaudLPQXU8hBIpjFC8dVx4gnQ/GDT1ILmETe/F7kWA75uGsxdk6+6fHp6cOJ3iWvVEsVeOkU
lT+gmHoaqBHCAhjC0pN57BG9KJi3mdCw5G9uerBC2w9B3KtX2O9rvFgrAb/iNTR98aWnUGq1VSzO
d6+CdAuT/ag42SEVD4WclwFuhUbewe8x2ovhnfA12tz32m+AWzL5dpWoob9aI7Z7oyAza+12E2ue
hD3JC20JO0RR5b8scCguJ7vjJdQODLrVBV+Gwo+58JsgxZ7zDqH8i/pnGvwUmY/2XZiSXFQhLoZS
xFkjuRYQR7yYLgczKfHo6r+zQLit/KpReqSyfm3m6+vxOam+YCzFEh71F7PEr0H+lICSIOsXtGsO
1pqptc9psTONoQjXXy7IDsCR21BIMWt9g6T2l5Hb4xmdZHQhfqiHphEwOHouTtIt31YF+eNpjJN2
hx/1SxYuS2MTjUpuUeeiICOSfcfZpGJo1wsL1hw/R5iYvK4Qq/sT5/Klm22AdSl8nGuSm3NwANW/
n2Wcy2YwgfhUFmamCBSqtFtAGELLeQnt/OxNG+nw+eHstXdKSoAh430uZ4mQkeAxo3WRsRn03Wds
m5EksyDXXxP8NCUNLCDZQRmNNagdkocdOrt4hyrKCVIDglBCCThB4qgx2dMZA85w3rW5j3fBNfwU
wLCdxaO8ilDWCKS/XyEw5815YL1AsB6QKUi+mWx3yQeY4MK53pcwIOo1uTlGmZqp4J4M/R4FWFxp
BXBHPBI8B/lVuwtbmw+D0mXPb74/Rq2b6TcBFgYhDog8Qmsyy82oHcTtGFnbFWn7Fu9gCvbT7bpk
nFTw7OqZCNG2kBSMMZgndpUxagULSsfnCVFzuhill0JgqSq1FOYOAmM+P7lY0OX9PdWmUlQyZ4KG
8i6RIlaRZOCmj1oYucKTwZ/EI2ayLno2bHYc0CxrPupNnVZ5Jl9ju7aoR86t5BMSP5xSyHGuVh9d
S0005HR5XCwoJt8KA5k1CZ0/6sg6UswIvWMiULFeoW+vB8BVu+GzfYOTyCmmJPmP1pLeUR+oNaTM
TOrl2EE4pzCrcVEJjRaWcC1rk4eEu96muDZY4B9bfpQUMpD0W2xhg3b1ABHPYG33hNaFMsCHVw7T
VZ3mLWjrUKGSweXkjIcwutd/+4IDahwFLZQFPGZzWRwAuKgSxRU0mFDXBOMaPrYBo7KCmjw6YmwM
DHZ/FcWdcWtVCo7ntYYDVARsXNh44WRs27P6g7y6Q7yxBpATOMm/VR+BQ3Y5kRaJODf/nGKYwX6Z
zXQ+irS5TlKUr3J6Xa0EdHmY9fjmnTkvNAy5oeAWccmETxqAx/CTy5zBUued7IlYEWBrnrspj2n8
Pt47dvWnC9ZQBz/vvakBytPom3+Qw8oFskFn1Pm5dKRkaJ/Iz1zJ8apcLmHAaRrGLj4q62kH3S/V
FOx6cN7juTflZzbbgf1Bhb4TKCPXIBaG933yDw8UaaapXVoFsCnx3KV0PHag4/M/0iq1f2jdnMXV
AuPO18dk0egHHv8bqSJl/MziMYgNUUKfY/C4sw7jBRyGlTPNytGBBls26U4U+iK/HSSVYRVuvYtU
NCuWRDOt7KCXrTU1l5RTDcGYhEG4W7wueHEd1R+KdO0YEEDPpFj1fKW/jSzbNM3bKyrHnuIDKuaM
+QRjWF6MUjAZJEnseY1JDDkw9vjipRmU9RpqHAt8zyj9Fj3bwj5IRVPH6qyreE4qgy1ivvWvCmey
xTmGzf+6Go52a0k5PANaRv3qRCk8pas5zy/8jj2FFWc27BFc9AFVGMkRcRRu+Ku+eGuDpRwN9O5R
BlYDZay7SVzkv3ueAtD4/HEQJAXW5kS4+MM3Ykv7fQ5i1jeEPC555AXUwpUPBt7XPo0wnkabOsQG
Zhfdxlw0lKSKnE5BI4xaXetyG127zmEGLti6vyDyj37QPEEtShKnk/bF8r8Merl0X8xWutJyBuhv
VmrR1AZlS+XcOKIrnyRce7eVrzqO9DitEZ4PZvh+FDJqMWNGhIpBpfejO6rlNYKm2FyFd1HbUNC1
OfYn5s5Nj9rzIgbpptdmmz2akUUZEpW7azy77r1FzQDxtLkSS8u84O8ffMpi0beYtG6VQtiC09Bc
a4FegV1LxPuqX9Fl4UOk/R86OkLk/7Y+iKg09ZfWKPRCq7eG4yeGmHghIk/+SzT55Epy0ANytt8C
K7UqNd6uZZsbFYxBqJgPIn2ujtbWS51hY0gcuf4RalsvJzPmlr8X2QFKHhBKhDU30HjVLHjUVREV
QAOwmzEgn963LXFRxG7G0zfDQOtYyHEBKXYeCWlbSJRMUfFJZvxUGn5AUeRuV7poEqnUWxHrOybU
ImmKZdHTZoQffFIhzbS1Pao8Aph1eJVmgQX5gP37t4UXJ6l7Tr0Qr4GQzmgMpdebkyzJMIGzAevm
PoyqQ78ugrKJ2OEhtzxVG1Wta2GWcrBatUqNnALUEj7CnEhbvxufDBn8A0rrXkuZiyEq4w4mqL+X
Xrr7pXgSzGXJs12F4peeqJSR+h3z9PP6X/61NttHIcwSfQYUVNaPNmzc9g99qIQ8YY8/w1M7ez/K
BffG8R9dpJX2Eb6br9FsOIMpTw5Qo6KovKdkd1oV2BCz4AqZv4R1thAzSwjqxJYpNDTWAsTqMBEI
uWYlC5inpWhgl4rIelJXDDyuSC7bUGcs4cJDH/ALdaaZDwj7i6tm+DweyQQI5Jmyy4ycOeAH7fvy
9NFwqhdIcMvqYz5un9kqHVqOJtwDps5zbFVBckrI2qFE/hl1psfptaJH/qe4HSXaoM1gRkkJSrRg
PL0bq59QkE6+EF2Umt75FDiQzoZgNzx/CpjEwwX/4yEw1BnpHisKDW+QhC8C0DMcdbq0lJNxJ5ya
P/2pWC0nqUNi1BpT49y4P0cqS2lxTctClnZa2A6EvdKHefvz7FuxN0So8w2rnytjYyVSWQlbBSNL
YTSXjISjyigL5v07Ws6gBB0MyU0ejvIARoBGPY0hRondF/mm2jvRbGSl+HLyeVTzlnXOOTVr7ivv
92Vr2QpclzdoRboYVmxdK1oIgZiRxCUuSVNTiHb6/5uRgahglu40KdmH5wzygFBaIKBQSXwLsgXd
6zbIo37xIQDz/5/+OSccYOq3IObNThonkgHqaZNIwtG5NcHxQdWpuoorWdrN6JpkN5Re2hLhPf+5
2ahMBldEqYiCWXAUxXycsIWa9vNaFt2a7KabOHsqYRugTqTGafImmM3+s5eYrHACrnv9erasD8vQ
oj7nVMTNlDHoIknUPzx9PCqOMQjpb1x1ZIdfMlN1Gt1YCswKPKsrY9u49256VYCPA5a9WdxO7bPP
+tHhgzujufguZ3z9gYN6r/zAQhUgUah27PephlfTyOLvGTCw8Dago78mOcypVIfGQVLWHLdRNeQW
Cd+4YDxIb0GZs4TH30TCjHaF+BT6nlJBtCWjM0UaWXZzy2ZNNxyaQJqiCaVXmYBtThnBJuxmklt0
cmm9xhgwJ/3hQ8UQYP0rZBdOVpckOAqxdB6CNkqBWbv/RB8x1Qfku1o4TPHeX6shZ5E7hMjpMN+8
YQwU0KnpZT8tLI2RYUOHG4giZjlqhf/KQsFPSPUrfaPl4rmYyvVc2xGyahExQuChaPl6xV2anXXv
87G09ji0bFeXjfvP7BSrzgrHPXQkPUJVr2u/sny8n0a5kJXO+oVBEKXe20uiN4URin8RbdpIz3v5
ZH2mTiTsWLG07G6kF/fdXMvenXSOC9ywGYgyCEmTWNG1r+YPXqqhUosqe7XjXl56qaprC7TkHo3C
MJ/Xk4V4ojmN1oZO4xygm4QeXqaxtI/CVf/0doVW4MnYuA66hxHeSZ7BU37Y3FhxbEqfNFGA2aUD
MSn0JwAEOWY+jlUbW5VjcQoktcZm222eNk9mG/eBaPAALsH1gdZKBwtNzdlaRfM5zXiPmFkD9yyF
3L6nNDEdIlJxAHgnTiyt9OktOLyIVrJKCDDx6TD+2zsJki8k6XuJ7EQp6Tbwo8n9qzzdHLDOYFyd
OdOjaMCGJDFKYQ6IzzJrorpnojzvXa6u2vSqqoNI6C4bFmWmCtbDDWZvhxXlZ2DFT/g2c2OKhQdT
/J88EqlrBuQSeV7DeD5U2Y+MUAC+VhPXSuT8zffckIKu7yh82U9Oz0Ktbi4RFouTVaCNz6GB/XIt
8Ks+HMM3/WWqmM+GYU+F9zT06ifYCoL8B5e9NaRIVqC+1TXdEBv5i5LTLGYabfuacXa+h/KY/QWl
zBRlKrnT/tyl4YUmKVLYfXeitigwfmvZfe3Dy4i7x83q/SzpFtKMQ1zkucd8IQZXa28DHkBfIphO
3uhWCTLH8/4DB7sLKmVyUpeZn7sG14Vmta+iP2Q/9aDP40vSmmg1JGTDGezCzf9YhK1OZ+huV0y1
4Ewlq2tpn9P1oS/h8aYMo4JqcMxKlzbU+doxq8t/T4dPDMlgvGJU79dCcoKtG32yqDTmNUbMa9dX
buI74g33hNexnGqxXu/PE8OthYUXkhZqDqFb6rLmlYICT9kjFSsERJZDkiU7Uc1x7MOwqGl95qDZ
JkYGgEx8A11HlF6VS/qNkzm+d1z1RsXRznHzfLUh975HBkkTmLo7diArir4U9L+diakLK4VraYVH
qHxnXhu1g3Nr2KlfeQIRtUmfGTwxb6UKCEV3PZbss5Qx1Epx33YdyGKhrhzUqEZ55Rn8lP9JOyxi
nhi45NyZztYrON6CTL81/9sOXLvOux2BRn8uGR2v4WJrLWEHmVeBBSS6dPIAY5QMXhn13Ldea88m
aX5ZBiMKb8NEgCUpR7tv54h0c+FR2Z3WunRRQo2C+mdpqJeY0A5q3TXQkpDvGL1QD+MPNG1UOeV3
8n1ikDid9ykeX+j5uidyRln8FuK8mxE3zLRFJlxVM5knSAIg9RUWmzUelTjWSeRbTKaVRURtTfo9
w/WnvUsgC/j7jt4ptQglGKubbaeHGSrA4kxSN81EIGmhDYnHnzc3KeAncUCaoAOUhiAgAPSeJp0U
gtbxLa0ihMsdbrSlOS4Zk/4xrNZ4f+C3nqsTr2l3k1jgZZorfnLgiMp00sRr20k5dEm0oSQrGKy7
e2mBTL5UTFj/j4xCPmgIb0lZA3rvA+Gq+HpYSiqMpQJW0aDx8O+oDh0jXjr5kyYrzV2MwjGVkA7A
QWSyVzfzFeNjxjZNRhExLhmjJTI09hRQb8qJH/yL/xFzvpaXKR3OEH6GT+zqSm+jKWKYPvMI4bNs
St9xrKawd5U/p2eIk/WCCLdjz9lrjTwaDH7y/D/ug42c3450wLy2zlOPt34jpEwjvC8VqFNcZaYv
lT7RCtHzHr5uTZcnJHaAGXYJbm23OyeQkob11RlF6c3lwU6YUZ/PwRBZH6u9q+LdI7CpSAcLveng
NinP5srlgXoaIGnb75OobXBvcUPK1ZWlZePmZKJk2Y9eN2ybhmVWo8+q5jpx/ir718nxeoJ0/YAt
XONa2O2JO7wI6k1EjbOH+sv/ww1JJeAln2FX+FqNBSRDLU0iEf56W/tp9Lp6ROHQM2tfadkkLUvf
21iLXp70f9J5hzsjjNxJf35o4jQYl7ViE60EdJjFLuZNvmDAAZK2vGPZK2Huv+yvTbXhKbWSkLKe
lNs/65lLXlHjhUmx0BfusLHK+y54E6euhcBdUc5ZpPCuJ+GQenovZLknhrrarjeZChomC+l5PbGp
AP9/T0vcbsdF2w+fKQ2Saup/t252lE7xDMBVgPXzDLggtfs6PICiyKwvkMF+xcl3sZntvnrpF3fd
zbnNbe0V5yhGlGKIKg2hhhvs4s4QCCfbcRnPD3MfsYi6dR45QSaGHIHNF2FHjug9sWO8J4QyGM6q
DQ5yN4mJfHkCMromwdRUnN6u5CMWFvR4tLG+612wXpSzOCXrtNIoIu/zblg5oHk/HrYqyVEVUszq
NqyKGjzxxUei1m3BmjOejUvxr8+z9h9Mk8yVBT0rPjbxmJ3PndUksyk+aAADk7Un5kZZ8MfYcM5z
z9FBXsbzGLOh5fv7AA3PtamGTal+b3HFixuiO+ln63f663bpwmc6ey/O8uXnBfrZdi6R5rA+3ovV
5J1N6sfA1FU5y+nGggGG+/41FiTLGeWFOudCwUcmaK87Vpnw6YGrzofSIC1FAFp1f613QJP/QihQ
pqgV3cBwYb3o+GkTmrU5tV2CATox9pvpLv4k3K2ydy96U0Aeg6lR
`pragma protect end_protected
