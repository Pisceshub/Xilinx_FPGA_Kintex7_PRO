`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14480)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NwSWU5ugpImxTvhHi5qNlzviIOPaYEaBLMQ
l8d4cz6YAoAnyt2cfURe9kvzqBSYCK5LmlDxhs73VItEZPMbKlWARL8D/5suXiwLKZ4bO0/IHdyL
ZU//C2HZ6/jUbRCkExHFVKsGlH0bkEJocTA/lgw5m69WO8DCS2RjECgGyYzh68isdeKErQXV496o
+ku3gnin/njIpsqnQVgKTy8mJabbWvhikAJgoUjHah+ww39Es3z22JRTz/AJXol2HHCddXCSVONK
HsLYFCOwcBMcKhMqtmJKOZj0YZOcwbjf/nORgoNGOaGCt7GBIF6/lZwflaI/MYmWLOMWnB+k5NEj
lPH+gPb+vHEyUxf9+UOeF/Sp9n/aRPw5IjtmB2Tu4KiRZG7I0lVNha6mcQcfIPub+zjl4sOItkIo
2wss/ESkFioD18bgGOX1CUgU7yKhChJ3bTS8MLdSdHVtzQ7mPp5ReUrpeL95KYLtZsOvF0ow65D/
yRI1hJm1gr5vUw+EUdxRXuqPdJ/eZzO7OqiIQWpiEqjHwTmgCwkXni0fQLrC3aMf1S5k1fNiyPLY
B/SlnhQkw/p17SJea8YxI3W4nD4VcpIv94TgPAD5KXi6JdNaB8AKOsHPjVGqsgGaHAJcKz6gcE8k
dUzH2CZGLgANJut1ElNCwl+kKPMgVPqytMObBnowEQqNuxe9HNbCW6/E1Bmr6zKELcgTtTfw+uFw
m72M4lagn975tOnZMK4ofUC5DVf1NfyHf+NNWKP9zVs7Pgfb64MEmqiEb1cffwT1FEcyp58sKZLz
k/EDF0yzvFIqeoGrYRCDMjoo4hQ+asRdhQ7bv/FGYgYGBGEiemzMPSpf+HOPJYJ+YL42J5fJ6dJV
J+WsaCQD4we+4kTkec27Yy8rsKmbpkMk68scuNslPpK8XcALq3wIjtHPPad6XHgly5CgegsMbp7t
aTkfq/QqwIp5hHSTjpbtnIAa5uKxHrLSEjrWL4Ogw75UF2PhWG7VWI67YnFKUUEN2rh3McpzEEJ8
OzyK0T0s+tLmhDsx2TBvQRUgaL7tnYWxWSruyGac84QV2tjGXxPNmEslHlIRqA6gGdFlWkyRRhUX
RLg1cKfTbykG+P+GjWFbEj/9SteGjmqRwLf439nkpnVhGe+5MMxHb6N8z/bgIc4ndo8dbTRTF3FR
Wno3psYE9qZpqr4AbAhUDuqPB2l/cIYpkcC68StYuE9Q8Lbw6Z0gO15rni5TyoSY/gO7Hjde/VVq
eVMI0/RPFtw/w3uUa0E9TiTJL0BD5l1vVyj+da568nQQP8vtkIQxY3RglTKXQcS7LXwqUKTSPfLw
JxJQl6b4BI4mE33UWQpKLy30wWsnzVPoC20duLSqxUjU8qw/q2BED8wfZySgVAbSGUgC9fUsRwqI
RU1LpUdG1g7mih9XcsrUtlBT3JkCrkKQVSCxrx+IrWEKGcCE64HL7EOkhs5ysT9fFXNJiGvXjyjD
1J9Scgk/Rv/CIc8SoaRlaYqtkXJWgT2o1p5GFvL3/zNx5FIMPjf8SLgL5GbzvH2g7b0eIia8kRjr
FS0vgqF5GetfQP/1kWDqxF1NktYwhFfiF2GnzT1ouYftdxxLtmRST2KuNgCfhWrFhrXbby8gpvqM
TnamCd9ORQqH/p2HiqRu/7FzUQvDM9UJXKCgM1X7o91Qsw1CMqx6d3GsS14shlBCnWHhfVGTfV45
RpRfC0opUCool5dlhiqsIB3okR4g5ZbsSNZTZW9VH2baqFJfoXYviHXDofviEqAfY6dY2CDgJX4P
pnKsytnP0J1bchFUJZbO2EeXbDIkaDiSZh9GrBWkJeyR0DdIWU3G4HdR01zh2GTclXceWBM31YBw
PW/eE3nkRwPSaVANKWIkZ9lIgv93U3egMuFrop6lsktvygPNsYSZbRkQ+0HTyT0veQKdnCmnuhra
J+LYJPc29QW8uJuxxmNpD+VzYP6Dswd1mn00mwInA9FDlk7QuXi6ydwB7132uQoZ9MLDySTsLZZT
2H8MAoQxSHYKd4tmQn9Tvufnajq6i9CHoZcQ5vsAGIP/SftP9bM2tAsXzIwGqxxYPZZ2XPPiGhxQ
WyiA+MHeTQKzOEThAXIIXydiP37cOqXruBSBqukhhj+aQ+XEp/v9VoMxaKO9Hd6pLxibdX21dCdj
xPOwsY9R7oeKXG2tmZkWfzKP6qz84GqSgIx30T5slrM2U6HeLcckJjuTww2VCDR4qqQZPTdV+tUv
JQYY7yPTDMqhnCBaKJHYcDVNGvXEpoUhcDjDpeyvK9wesqv5c89NzHU6lylxtJ99xCk4SOuYm5oT
mP2kCiT0t1tk0AHDWT9FsMBpQWrgXZ1dRyVhiYF1ZgXIAu8EOmEzYWqFjSuLXsVdIK7Wg+L7yIIO
d4LjBFCJH+nFKN44HOOkkKlDcdzOu2A6m+k0i/l6+dm6ZBrb83rAgaIGbyPh5x0FGV6rHsrQ1El8
MGR/snekR56FKv+ftg8wg043mIaqekITPe3I2LAztBO3FQz2gKBYXElFsMyzdjPXIZKd3VQBkNLR
D1iXfmUKK5AiLX1vcku5Qu3xQ4U090rn49LJ2fRU18mm2lqXbLsJYXfGnTRvq75fZ46TwQXDTrQG
4I8WcNSZydFSgQS5go9TUbXNYjO3QjxWh7EL4BXrt5IXvb2f3TujsbY2jE33KeVf4scB4IMzDNcL
HzY1T8KSWkBBHCbwxDSy72QN/lCiy8YvZNuPk+P32bJKeeiJuWbb9mavhQd5IOERkcm5QQ9+WKRJ
0D+oDsJihgvXLwmW33EQ3u0+neAey0StbhVXIfIUykac6zPwyFezEgCWI8GcpvHHCP1Dw+piObTC
EeRpCFdwAz9NX+IltDPuSMAPAMyYNwUAXQ/hrk1L8Z/NhOpuFzrif5ZBqJEFPL1bnCneSrzt4hOy
rF5qC5JlTuc/Fiup5aWkiDtEWyYv2YWmuAOHPFAtLdlG11FCEAl2ghctCPmxy1CTOHHcpszUTnNK
ar6VPgpyrv06exSE4DKcSY8WlhQ9IjfySaQBaXAZxvpeUKmBeHCxo0RnezEeuBzCOfbf4Hv0crOS
aBbA5ng+82MhfxMrMUQxtL0CP0bgHP3/z+htUOHCarde6oa6DlOBwkW25Ur36VpmGPZEjJCsUWFs
QWbR7s8nBRxT6laabirWbHnD5KTJioinbNEUqEOaLammZbMesAaaDnBaCgVT8cdpXq8ojUROiojt
PB+bq9vzYWL2NSLKxffNwjTjIG+ij+DsCBABEDGTZ1PUyKr2VdOQC5Rj68GlXmgkZI6pnbpA/Wca
2MbZUSX/XHSbcXp1a1oQE7hA06nA1rfSAyioOfck4mb8dbzKC/VRWG22ryoSrxpU7zNlzc4THUXR
StQiyWD3pUzHZhXlz+9GkKhNDYAXPTgeei9chC/MF9XhwHCqmMEFNIIuw7upM7mYAmABASu/kU2W
+SlBgqb8O/bT1rJ9eJi2OVYLiHRm/3l8ddbSZMk9ZAwCohgVmICK9+c/RdrISs/d38K5YHzTelvc
eqs3bjCSJjb3xPBYdp0d8B3G1rhUGzcjdcUx6e0Pvjt+46p9WQnmXV8X6kKanQcry2NHUtJE2fK3
Ip4gJdDM/HxEGHB7fa73B1qEPveMuuv7E0fJVEc3hrocpo3Vb0mXRCsLhRAbbn1k7sb7tEXEYKa8
HHA9AlT94NnW4OUJvHBOXhhoAdA871Zab1nvV4R9fc0skQWsxozm9SGp33zsvUPTndqYI96Vb5N+
oLLMRaPfoA5NtaJENKVCyRfeADXLZO0e9qT3jJGV3B6Ip8y0jJuoUxJSmCRGJfwVyH9ndsRRHSA3
kJL2uflOsNOZm8JaDz7v/24cj5RROpuMkL/2DdYnNhNaf9Q1BfDiumfHoVBxWEZXwun83kJyXGDm
R1LWhCjg0ClbrQHtfFP1FlD7XxAMaQ/VkuXYz2vwrWQDg+2uZXtknYNDIEiGQGPyp6UOnt0AE2Uy
NfTrumjUPibbNHaTTQxvJzi1Y8CvnZy7LfnSnecAEF7FdLY1gilOnJdddX/EbW9Gwi46h4oDkMQM
hL1lb0Zv369F0TxgIocTlzw3VaeltA1UhTrqaxQNacqdQ8K7+dbG43ECilQt15aOeus7OF8+uLx2
wYBa3v88KwY4lSHtEa4rObb8Hp9od7VxrxkNyS3kxwr2oJpTQIi8IfHFyIXiZ04Ll70bbzcNjTU2
M61p+YxXGzRj3fr+MW9NJJ+zRENVa1tzqhO5NlVpuaFjSrO9hXgs6aLFehV2L3xalOIfVmEMHfzC
EMmc72pJePcRO/EkxawuGQc+u1fX0vYMHPnNsR+iNIKZh1Pijta2CSstksOTYE5jKsPDQi8V62WV
PSAfCRmVaHXhDqmViEe3UAaY9JXFxZzhRvCD+CAS6GsXEPCEojXC3v0i2ArP+Q4tl+PGGcGEi3fr
DjSSACTcoYYyFhNAxue/9HagbqWVFNHqDd9fyQAcqQ2mseERH2+HtQxhV3UeLolpAcK2n21OJttb
84C0zwQZYkaHW8we1Epw/JCyssEM0THmrX2k5eH81WkKd4zVzVl6ubMcgegcvdgnLJ8lOXYGHEUI
K1q5HrHfN/FnBUhDplAjYJblGGj89sMnAI6b6Bht3rBZgaozUwUNJfKlViwWsc5XtRmUiARBDTpm
TUXla97rdufJp0WMSoalH63z7Xecb81ojGO3zCDKigfxX470LM9DcvbolC/6D8NC/w5r/bSr3hlF
r3NwcnsDagBmFRxL4qc9Iv1VbsHUq8INausXuaElkJlDOk7GvcMHrm5WSaVhwkmqIUSizJ3Q7IhD
UElMXAWgOiBl0YK7RniRncrQy2BXGrdRYO1u1sFcLpGPKqPvjyhHx7SA9IkAfkgCEyDLrt0vBjfH
XDuBvNwrM2TcmXAp9HkEtrgrxdHzDN3N6Z2YukA/CrFfBuq3IqHPQzAEQ0FifDvGb0f9HqmgdOJI
gMp4A8Cr0lw1fXsIbp8DWFN6RE6AJXy3v5ys5C37oWSIZaXIA5qgn/O/2RdbAZInodnerMFPwb8E
Z+X+iOdb7qa7jAqFNcSsHjZV2vtbQp5SeoTkTRJvI8q5hsJSksZOkEhHJc9joUcI8CPitXUfWK+w
miIVpN/jTvgPig6RTQjmTMRiG57Qv3kn0LEvD8k2NcQhzJ8LIN3nZBgBAqNGZCpW+yfwprV94iAa
UTvqbacfXWjKYnLp4ziosJxlGY4EahV/vbaGBAPykGTGr4QsdsQHFt3o8npwj2d7aWgjs/W3aNqk
ZA0lY7h35yaY3swTRh9CHF9iIoiGU9o4SW9+ZLIE9/yHxnsfu4fjXvL+7HlIog/Oa9ijiEMPUnID
Xt9lzF7JzS+lZnO3T/QZdAeEApTlhVIB7uDDi9+kK+SNJHLT7bVKSrfpK+vWkzLFtHy2nZebmSam
mrwP3bljDhR8UQox5+MrTmPbjmX9119dxIN/dTXLt7cyhG34iEwK6eMup7xyXfUZ4etk82of1ZLC
PkJa3droI5fflHaorDO1IlI5mgJRkeYThcIjStSOFxNSdIskqlCLiYRYNokvBlqoSRDY4GTll8+P
X0M9NaRNUm5hi566wkD3aUgB3FBmTw9MCAL1GptKDFZUaVowMrHndCmJ6zaHIYLOhKr9x+QjDJnG
ir+RiKZkQSu51ZLnIQ7MphRVZAbMU1SAeKuFgAseENFgx01ZULGQ4WOIbgAbTQfH4/fvyC32soxI
6cCjEEEsYuiJ4TtibGNeZgDqZmND8rriB57pfmOeXbtfcXSezi2xVOxQFFwsxZOyBF7O8MoC69KP
iiNnaYzMX9xH2zbxidR99XbzRNkmo1c0HtIHvPusNO6YEqwGYrjPBXVAbNmfSjvWhcUEYd8HPFjL
5tqSobtMfWJKue2PtfBfMa3Sx+Tb0qxbj8Y+Poxz/tnT+mBxeinRYz1fgY68H87eVsOmHRHZvLb2
hKm5RG5KNDgx37gQiPGk+xz7qPFxY14WzIiLbr9eb3EM92HbwkH7PBJGDGXSVGIvrTjRkmKJnJkb
qxT3qkstZTB/ZWsIxoZ8cPgas4h30pvFg4ssfVjxHjCb1qJWf0i82S6GLuoop0yNPSosuAiT6CyZ
wocqUwW/e6kZ6wBzN0w3GLuWJHKYMqxpi7oV0K6LIyiI9p8h8ZLSgTDIa9c/hDUAuSCsJgAKicWq
Lc1gOcIlL74ZM/D7YdWSnLHeIRdrId7vyCnVMWDcxK08qTavJtSWUbiy+ozVnrmnOkdcY2cJo+81
3kKYM+/O1jpewfRbxy+8+2xVOFo2jb3YSO/tLD5NlsykPFE0IIK/UqVk9RpMkhonogv2Om3Zx9TJ
6eWqrphARTRyEP69WPzEovz7rM+FHrP/FEoWOd9ihP4+0A/TZILZh67pTZ/IhKjw2vVlwgrN+0ZD
60MxpfQNHJUk65/zPr377Kp8B/Yu7oSMdToQP6HeSVCp/MK8QosVXtMXAgr9TH0UtiWavb66krI1
cm9SGxIow23JA/iMfwPAh9ngfhPlme28qPkjOKQ0AL+vbh239oviRhWbntz95zfxSAV9m1AO/SOB
I5xA7MFymrm666Y/wGPj48K9x9sHUcrL+dA06jdOOfBg2f7rgvlhPtObxqd30wHsrHRotGZylLBx
+v6WXq+mhbFqqxjaV6UtqwC7dSDoK8dAvekVEWUAHrK3Zl3PqURPK+Vtb328FSj0hCY26mVuMsTd
cuiGVLcr2pwZ3+7dqvY7U/UAvuxM5SxJoQc4JrRfECVXtE++pnT0kuWrrdV0P32bP/BgZE9LfxCb
M2rIOt7iRCGOsIMNztlgf+dhBMPSB0REBetLl0+fOgcckkwtzSUq7Jw0uPOwYct/9m0Lg16H8687
XsW0aq1AnrUDWhsRAwEcFKhCUGLB/s0wAaXzo8FJP2DT9Y9+b4ulo6GoD7/wmgsDTGwKNzxgurm2
y5AQI7gUJBjz54qKemauvSPdzFZcUxucFuabLKuHTIzYjVnHTRjB9EAMilFibwAoIP0QxBrPpIZ3
QL6HrpNC8CZWQNNffaxKLGwiD8MKADqL5yDO0JAbHP5gi1y4fu56DNbdmAgSXzyWAgTgMHhqgyzG
p2Ftz54IML7OIPCUFAMLgw9Ke6zGC0PBzSpOfZL18Rksu/+vmAlnZdtKJ5EJ0Kv1RbCRNhZd5cp9
mW4VJfRCzca/rIzQPZGHUCrhpW67dRwfMYd+p7MShKNNCgaizfJHOJVhrDmMp34Mad4Aq3/ALQlC
4x3QMwVrgvlnW02P3kyfvq4W94O6uZDXU+B3KOHkoYAInekaGnq09Qi8104m1Tz6XWk9QrsU/Ery
5NeE+5HyMhretTKkse2l6Z/WeAEiEvFqkOkdUFxov/iOLldU9rjOyHzf6W5JYKTs2boJzHDCdiDX
QVrMIBiXZAt85mUD24znyPVX418RKwTvqgIo/BPcq3kEC7myRTBeX+uOFMzl1BjcOAgRGPEWSpK9
wNrK8EhpkLb1+SInT4gh8pqp1X4Uducb59a9sSOKpSVOzUHfrodayVGSbE6VIn82TCD6AjhPxQEk
b1QVGRr4jENlbehbV4kRVKcEA9i3ccxmTy0PR/b2Jntq4cMBl6lGx3cw9XTMi3WiE5x4E9SmHD49
BTpo18UZdtac3fxlqFUeDF+2SLJ1v7TU6O2MUUCjor5zc3I2WT6QkrUafiHXJJ1UiJhNNfCImA8p
BK7RpObxFMthe5x/fWOjxgGEmdPzKBZBHm77Cq+ep6nIGXecYc8hZC7+UoAiVCQe1g66DvxPtMU6
5AHXANTaPBv+ims49NUs/74pCoSWiCssoQhsRiEP6xEdoCmUb1BrDqJQFZuhT2j2Kt3HYf6X2x2U
N7wg9OTp4OBO3hJ12GtjvNwOYUSnN+fc0mLnanNDXQtLZyCVBHXMdopLn44Kn52cvQlnV1+dmPUK
dMI+mGNXPMVgSDDDbQ4oFlHBqowkfJ+bhkOp978S0qEAD1wtvVtEZCaixcx6opPZIjbOyMY8e3Tn
koNzxFpXTvbzb1pz1BaPItEUqwNG+OHXMOAnXNNxkJvGBu1Ot8rI9ubwBRVlLaa5UbKSrLgCYNuA
alDD7gE/aY/uErnw+Cz2rQvmJBEc3ih7S5qHoZ5hkZASRNIHul+tjR2v3vF9wCOKW5l9r/WGBsLv
7dtXb4IeJ1NzCifppQBj3s6gsg8ihHM865ph4TRLeLh1bZrUHhx4eL5kM/Top1mVreVp4AscNwAd
sgT9GM0n6I5zon2LuWVCGjKrPgSFiRooOhiKXLEhDWT2wkhYyuBK1ry+mVIktrIAp2ItJG9G1xxE
TcXgsy0YNz6P9FyqOIzKtdgsOdzeCr0tt5/h+nDd8z3/eEYBJe06asyu/wJUAMrXi4kTj9SJiFA9
yq82jjyCelY1ci11lSN9Gq1ohtwP04odLu5t9Z7VsXy6hv6XHgG2ly8JZNLRFmLtu+H9agojs4qg
53h3qJMgGmnXjKOdkmomTDV2vltmrUVoim+wt8VgZTrxbK8xN084zW4qictBMDYQc/SKa5PTSV8z
kffkzpypBqptr96rN7foNL18dmSeHs2WmJBAEReTUQFARzVldKRX15i1iC69LSxgJ3WZRSwycBcK
tiMerNENe+ao3KCwxnApAKbHEKHnrHJvpYu8jU+vyXOgQ24U4q1QhEHnkOGemaYzA99hTpNK6lWt
ynpXJCz9UhWcr0FH0KRvxzlfO4xR0whhqzhQksfuQfrf4CqKY5mosuU1hrItQeBCLoZ48cBaJBpZ
SkP5oU9KmcVXb9SMA96DBzDVH8a1Sno/W4Q3p+ppBb6IyMTB9376pWPVFAKVsGPsN8r7NyJRqqf8
b4WN557jJfInK2RiEqPKl+8GpUrmAJlDRtKSpABDuKjdeYNcovVJuGkk5RMzFqHczZhpSTbJaW8x
8oHBaL7eOeRk6ahRd7EZk+amSUZvoy6PpXG9IK0x8NwhxETsYnpJpmhozVStXBIagkn7msuhHbo/
hL0VImVrjBPmh0k3pSTFxKP6cUwU7qjjCC8GRTf9cMZKLEEBJExWuF/+gIoO2YKXqVAmV/fbecBP
StAnwAAmjRhgQECHHkoGW7k3OK3l8wA2jy0jcDlUuyy4uA0WuY6UWotqWDZGP5BeeRCDrrLm+wX6
e/6DNzQ1VqWqCUyca3Wa7VTtG1Srjy3dcgMUVO4MeTSYTCAYXRgWWRiEiPuA3h444g4B0AYb3THe
97VDGgvdUn4YUxgV+O6W2qAJfAZrTO2jsGC9tNcSwhDi2Bm8bCtC1L0gEP/HDnFvAObOnpgMpYRw
+XDawJIMcUjWwAt9SzwvIvPKgXRS9vrOeYnFCBMGYPxUr/xHCwBMa+jwH6XnOwS6KgzoCt6SqnQT
u5Vv8N/CbiiWgipCfSCvjeB+gaZxoUmImT2el6r9kkzGq0fapdNC9CGMIGFY3I3qLy1MomIwhqX4
y9AnGnVHnmhAG6K2zkqauh2gGWlkaDV3O2nuAxAyfHeh7wSvHckVkGxWGUumsEe6llA20HjMQeLE
VHZcnMnJG/NFDO4XW3ABui8GERLdca3v5gbFfg6TAE3VNa+s1cpqWUq7/YHMbksmXOG8TQlvnu4S
H+Bk0lO2zkQcoV4x8cmddv1eOMvki1aPyEm3aNsHzlz3U4FtoMoSAxfhzA8u5DY2i3Wq5QAaV8Nm
TPvyYGeuGXE276axu8j/6a/YG0nCcq8fc5RZC1FkaPlf4Zfh2cBv1BhKW2Z1V4+aoSsffbKUuRIF
ZHHmiyzCafDSv8yDMB3r3XmjFVoDpPWzndJrJ5nXu+x7376fjJsfl5Wbdr7PRxO+v3HvXtvkdPUy
RM0L7AwWkEG5hGV5N45lGhlK44MtFITixaFv5JpzJhrr9EWoCOSCbWZN7HWSGfZb37hnfBXnPCTQ
5L4+3c/gsxbEbbSZ2h8e/BcCNTKHkbhGTXlQ8d2AC5YkncfbE7JkhfO7Ct+JdLpOE5PchNTLFpYN
65a64xLRGq4ig0q7MdgBSsA75obqUq1Uz8EQoQZY2FnORp8/XSL2qv76/N2Aq06cGuWP7ZN6OnSy
kl5j6nNajTwRxOaVQjjVzFohHf5d3ayZhVCRxDzuzshmgvUCZmOSAnrsqJX/K2+SwFmCI2bdxgGW
R5uOb6ErK/ljoAKiX9CT8u524Kiwn2+dWluCsUn6zv07XjYjv6EuDEeF2EFCk7wYUVMqMl8PzEFR
K9kG/P9Vqdmmkvh4YywomCdcIa35f7L4lfSWUX70LKzngSI5UfQCWyY6gPvlEn+cAflPTh1atbfo
8eWmf9PUzIfOk2BgPhmI+eR+6zT8JgigrwBBq/ROPeCixihwBMTY/1H9bvFqXA8e472SWkUo5GPd
t9xh2ufv8pthaNMb0YEMsKgyJaw7y9A90YdFrYPCbBOC89Xx6z73Fg7y0UAlz96O0q0nUExSDHA7
dnOiWHb6hSWhAiJcjOZ+P9aW5gr/A6RRhGC2JUhqM1G2CkD+P/R4aP62Gum20CmQ1IGGIy0Kziv9
5W9MFZoyBv+JbxJRm0DwOHXM3RoSSJZnKIUPwKEVC0aKCPI5Ytagb9h6knOyXUHxs4MDjuGZcXJg
d0o8BGZM7KQqUVE5xZ9CW3F9JrVMy75gZM9+kHqzXf81DLzL+1HXV37XPBNGgV2LXUnrpg4BFVzt
2m5tkDYfptQO0ONI1FwS4BYmf1QetvO5i2YRFmYAFJMB+1Bjiaffk5AVa8FK7CuYJ6o6h4aLaZ2Z
e17jjRYlv6YtWv9cxWOhvfo4X3X3R5kRyhbu2rRozzMMOLJd2WcAAYhyOA4S5Q4/T+phTpvwxTQ7
iQUjpTvdjvNFifj4jjzKJGPYiwACMbFux363Fzj23R863gN2uKgHzyazjhZKMBo6qMy8kJUyR3bR
0enER5F3TcWmIgbxzP9oenW4Yj0UpPx835RPbQMoH+vWYaX8QrECt3/+wk2SnggWolSh4WEf74IS
c29MwbqdqlAvba6lXGTm0ES95iw25m2Q0G/boKyUJFNwfk+F165pyeHrnSoYZh/1dEcVB+N7NmiS
qfsfX0T5aQBQpOD0HnEWfHlfKlJuicQEfvV5sWSqHxizidYyyJexuBpByrkYsJbFuwituNNrU1XZ
kadBd+EydwNcEjuD8NT+w5kaZQDjfUym2vLUAboSpjD/oVUTUCX4/RzD3GMmPUrvX3XkebcvjQiu
l/QBj2WTQCsF+B5IRZZ70CGC3Q2M4tVd/f//w3uf5AE+VMiIbnlQbwJOTFEPqY2vgqWZU2qUF8aZ
LJ1H8AVklpBdXfUigMyAe3w+gBUEGXSzvjnZ2mxQO1vpGNy4DluLe2Zig9PD27uB1yhfcgsI8k1Z
y9N64pgh+2vzj1MjAc05QDy7AUluzAjCExfb7O+54nj3MyPkFXTLY0vJ9tuII3WhOj9F4tv59eEE
loeE2NXFc/d6qwNjhpLLDww7Dv0VFb80gmPtzirAGun9Kx8iYJ9bO81VuYUrLsPVYu2DVduW4ruR
y06vPeD89Uy7yusGNQhoCKRw3aTHh5m7qUu5J3B3rTbtgYmthHekhwBLaJmefI9AGYJJGTRF8zuL
+OSrLYMxxnw3Qj1H3GPltRgEL8dQpuP76dk9qfEgwCjpeDmUjVlykM4KH4XAM4K6GKhLOmIuuOC5
ntnHbaI8+HYkpW8fmr/y9D63cVMd6pqzWt1Xew0dqOOiei4pxK9m9vb3FWMjNPNOYGBtJOTtOnDU
hAVsWQFsvq2BtwxobeBDxlk6B3lgZEF2pM3NO5Z6O4gSifLTJRv1uubYhAPvsQNbNn7Sd9L2SDDd
yNsnzV7XgiBsNeWfGhQUf+GLiFW+RQY++DSq5OMDXXRbgPOx4bS5HAUBWJ5CpeXVZlsyyak50pt5
YxeX2QHwZdnSDtPE5LKnAJX4f31AlRvFMF3O+5gZBRpLqSMjH4EiZnntyGPwEpz2OJrlc0V53ASh
boBUK02qV6wL3WBJTQEpLG1ugrtLBFqEfOJQEqt9rwlFOS/rj/Ijb5J+bbT3htt2YoMgYPvOGWbX
G2i1iOCAuX7t4PuDQdBDp75iqDkxKIQWBvJjX/xf92M4kBaklB++5I6CJB4Pmw06g8NpjtiYZhuX
B1hLuIPj+S6cux9SMaGTV85cai2GLMhZ9QW+eFcQCWW7gTklYHqDnRyZQq7ON4ig/anmXkF19ZoO
8lj0n9Rlb96pAciSxS8sGuyT90pjgA0QZcb28r07ZVVgt+/YyuoxZtLGvYMq3s+hLcmB6qrLK2Aj
4seg/kmU3jmo/6mL+BnM2ydYuPbihIV/u2CM9plAhdf0rVV9sbyr/LPUEc9GEgnHXvyR45UhTgto
9cKQQ5XVNx1e7ptw8qraI+fATI6ZORyfDKXcI4ySUqo66UEaN9CnXZcFdrPi3CUoqlQwTHsLaSAc
Ejqp7vXFjNwkpAC24+bhTHbfADQ9tqj91Gjr38IwQ0S0l7KPDK0TfvwVDq3/FiimqWbDQkGBb1hR
0ju7dlDWBa0GLcfhIjqpqGjXB3BDjTP1XRjHYQzX2oIctJiED2I82cXYZ7hsLFOiRPCooC71U6jc
i2ezhCi6oC2WTzM3+Kh8RQY6C8/EkwHIjpdkJ0cVfBn1q+WSAu3RpsRl51tSRtec5YSA/M7JBXvs
mlB9p9dqw9BHBLEdBLU+sxFlMNFrSV/O7CQ393cR77XDALCH+KemzeHCAvrL8kjhmT/YQJt67I2V
1igIbHSU6fAhRGvm3hcKDWzsAPShDfHjzviWbJPxT2AOmrYjEzvBau1SprKZsSXaR4gmKcHnJWso
0WzaEuHYJUpRQLD6Or/QgZve1azZ5I3gBwFhlidk2JN50shXzK2D8IXugFUTP1lTGDrV4sZxM6n5
Ff1o/iuBaKcEbZDml8/MFRyVv6o5M88lZbKmZs0FsWOWoSNyD25EoP2qq2ivVTYGoXTf6SE02NJZ
oxfGgZjwtBbJmcev1He8MEtodJQpgEYuIwzMJaUGJ2khDkau6g6aSLaSvTwHzNPpMHdOap6qXYne
lHdG3UbqRublh+pxD0/ZWDAqazlg0ukweHqDqyhr/n0NLs/rrKpX7mNN61gMcfSGLCvWHIViqyVH
sWhuJryU0p8QqzxLefmaR1wPgEZ0iMRwhVog7CQbyLR+i8715NKpTdFMXCvBjaQdlxPOi3/NuUMX
dNfXNGVWO4AEDf2/TQZJGgMMHBazFGmy3V47il5A3oSoYNxxg1GFBnV3OK7RoM0y2SyOpHUL+JVy
p2BGWzHM0Yc37pF7JuinN28OWbjnzNuhKFenQgJT9Zp33J8o29SW1hpDO+gm0y0Td1uxh/ZKAzz/
/jiOeKelubX9hMzzA6SWJZHswLc5L5RowZ54FOsgIMEC6+cUo1+b8oRkP1S/eqWTBViszcsMl0qC
j9eQCpfHh7ISqNBUgHrSPkt+kqEwll2wNg+SLJ9Zei2YyXgCRxl6HVD/FfwNrdr+RU3WAEtd8c8H
YT23mOm9B1UW0cGLWSe+n0XCtUmYqiQN4nmid7eAD35U8oPt95JlNDvQi1+4e8fjwM8FrwVJ76gd
jd6bZoW03U/GiAtXadag8SFfXQgTDZAwodZ0CQJHAEULB5xQEu3BJBbz1K/ogomsY/KnroyD02mO
EkS4aefx5uFrAieKx+WoVytwGRbMNX1jYShCZvNaEa77vBnm6G96weLoGuALxwEbx0f4kfCoV9gg
Wnr7MQoa2kY8a8zRGemufXZ6UUZKMP2IKCLWObxLQddgKtz8ZEED8Mogwo4KG9RD3uVKwfWNt+wU
UFRiOUY3NpxYoUIvKOpsuOQLB3lmUmnt7z6s/P3oKeqbaVWqxpgM9rbuUP7IolgCWpx3Z2k+Bw+a
x1lhRfD9EV1/VdfXVjQUF4P2Ttv17h04rHKFze7esmlvSWmkXhJ9s0EDdRG3x1PnzhjN9BBTaVkM
ZB2zdwdRjc3HHX8mylKhgGgbc05Wcl04XHzrej6qvoFDFF/P8WGUFvkSAwMbjB8RMHJowhfagOdi
sSXySVggkT2oD5/cDsCXPMozFIjKBahHJXo4Q6EUeyn83ra3yi/kOPtRIDuunt+YlCYhe5RhnXbz
QfyfTuQ/dzfzOFFxRT/5Ed4BdSIwwRD/gtzfk7x8HHYhxgpxdL4GuRxmV8noNqMIZ6SlHR8oHK4u
eLL6zyXcpTIj4N/1zk0B3N5CC3Omdyph73lNTrS9ZjX0H8Z4saY4qMgxPtby9NRdOvGhA8SJ30en
YjcogzJtjiqhDn4QjL1uyY6ZuRevPs+NCJ7gtWirTeb6LxQr9+cpWwZbyAdbpgzt+8Z+D58q4DiO
UwSvbXP1hiwSZq4tRqeO3NBufE57RvUDhVnC+fRZvuA6pGyvVANS5DQutUHt1Tnss6LMH8GzyTxi
QekPhI3RqXiFZpYA0GouCtE6UR46QjyP/M2s7RPPD9QD4AYS6ykZ0IPiPfeJMwNozfZvxrtUj+FD
IFUzwfVevH0PJtc8+XchQfPKzDUuUSkRWECt9R22rcfcmUC56/DTNVSgYpagDYfyQoyCTyv6lAtz
dXrlmGBB8Wvn7pgWKXIjfg67Uo/f4UlkzsnAh1SIsNiGgvdpaVHbbejgwyzYNY/ipeQiJGit8TsK
DyRa40I7S9TImgQM8S0sBkybRpE57P0ZyJBY8GimLQFlRdwC95nFaZ/B02WIxJIYOEOlYzZpZ6xx
szhsyVLz6kiR2EG07iWEXD2Z33G3IYPpOxH3TRfDGykAf13Nv7qljT04op7bcSXIhS3DMPysk3NZ
76RsA1Cf7nH5WaaAdheCEskPvSXu3O0BOAUxH4PyHBspAwMCPkyog426/4kvlaQVxRmPMcHMfOUo
enXhX73wcNoqjTUQTveDENp+DWGTknJmFrMs8z6h/fTIfhnGpLnOJXGyHVJgaWxdCjr6xwGSm+QV
aDJL1Nw8Vg4+cA+mQIjxW+ht9Qw7jU5uzKUbCmtdo1MeiUrj/ifDubljIKOVcO4tu3Apw0isorLZ
bPrGxCSkrzW1mq8Q4JZVMM3E9Z5UL2loQOMgJvPX9sTjamOdJz6zfb39mV17SjXpt6MP4JreSwG1
7FrmXQSycwp4Xgu2KVMkTq6cRYcsV44lpbHPXr95KC3D755XCvm7D6Wkc8940nAA0SbWrq33FWez
ibVq+lPWMuJQxBuPjOHe6lX0F6PoMxxwaj3VUfR0KmP+Xlg8sPYsbtYpS27Hwc6Fb61Xk2JaFyZL
SK819qweVezxu1bk/zDdyK5tfV6c36sEBwPfhXtAsoAD7i8Phb94LGfWOCODkgF4B/z5RG8R70j/
wFCdGOMoqGroaCSGhilkisYzLftm6vqSATtIBsqqKhyUpWoBRi0Z+8x1Cjhy7L7vcVnrxtggwKCm
ifxMdphtCIDgNifgiSRWWAD0jByCt/3bMOVWlKKDEKTQdmoAozpscQBI76tsu5jvvs6Eis2/rfF/
nLEC7Js/hidJUjpLOhTP7omO7tMSfHp7R+HqgptB1AuQAvqcC+ssmlM9mdrRKmA+nPnb29T79wrB
IbLDVM2P3WYTIyvSUbFaukkbrEwTghyhleytqv2eEQeVlZMXSgLtLo5PXHXT89B4VVyJ3ctr9ZU4
EmB/1OPoLULysbZJkkYwANIOPhbD1g/GtuNy9JlpogDrJOmW/beNeVtBcy7ozot7m36onUmYSoV7
kg+NVrlyPHOEVKa5DTVL47nhXgcGe3lWwgv8FJ29KtJnUBU5j1wStJiyorFvw19nnqDUh9gbcOOy
egH8wTG7pJpRURyddsyh41I+trILhUxcC2WC8gsQkDrbU0JLaAgic2PQ+1ky9QKsFdp2QeyHjIbH
nYGxzrh/rntTu1250G8NSGB5PgiFjzNPEHlZ80LApNko8Qaal2n7lgatGFWzCTlFlgYucm5q+0L5
oaz8Opp9HpG3Q29c/8i4b6re2ot7rIYiAQYa0fS+vN+Sr7ixLPxDVES196iDhH+mnV6bKVuJhZ9a
SUbnaLkwBlOrzNOwCqHfdeiuGBg3J0E3oRkSlAjAUId2SQNOhe+abJnKT8zayaaHQt8gibOiMLN7
qEMJYjLYa1/eAjyGxrV+lA6QI5XOQq4Pt0hnCipzXW/RWYdnluRN6XVQEZJ08BPx2WyfayUAqOno
mPX9ptgBC2bcpEVZQ2DekuEPgkbamlL1FOfQjVvfqn4Sa6BMH1fFCmDYSWsY+92Y7qtCZRQ6D/iw
3k5I2fJ8OPxyh22iUfC2v6D95WPaGno579PlO3mbVbgrcmV5qLYXWZ4p9a8q/sltbAXwETOBGzcH
/ES9aHM9gCzmtmS+L92QOqH1KKBpC0pJ4l2/NNLG5L2r2jUvR6TuAHD3lId6Rl8oPnzgAYM1wRTX
8sMK4nrgvKS0AeC52w6L5jh+CHZU59ErtpNeoRNTzR4ZUWY09+1J3uYs0WI7h4NGSzMG7Rzyd1Zd
H6o3zsM6Atzvqtw5g5+gi5lPbHmOjKz71ZCgZBl5/DHZidlCKxe+155VJ5ucaNAWmuHebzwpYMMB
94QAg0jy/EYfUnKxOQKzlH9+YMpQprx7y6+gcQ034csl9gAhD3I+8HrxugMHNc8NFeaRsUmOjxwN
UF645Mj0AmqmzZxRNmQxpuOX/QeFXEylWTThUFEk0wcE/QWSIDBDcsdhG/GDKW585WXeXfaNrBvb
fXDC63GpHfknPqO0hM9Ei3chrK7wj5h43t5NV28iyd34/4INO87dlSPoY6l+q8RbBrsfDyGNHJbo
s1gheVreYRSiTCDortqKEmShkGbCFinkqW9Kb97tPnWO9MdiaLF9sYzcq5PmhnLMh4A4yDI7gjyx
yt+10K6zzk5LZaxyiAe7xvtkI3kGcTL2yKXaZT+qK8g/6ZtjbLwNEaRtZX0AAVUEjXlc2V37avMt
Aa53SOdEZcN3QuO+9ubp/Uw08cxy5fzHlM3GhmRzH6c2ON0ehi0ic5JoKn6JpzVbJViSeiv2UWvt
JhLVMlcp2FsJ9B0iWY8HqLmEr5jtLttped1s7FFUQjtdvHmlhkKlFMbsDQi8JheJtAdo/lX/xEDr
8+9fGYm7+8558iOTUMA77OAOKGSxa2WF5oDzl3MQsC9lLhhlw/CTNiJuQThxo8ayFqy8lxIlfUxo
Ef42cXXLnkAB48SljaFg+WkhIoCENQ5dkvOCQmtsU8A7/UTqRqbHJDrnOR5MGhmCqXsE6LBDbBav
A2OK9isW3Abf1zGuzCVQ1a4lcaj7pyrz6zNNxHIgycGFSljo/tICAvbV3Il2LVMcfU3DQpnKXUZJ
brZ6piGbxF/G/PE66IhT3RKDNvyGc5S0eYgWH8L2PqM8SzKsHkFghTFOobt1ma75tMpyBUVt8ZJu
V73pfD8vPfabpxx3TeKNdd32yiJnqO2MV6K/oIOkuf8BYuUXyZYgrXZ/Ttly5+I2WexpWQUBYaKW
3KCEurddLqaqbLrUEiCnFlbME9OWQWYV5/aN6SYin2OTEMa54Aj8+LebSYuEFi3aggdvMKv6YzPw
J/EZW7mTUUjJP0E/NDuCbB3TEpJOS2qw7AeIdFF8fCOByIW3or8TvofJzQ542GCK/3/A9HTb01+L
CrR6CK2wa6GMAxIur7WLUYgcg6eUTe6h2Wu4U6w2uOIMj7AR3d8wkj7VrYVZsL6izvORwgBND5lr
BXsqT8DzQdyGH9tR9+6m8M/VIX33ZrSq2zgA28FRosNoGnEKutZnmfS0Dqr5mErjAWbeYZ71lZu+
HHCp7GR5yJ+O9I1dFN00gAZmYdr3zYX7dOqwJDBUZjy62Lksjhnw45mYZcSazx7VYo3w3OiSvLqF
fOFu5RpnqGKR/ZpnkhVj+O3FSR8nHBHcBUV2u4FJJxFLfMKYpv982Xj9zqfEQ+4zjZbE7IPtz++p
vV7qv4QHUdhu6Ynv1zitpjXaGJ8lQwkXFkdzBoMqYUgmgzNYBcNPqy+rk/Fvq6r9ys3UHqy4zUTi
Q8rBGpeOU5cWU3AA6hPBxA5omkiUmB2ThNBoyuEa8TJnCwa5E4F+Xm4AAOAQ+3W2lAO9OGqM0JLt
95oa2Hf7DpJI5Of/XNOwTLv85iaCuqd7Ts0bYzfCp6HECmQrSjGPoVWQHcATWO+fe5e8TYRtfplF
zlrLgL4ufUK5SWxT/y3xpT0BoJIAewWZr950XnnZSqqvkhyGy2EoLSBF/mN6uOG6qpeP12Zvhcaz
Jqh23kF8n88YY7ecUK+aso+mPAidLGLNdDnLp7k972tuB7y9AnQnL+Yz70hIhxRnxr5f5zlfj//T
DgvqLD6rQ1WMkf2kCp+UPQ68letnxU79BqrNoxoRzTlzcW6e6Tzja+L+BDdnj268ck/HS1XSrxfD
Nw7d736CCRTXPbNxY0+yfU2GRm9UkqHqPS+EdPqjNeRXE2v0sSE6h/aj1zSkwWvdN0w5NYH5nY6a
8j2Ho2Jeyq/cE0sk+/qqx0/XV6UDz5d0R+tVhR50AcwyQ37YMn8HaUWJNPi03BI96AQk6dekRIRe
+Q4jhpte7M+uqYdLl4MI9E5KEJ9njJEny+dsvs6RN/dh6HJ+0Y7wZnjh3kO0wlBX5h+uWHoH5Xbp
Voi5FLHAaVT0JCnyEKGOP7Mln9fCaBCbOqFP73XTLxXnPUZc8rpzOd2fQ7x1NpTIDjSCvG2b3CMv
FQPYg2Wootlu/nnGxBM+LgNEns7XAkZTFGok17Gz8EarS9IS83YvGHYLc5HVDNg3GXUdbyshOoBb
9/Kd9bzE3Itm/bc2bMdnfYMtaQJBB961bqPVnqvM9qF6rS1GE6R8mKAMJ1IfEHDCTNXIxdz2TWV+
bPzDRrpmAisuadf/gXquQjj2+gJFxvU2BUwQnWQr2VwMen9FDS4TWd507/1bDlCq5UfJbuGuuq/p
2X2LEYXCGCIZ7UA/Wo6OWlm0Gwav9QsSuN8ZD1fsyAo3aeuz1F27VDhyHTADPc2cMSm+Ru6TZyhP
Zzxnb9ZKkikueFH6WWHq22de8t5t3vTSac2Xi1q4OP1KTcNBUBEUrsZEeYKvVYQ2T5UMFkXaDtkE
dlWB1LlHHGwyms4JwUJPSOdH3B+TS6vJr4yc/EcUUmPz2W2F24F/zab29g5y+UqtUr1shzqy+JxW
dVfc8jbUwzP6l/I/bSBwGqDPhyFzhC3twkb4SC8+QRz2DbH7Ue6rKwFC2FpFqEPSbfgr1bBDZofY
2R97zT3oLK0LRACTSYU8n7tAhz+t7vIcRJHbdhzoTbyGfhw6G7v8fT5DfLl8Bc7tE3ogm6NLxsaC
O9c=
`pragma protect end_protected
