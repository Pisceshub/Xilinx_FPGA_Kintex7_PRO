`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ok62VGLnH0bGsShrvDxmMQc7W88hufXDwdHESsqXG3ApRNJl4b2UGRJUXci9z7ycPJ7DEwEa5xOt
4XLP3KfoZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ChG4q8RpnjyX0Bdlu4jpiqa2qIyaEaw4p2at0f674/VEIQonbysAhpHJWYooZ1oTRlleVIwswWW/
da0RVJTzly8As+eVS/tYhb7TB/MIMJiP1oMnY1gWvviPuyX5qDkTN1GajiG0vPoOQw8SYOGJvNEi
u8nAKK1Wcw+JZOxpLQg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WX2XZsDzfmk4yEJX9VCAI1sEsTG4do56hJxTjRaIOloONJAJdmDYXYUKxlyXht6S2wTCWhPRLtPd
PNApmmizFtyWwJ3mRwIRRJo0JqkJzzjq7toK5Vt7o5oTkWNhBKiaoU2N1jlLnRlSrOfBRnbT0pbR
HvsVYfSiuf5CxmJmWkTTO2J+p2PfnmaZZugH54GX7xr0T9q+dNgJ07ltJJQ+V9vhB7U6XbTavAL4
AMVuDXKavuIcEXeBPfri6WLSi09O/6tWPLZ8Yo3dQevEorre+uK5eEiPFW9wNgOCsURAxSV1bEYO
CPx3Vd6UgkAqQpLSb19egrBqiigAryuBrJ92VA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RzFJSzX64wRgI9o8JdttGtN9IrIRkl/WJULvzKwWt87fjVa5GOllG3GxvtESknc1eFAVJN2Pk0Rg
iNuziK9Z12B5bNtoSzoCJmM9f3pSNF5LssF6jR50aO6mXaRNoLW+JgyvSnHV8xxA63Uzsli0+ilM
+vtB9n03LTungEEVt+wronwdop9zXFx+NvH0Sxu0yXF5mHC/6YoS2KRD9aApWwodOTy+RCTxQeE0
2oyQDoH+GIyQtDyI9kq4EBaxxrf7G0dBOEQaEHB9KtwPomk0vRQxC6/JsCls1qAqvk8qBQ5sIh5d
drXSN0wi/F6pzMShCPvLZ+NdK+SOqV/ZFRvYlA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SLPXyGx0HwfwkogKWGhAAc4uSd0TL2rfeXBAkpuZZtxgxStruZbLvkVx2ow8nz5xmVwM/4748Ipi
lFfBacKRNYs3VZVufbd5khTLiiraX2EBV8H4Q6l5LYh2fb1suo90vwGoiAVF+/Qrdno6mNyZz2M4
x+DT+/cXXOFS3HE6gZ9IX60N5YbADyhGlktfXMLCQoXNpY2WHL87qfVCKzJgbB8bmp3PYxI16cpJ
+pS8eWLBmldd839DCPlYKP1Il0ONl1+TRFOOAt9UQV0T42WRCimZuMZlr4hkgWmpsC3myzxioPHi
FXSBRw0ZUhjqx7B0Z+1oclU3glzUvFOi1VRksg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jgv2XhgfqZOwrqDWFXxX+cz8e6r3n6Ma0Gj1XMqAb1s/P5AiQKNLz46+xDMJfdQLd5kRlKk2zMPm
IWJ3Uv9GhpWdstvYGoEJopM4JgJPmFL/b5ofsNHsFbDibAAX8kd6q4PcOLN6l9r3aRDPnCHF/ii2
qmOAsewqAxf2KzUg/5Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e+Zq7fugn2wn+NfK5MiyV4wTKif0oJK70iDNbPgK9Tu4FyFu07ueWrGS5pD2q6K2tu9WtojoIChW
uICG//4++w6VSxcfgkBx7eZaM9hvR4Y8gO2p7mS55QvjOtpNJA1gNRrLov8ye17vOZSia6k6oLES
ua5ykV+u060fAK6Ky6zybSpGuN0/aRWsbIaVUG4sHjoSdG0nHF0DTJp8yqbDMilUcFeGiJ0f6v6+
O6cb4N3YlgTJrbbLpV3qOQmRJNdCBscqnWMXx5JcE0ujjHQOE2NRC9BkaxY/fC7bBsQIY1ZpnNOG
CwsmlCNaT5x9TTrVasF+4aqG4l1M99iERs95Bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`pragma protect data_block
3dBDzv38LYSblodwRBnvEANl43nPq5xQmvf7PS+q3NxQu8fzKEq4KzrFhfqft+S6kup7sY38v3Vt
NFbHGpAIXWkx98cITn7DEDsHq9V9mE3LOUzl4u2ujiv+DWMOVKXTjbR6aw1I1o2oCCYo3DMr3JxN
/PQC4EAuEKjsggMCvAyLh3FiJaxw5U6oBefgdTtQtLBaA4mXOyChQCngldFWZgNlPtgYRkNav9Zv
GFJtZ83/B7JBWC1r81ECoiEIqRMkhgSv+lxoaXqqkWMeM7P/XB7c74PFZuJr9K78sF9r3mjVJlit
yA+a/z10R4lbp4hbYcwii96NlBnqpP24LROz+PUEqYlAyND2FLmeGh0LTzEx3IFOGh7J2honTyvT
U83VkicOqfXWkexASnkT3bkjmUmyVM7qCtsukptmdOyvP3gX/qtTgeBwFxOidp21Im9kw+fTpaFb
HmifCJK5HEr3kM8zDrtWjUECcPENMafwUe3h2VYcjv5sKzMV4V+sQDyw7qNFgtjTHJv1VQkyuRKr
r8XbhGA/DZiohy8JNgsKS/tiSyiXgctTsThqD7NsIw1/ebf3LBVR98yydVVEnfSwMqBH0xQrhYlN
ev6zCJ2sLkzK6IyAx5zD2tcgV8uPgYzsIDzYq75VPplgix7kX8rpuUnDG4pdiePPNo4ezbuUL+9c
wQ/h0/M2AQ65ZS13GbW3ivdLy8NnO+kZ0VIprDycMK3w8ROKSgwz+eQ2n8WjYooSIqr0ZSTK1VKf
TWU60XncAvwzTO5nAeYR14QLgVAfJZTWYMXKZqZ1n1nx365cUuhpN7YuV5Q9cqEuXhQcx8nSAx0S
HPKZ5Ql2PX5a83vmmK/18Hw14OwB86VLmYziZbOtJOCEtvgtfLoYp6/bgI4RF+Reu7rGsC9LAalV
ENegHGJwDZ8oatpt9I3KuhwBX6e1ov8qiF7BvCDKUI7KKL1W8FsLc9d5OPjxdk963Qr6xrBsj6vw
C4T48QcPEl9CgcxTAyxHGB7UdjFog7E+tZbckSikm3LEGh5znU5AXigHrQyQr3CQCzTj1ISxoqnn
62J4CQt+gYURCDoeeVFYrtNTmvbNPziMX/Vi8NhVbsWV02gk9DK/Fm37QUbsBc4kp3GrqTs9zAsp
8gB029N5HuIcXRjLrg1+dzV/R+tYdBukmUS2AAGyL12FAnyrcAzzO21RHwqwpvCv7WjqI/AD26sS
KPEIE3Ai5imXJzRnrMfcWDIb4Xwz6M3RifryaWUVuxPqGIan3nrGoiFllC4p3JPIlFOki/De9WoE
R94TIk7hDkdIy4RZ1N77wG1CG39rCg1g4Pgd+D2lSQVylNNxXxn/UfXzU7WJh3PmMHayF9eWcqPE
LSL5XYwgNc1dGMAdXJCJDPAXocecOlL1/pTnc+ndo6vjBkRbL4yRJ9iW4HEnJAHbJ6pug/xzw1ky
GlqTCsuUhY3zbfB1kxMlI9zxe3PmTD9OpxL7OmQzAazZeHFbi4Wspa4uwxyACkDv8Rkudyc8DLOq
9nagLXNViaZaK49uiuetdoxUuktXiqQnbzwp8JqJBmbxrpJlTdrBGAYfyk1JgfToFSTYM80fOgK+
QEA9HsG+Gn8KLCVrygG0FJG8rtkIOcMDnUemvXOBnvbOmygnobf//hXzapwBejcyRHwhg6VafBHL
66H4KZ8aR8GeEvXms9E1fCCvNNF7hqdnQzaQbEEiiQrk27wbQfHfZ6XtZ63CCEnQx9iES535nPAE
4E/4/oa9asvYGzgn2E14dJMk+YVIAvjYOxgx2Vt0RtyHYNbf8i50euQ9udo2fjkg3CDxrZ2+kEh3
lqLWBjdAndEWNWBEcTpANLFGUBsZH3D6sdysDSYBs6CS0Q5p4SzDwR9Kd/uHR+UoH74ho1Ws52A8
+lY8j7Ljz1AQiODXw3t57RIaTC+GdM2zmvC9vuklZSrYCVsM+T5IkZyJrSrhO2UW103oy5PTUH7g
3xDebByEkeJlVk13rOLJzK1Owi+dqWPGUYFOTGAl8PEdCbqvA14PXGnkxLQm4YgUKre0x4JgUDhi
2KcnkjoZP2ne84xkNhM3LGvdGVn/UHIbNqAsUhc4Zad7/c7rYsuPRHeKqwqt+xw02DtUkeDjKh5F
3DZZm/SuYL4r+e4TgOABkjG85hdWCydeNh1Mj2wB3nSFIteEI7CTnTh0+AqCayV+Rw3Y6QSZw6we
f11FSSX3fUVGo7MAP56tdY/FyapnYFqbiuBEe7cwu+uk44+QYvThfNhBxx/6gXEreSSyt/1xK8pY
6DQ2p6VhIwOtI2XGfihCmSDAEuZHHu+ij/V4Z0wt0FVo8kemwDQUKYCLhVcaylP27f/iOGVZflkb
sHfClwl6OnhWFRGHjHn9ibE1i0db1J0/q2Ei8YxTBt/0xJZ3RynBrFxuXU94UH2JRDxf3w/TfNA8
KBBoLiECp0q6ovtikZDa2FjG0xgsTzkZOTbuEmPMxAjvTzk/VoAesVXw0qpOwdoA/anLbqJ7iz1S
vmWiT68I9O1+wkRsvatf7ChovvcKg7kfVFkJJiBvvbK2winRA+IZ4vWPuz1/LImO+deqWsqxrbv1
URQbpYK0V+mqfiNMqeKwPZ2fCzTJhOMUlzrWxET3XfPkRTh9qgi+H7Ww3yzffpVGhx4x+/YMZ/+0
sTlVfIlfnlSx68Ac+d4TGNJ9a+Mz+bhT4z6oBS7tuYdhosVbcAR8KICbjvpKXCw60tYvio2QwkSi
dgTtx6L4+Vk1ZZ7u8mQ/bpnXfCM+LJQQVo5iy6YHEHh57V0vsYuiJvKjBNARmObmt4244MjAH4Zk
hrbOWj3BlTMfaNIQ2aRlVQZx1+QvD0TutikFi3/lcthqjEHSWbN8VBTU+Mszn7yHUERfvTXN2InC
c8Xu399BcMyO4qINGPa66r6tbN02/kwWkZgJhj91cqhsS39c04wNG+o5pAcFj/xB4pRIZgDk3yls
rTAy0Q+3aSBdyVYC7GxkNx7VpQE1J/59x2c2IqAuDkBjJx0hm6nlDF2dSgIDcaFnZ4r0vM9J2dCd
p6c9UuImoc2ZcNfxhnpZWXBVoBSMPUltKBmWF9iFR88o3um9KQIDD7uJ8QD1DX894nN6syBlzPVQ
Oug0i+Rb0aJ7FOFEu4TsiyG4c06zuftnR66Y9/NDvdE5LCTv6xnz/crdnMDOR2HLRsnxy2xZ3XVe
/a3GRRBg7jY+it3/QQyl4PEJOn4v61Ix9wKWVGFyzuNgCk9H23Pm4NBasEce02y66ME5RAneFnSP
FictBXxViscmfV7RqzAzNp1XizFZB8Jrl2msfOH473Xv0k413ZlInEw3Nj2Rryt0OsGfQ+dtrPhv
Ht8AQKLCRMaIFovUYi4XgjVfF7i0Y669jSmp4JaiBb6usHHTJ1WLGP7ohJFC+0ku4fw/WeydZNdL
lKv0fs+oIUS72MjZYCT3foYVqSGPmxHaEEK1AU5DRPa/OiO23HIxfDgXmdQv0QbeOrtW0kyl9Uuz
9UfwNidsuuedDxOjIr+Dohx0fqMJYUFQe3/wORQDlEPYrILJDDbGbzTcVHZQYuSelgr7v8uQ5UUl
nyJ1DyIHXA0+isZgk0disHNsDzNm3M0QoSxrE4K+zV6l0/MwD1D/3On/EEmdkpwH9lQWyFt8ovHT
4yuAJkeiU8cJdaL/caDXSdqtVWtqN31nAakgfkYiaOB2VTaGlmf0GfmiJ8XiAKYo5BcKgDyEwfFU
ZSzCLg+wUKRYuY/U0+dOcvDNimo7eiszt79h8XO4h9JEirrmBiYK/JCvBMINnr71/9/Mc6NoU1Ne
0hdXLqf7MwOP9+g75CZhmTso0zc0JsxoeLrK0Y/Qb5r8Rsx71hHb/2/iKilldiBukX7nJK2qrGzG
h2PMD8Sfobbu5Cs6EV7y7TOLlOx8kCCR7TqXZ4G2KF1Ljr8ehZpUO9HJckpsVm339xrmPRiqxGbm
pdLN+qstr+B9oKu6XVmOz29S4eRlNeumGKaq+2KpT7E8O44eon7m/+YEpBLsSBBGwEQDqHmtvuf8
mNEebl3yDbqo6RaQqsqtV2XD2xxORLzS58yKgo7f0OFgwQNxQNLdFDlh3SWZzAdghzwXlYgzDmzW
rmVZHB8Z6L0D2Kk6TStn1W4yP3kzncL0U2+f3K3pqMzVAT4qb3QoAs2qIEDtbKitoCLinnP5X9VK
uQtYJTQ/I73Es3NrBfqJDIWZXq2CRoLERM2QzhcEuV7/D7FVMR61Oh8Yndon8Mnv/93zk079HmV3
2wXTnyiSJcfyBMkuN0srGH6i4SsD4aCq7/B70GXqS9wVVj71Jtj2W/asK0C95GYmZw0PPeT3Bod5
mBwP0vPk5Id/SP6RhAFaDgCyfohuqHjG+7EqvFim9zO+F0oDaxOIXgJZf2He77ZzJvZ29y1g5B3X
qt/55RL4BB13PJ+eDzpXBOuxTr/MbKG04a5tIXlMiZBF6jmLZRNlRFguxT7C7IEFdOEYJV4wqPY1
h4VSVq+mGCfC2oYhdw/WCBaQLfG7ovZy/qBCWlvlEa6YOGIKBbTdGKRSbravsW5jCEI9pvXVy2sX
VZTG90BdsRkKvGOIWuApJyIUrqrAXjvsEJNsFji1hK3EfimXQ3Fc15p8io1895VAj6Q7CA3PcXrf
+LS3VuFZS9YZuaHSdCRanLTZIeBRXK3inBFssP/q0cM7wHfJXWc6STkFDFZWcR9JHSc6VqoQteSC
9keutXKuXdaNLw9JRMN521Y7fD/IB4j3hZvSW8W4KvcVNIyFQtvEVTZQ0SxZCRdgWPss+kPRqrBg
DWGiR7AqOMEd6HLOiQCDKfmexdUmHRL6vhNBb6lEEM32VxmcFWVHyq9YRCOSIMpYdnsPJsUqXHwL
ca3SpGIU9mtRplIKqyNBmUQc67lmHuXHUmel/KdoC8Fsya2bX3YHc7KYzLyTSKNC1lkEngGr4KXH
PAbOGx/fJt4eIS6DXvI9eZxEp10SoxKK6nnE2HUUYSniaLUhzuSAkwSfGBJHesCzkWq62DOG6ddY
OsLeycRH6hbqZTQaRUKC1jurMQ94i9w2apOHjvuWD+uQ9+BMMCDroTzF39xRR7t3WMu12n526635
xNfA0gXGfEbTxPCqAGkJnLzKryZtN5nOovLDeHbz8cYgOZCsYpKdF973evgQuN3Eh+rrdoW3ubIB
y82P8RVasXZAssjLQx2app+iOmOYJhkBjcOkKsODwCARP2amJbHKt2PV+uP+5MOLUU8l3YcpTc5y
8J/BfUBlLmBguh/iSpIgbwFFV+Ml0vz+iQl0CCY2SPe08RLnAwZRM9bNuw0fASRS0tDVepI7ZRR4
pF/R3mDk00OZGAQSCno4xY6CTnfvP1h60wuIQjl331DkgGHpjSKu8sgKG0O5sn2sWHm5K7ZULN63
ruJyKgFppUrkkX1eL7RztBsrP/fzBQ8jFaa+5EByzR2pv6x8xQoi7R6OciZ5ltmKKAdYoSQD6KYz
FwnL96SI2KeaEhGJaPKAsiVDTpLQ1g5v12ATHMJmHVc9yFY3EsT1sxzYYwtAq0GW17FL1IyStB3u
hqErBpflyQObwfSwA8SB/HTZWAlWjYHumTFLhwEzN2Qcn/Jynq477bXcL6PiFcZ4RnKq8wMphaIz
Ed9fF69YL/HcxKFvZ02Zxgfo5tWbucC6jKLL+YOr2ZC13k2dnIYj4YdDGfQfjHB1cG9dOO908qrm
bSocYLSljlry2NMapezhuhM5Nkf4qPnOv/yqz8au0VCfkZ7RgaulOwZUxIXiYH8la0ObhGJDRxLI
fe7NhiZYBtOwEyn48aBhsL7vQCoaOAN5AxbgAdUkoJqAg6xNp+mUurDdSRIt94kUDy2IQ3Z513WN
DcIEu/T/xGS2EzOJ83wm9UpnaXs1SpMY866X6wf7LjVgDs/SkvUOYXmAtANYyX6bJPbmv3LigUZg
gtbGSWXgV0am4sXN8YpLmB0hOn8WBeOZh7IkSV+NTvxwsqFOAE1sf/NVUOpUDRzrwquvD/4UtD2p
JdiqEpQZijW3QGqnPsdvPPwXbZRVPJQu18RegXX8GuP3UnXhvZeX+ySRptWc9sGPAn7aYwqItam0
JjU+x5HD+uFqwwmb2ztf+me6Vek5RxzZE7gswo3koRR7/m0xI9bVsryAKJ8/6vA0mkTPocgMF2l9
ewPa3khLH12hwFVbyKxBLfs8a933hCDeScdC3t1plgqFeh/MEcvuQcnB62BDWf8C/y4BNPm0W/I8
FW+DR5fpICBQh1SUaYTuLivnYRIVfT0wWlvlkTE2o+C6b7CExlUM668rfRwCohmTR/HQn1iJ/cL/
rTkW7/sK414Xbs6sZOE0ZJ7ZRVGNDi3zwSnzsqw+tpWVO12F5s84G+k0mrMo3VQkbkBcU3h6dmox
REP2X7TrMYQNOmvd0VWLDDBs0dlmOs5Sp6W+/83H8gcyBU02+28aEiesbV1KJpmJbOduelU48qUM
lhZm8aKRbcksj7B9muRGJrc9ifBPSjc0i3Abrzt2n8pG7JZBhkWMnBn3la6jXyuK1as0R9lXq2UH
f6co/8dock66HaUDxk9wSHBxCox9N2P+f5pnnKVcwxlcc9d3Q8frk0pYNUkkjVbnUN7Vrq80/xMK
qXY8Cgo952l0nvwnxRAmtdXtoquUkmA1shyURYcFqcXaTXJ/9T/oxqGq7B2bQ72V8P+k6MCtQQs1
TqCfCr7MGzNUq6aYB6GlQt9LLCPe9F12kXkrNaZGs+mOytBtOj2kDz1pse0eK2ceKPnqqhjE+jo6
k2AjvCPjW5Ezrtqs0eHLc6RV1webMm7ZJvrZSNdyevX4jaUdYUiPnkvftff17+aAGNNasPIsHq4s
55za2QCo8nphNVyMCE80tAgYwEiJNf8pJ/sOpyBNoGSTIQQm0zY/ozqkv3sXLSpT0vO15W37f5jG
SSPL3AAJJ8AmhMBes+Fdjp3o1ZnnOm3TegBuARpneoUtQ5Qt1y0M3cUl60GNdF0fLsldj6u2loa7
iyRn4Q==
`pragma protect end_protected
